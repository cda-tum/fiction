// Benchmark "b18" written by ABC on Wed Sep  5 10:17:21 2018

module b18 ( clock, 
    HOLD, NA, BS, SEL, DIN_31_, DIN_30_, DIN_29_, DIN_28_, DIN_27_,
    DIN_26_, DIN_25_, DIN_24_, DIN_23_, DIN_22_, DIN_21_, DIN_20_, DIN_19_,
    DIN_18_, DIN_17_, DIN_16_, DIN_15_, DIN_14_, DIN_13_, DIN_12_, DIN_11_,
    DIN_10_, DIN_9_, DIN_8_, DIN_7_, DIN_6_, DIN_5_, DIN_4_, DIN_3_,
    DIN_2_, DIN_1_, DIN_0_, LOGIC0,
    MUL_1411_U378, MUL_1411_U438, MUL_1411_U10, MUL_1411_U439, MUL_1411_U9,
    MUL_1411_U440, MUL_1411_U8, MUL_1411_U441, MUL_1411_U7, MUL_1411_U385,
    MUL_1411_U14, MUL_1411_U386, MUL_1411_U13, MUL_1411_U387, MUL_1411_U12,
    MUL_1411_U388, MUL_1411_U11, MUL_1411_U15, MUL_1411_U5, MUL_1421_A1_U5,
    U154, U39  );
  input  clock;
  input  HOLD, NA, BS, SEL, DIN_31_, DIN_30_, DIN_29_, DIN_28_, DIN_27_,
    DIN_26_, DIN_25_, DIN_24_, DIN_23_, DIN_22_, DIN_21_, DIN_20_, DIN_19_,
    DIN_18_, DIN_17_, DIN_16_, DIN_15_, DIN_14_, DIN_13_, DIN_12_, DIN_11_,
    DIN_10_, DIN_9_, DIN_8_, DIN_7_, DIN_6_, DIN_5_, DIN_4_, DIN_3_,
    DIN_2_, DIN_1_, DIN_0_, LOGIC0;
  output MUL_1411_U378, MUL_1411_U438, MUL_1411_U10, MUL_1411_U439,
    MUL_1411_U9, MUL_1411_U440, MUL_1411_U8, MUL_1411_U441, MUL_1411_U7,
    MUL_1411_U385, MUL_1411_U14, MUL_1411_U386, MUL_1411_U13,
    MUL_1411_U387, MUL_1411_U12, MUL_1411_U388, MUL_1411_U11, MUL_1411_U15,
    MUL_1411_U5, MUL_1421_A1_U5, U154, U39;
  reg P1_BUF1_REG_0_, P1_BUF1_REG_1_, P1_BUF1_REG_2_, P1_BUF1_REG_3_,
    P1_BUF1_REG_4_, P1_BUF1_REG_5_, P1_BUF1_REG_6_, P1_BUF1_REG_7_,
    P1_BUF1_REG_8_, P1_BUF1_REG_9_, P1_BUF1_REG_10_, P1_BUF1_REG_11_,
    P1_BUF1_REG_12_, P1_BUF1_REG_13_, P1_BUF1_REG_14_, P1_BUF1_REG_15_,
    P1_BUF1_REG_16_, P1_BUF1_REG_17_, P1_BUF1_REG_18_, P1_BUF1_REG_19_,
    P1_BUF1_REG_20_, P1_BUF1_REG_21_, P1_BUF1_REG_22_, P1_BUF1_REG_23_,
    P1_BUF1_REG_24_, P1_BUF1_REG_25_, P1_BUF1_REG_26_, P1_BUF1_REG_27_,
    P1_BUF1_REG_28_, P1_BUF1_REG_29_, P1_BUF1_REG_30_, P1_BUF1_REG_31_,
    P1_BUF2_REG_0_, P1_BUF2_REG_1_, P1_BUF2_REG_2_, P1_BUF2_REG_3_,
    P1_BUF2_REG_4_, P1_BUF2_REG_5_, P1_BUF2_REG_6_, P1_BUF2_REG_7_,
    P1_BUF2_REG_8_, P1_BUF2_REG_9_, P1_BUF2_REG_10_, P1_BUF2_REG_11_,
    P1_BUF2_REG_12_, P1_BUF2_REG_13_, P1_BUF2_REG_14_, P1_BUF2_REG_15_,
    P1_BUF2_REG_16_, P1_BUF2_REG_17_, P1_BUF2_REG_18_, P1_BUF2_REG_19_,
    P1_BUF2_REG_20_, P1_BUF2_REG_21_, P1_BUF2_REG_22_, P1_BUF2_REG_23_,
    P1_BUF2_REG_24_, P1_BUF2_REG_25_, P1_BUF2_REG_26_, P1_BUF2_REG_27_,
    P1_BUF2_REG_28_, P1_BUF2_REG_29_, P1_BUF2_REG_30_, P1_BUF2_REG_31_,
    P1_READY12_REG, P1_READY21_REG, P1_READY22_REG, P1_READY11_REG,
    P2_BUF1_REG_0_, P2_BUF1_REG_1_, P2_BUF1_REG_2_, P2_BUF1_REG_3_,
    P2_BUF1_REG_4_, P2_BUF1_REG_5_, P2_BUF1_REG_6_, P2_BUF1_REG_7_,
    P2_BUF1_REG_8_, P2_BUF1_REG_9_, P2_BUF1_REG_10_, P2_BUF1_REG_11_,
    P2_BUF1_REG_12_, P2_BUF1_REG_13_, P2_BUF1_REG_14_, P2_BUF1_REG_15_,
    P2_BUF1_REG_16_, P2_BUF1_REG_17_, P2_BUF1_REG_18_, P2_BUF1_REG_19_,
    P2_BUF1_REG_20_, P2_BUF1_REG_21_, P2_BUF1_REG_22_, P2_BUF1_REG_23_,
    P2_BUF1_REG_24_, P2_BUF1_REG_25_, P2_BUF1_REG_26_, P2_BUF1_REG_27_,
    P2_BUF1_REG_28_, P2_BUF1_REG_29_, P2_BUF1_REG_30_, P2_BUF1_REG_31_,
    P2_BUF2_REG_0_, P2_BUF2_REG_1_, P2_BUF2_REG_2_, P2_BUF2_REG_3_,
    P2_BUF2_REG_4_, P2_BUF2_REG_5_, P2_BUF2_REG_6_, P2_BUF2_REG_7_,
    P2_BUF2_REG_8_, P2_BUF2_REG_9_, P2_BUF2_REG_10_, P2_BUF2_REG_11_,
    P2_BUF2_REG_12_, P2_BUF2_REG_13_, P2_BUF2_REG_14_, P2_BUF2_REG_15_,
    P2_BUF2_REG_16_, P2_BUF2_REG_17_, P2_BUF2_REG_18_, P2_BUF2_REG_19_,
    P2_BUF2_REG_20_, P2_BUF2_REG_21_, P2_BUF2_REG_22_, P2_BUF2_REG_23_,
    P2_BUF2_REG_24_, P2_BUF2_REG_25_, P2_BUF2_REG_26_, P2_BUF2_REG_27_,
    P2_BUF2_REG_28_, P2_BUF2_REG_29_, P2_BUF2_REG_30_, P2_BUF2_REG_31_,
    P2_READY12_REG, P2_READY21_REG, P2_READY22_REG, P2_READY11_REG,
    P3_IR_REG_0_, P3_IR_REG_1_, P3_IR_REG_2_, P3_IR_REG_3_, P3_IR_REG_4_,
    P3_IR_REG_5_, P3_IR_REG_6_, P3_IR_REG_7_, P3_IR_REG_8_, P3_IR_REG_9_,
    P3_IR_REG_10_, P3_IR_REG_11_, P3_IR_REG_12_, P3_IR_REG_13_,
    P3_IR_REG_14_, P3_IR_REG_15_, P3_IR_REG_16_, P3_IR_REG_17_,
    P3_IR_REG_18_, P3_IR_REG_19_, P3_IR_REG_20_, P3_IR_REG_21_,
    P3_IR_REG_22_, P3_IR_REG_23_, P3_IR_REG_24_, P3_IR_REG_25_,
    P3_IR_REG_26_, P3_IR_REG_27_, P3_IR_REG_28_, P3_IR_REG_29_,
    P3_IR_REG_30_, P3_IR_REG_31_, P3_D_REG_0_, P3_D_REG_1_, P3_D_REG_2_,
    P3_D_REG_3_, P3_D_REG_4_, P3_D_REG_5_, P3_D_REG_6_, P3_D_REG_7_,
    P3_D_REG_8_, P3_D_REG_9_, P3_D_REG_10_, P3_D_REG_11_, P3_D_REG_12_,
    P3_D_REG_13_, P3_D_REG_14_, P3_D_REG_15_, P3_D_REG_16_, P3_D_REG_17_,
    P3_D_REG_18_, P3_D_REG_19_, P3_D_REG_20_, P3_D_REG_21_, P3_D_REG_22_,
    P3_D_REG_23_, P3_D_REG_24_, P3_D_REG_25_, P3_D_REG_26_, P3_D_REG_27_,
    P3_D_REG_28_, P3_D_REG_29_, P3_D_REG_30_, P3_D_REG_31_, P3_REG0_REG_0_,
    P3_REG0_REG_1_, P3_REG0_REG_2_, P3_REG0_REG_3_, P3_REG0_REG_4_,
    P3_REG0_REG_5_, P3_REG0_REG_6_, P3_REG0_REG_7_, P3_REG0_REG_8_,
    P3_REG0_REG_9_, P3_REG0_REG_10_, P3_REG0_REG_11_, P3_REG0_REG_12_,
    P3_REG0_REG_13_, P3_REG0_REG_14_, P3_REG0_REG_15_, P3_REG0_REG_16_,
    P3_REG0_REG_17_, P3_REG0_REG_18_, P3_REG0_REG_19_, P3_REG0_REG_20_,
    P3_REG0_REG_21_, P3_REG0_REG_22_, P3_REG0_REG_23_, P3_REG0_REG_24_,
    P3_REG0_REG_25_, P3_REG0_REG_26_, P3_REG0_REG_27_, P3_REG0_REG_28_,
    P3_REG0_REG_29_, P3_REG0_REG_30_, P3_REG0_REG_31_, P3_REG1_REG_0_,
    P3_REG1_REG_1_, P3_REG1_REG_2_, P3_REG1_REG_3_, P3_REG1_REG_4_,
    P3_REG1_REG_5_, P3_REG1_REG_6_, P3_REG1_REG_7_, P3_REG1_REG_8_,
    P3_REG1_REG_9_, P3_REG1_REG_10_, P3_REG1_REG_11_, P3_REG1_REG_12_,
    P3_REG1_REG_13_, P3_REG1_REG_14_, P3_REG1_REG_15_, P3_REG1_REG_16_,
    P3_REG1_REG_17_, P3_REG1_REG_18_, P3_REG1_REG_19_, P3_REG1_REG_20_,
    P3_REG1_REG_21_, P3_REG1_REG_22_, P3_REG1_REG_23_, P3_REG1_REG_24_,
    P3_REG1_REG_25_, P3_REG1_REG_26_, P3_REG1_REG_27_, P3_REG1_REG_28_,
    P3_REG1_REG_29_, P3_REG1_REG_30_, P3_REG1_REG_31_, P3_REG2_REG_0_,
    P3_REG2_REG_1_, P3_REG2_REG_2_, P3_REG2_REG_3_, P3_REG2_REG_4_,
    P3_REG2_REG_5_, P3_REG2_REG_6_, P3_REG2_REG_7_, P3_REG2_REG_8_,
    P3_REG2_REG_9_, P3_REG2_REG_10_, P3_REG2_REG_11_, P3_REG2_REG_12_,
    P3_REG2_REG_13_, P3_REG2_REG_14_, P3_REG2_REG_15_, P3_REG2_REG_16_,
    P3_REG2_REG_17_, P3_REG2_REG_18_, P3_REG2_REG_19_, P3_REG2_REG_20_,
    P3_REG2_REG_21_, P3_REG2_REG_22_, P3_REG2_REG_23_, P3_REG2_REG_24_,
    P3_REG2_REG_25_, P3_REG2_REG_26_, P3_REG2_REG_27_, P3_REG2_REG_28_,
    P3_REG2_REG_29_, P3_REG2_REG_30_, P3_REG2_REG_31_, P3_ADDR_REG_19_,
    P3_ADDR_REG_18_, P3_ADDR_REG_17_, P3_ADDR_REG_16_, P3_ADDR_REG_15_,
    P3_ADDR_REG_14_, P3_ADDR_REG_13_, P3_ADDR_REG_12_, P3_ADDR_REG_11_,
    P3_ADDR_REG_10_, P3_ADDR_REG_9_, P3_ADDR_REG_8_, P3_ADDR_REG_7_,
    P3_ADDR_REG_6_, P3_ADDR_REG_5_, P3_ADDR_REG_4_, P3_ADDR_REG_3_,
    P3_ADDR_REG_2_, P3_ADDR_REG_1_, P3_ADDR_REG_0_, P3_DATAO_REG_0_,
    P3_DATAO_REG_1_, P3_DATAO_REG_2_, P3_DATAO_REG_3_, P3_DATAO_REG_4_,
    P3_DATAO_REG_5_, P3_DATAO_REG_6_, P3_DATAO_REG_7_, P3_DATAO_REG_8_,
    P3_DATAO_REG_9_, P3_DATAO_REG_10_, P3_DATAO_REG_11_, P3_DATAO_REG_12_,
    P3_DATAO_REG_13_, P3_DATAO_REG_14_, P3_DATAO_REG_15_, P3_DATAO_REG_16_,
    P3_DATAO_REG_17_, P3_DATAO_REG_18_, P3_DATAO_REG_19_, P3_DATAO_REG_20_,
    P3_DATAO_REG_21_, P3_DATAO_REG_22_, P3_DATAO_REG_23_, P3_DATAO_REG_24_,
    P3_DATAO_REG_25_, P3_DATAO_REG_26_, P3_DATAO_REG_27_, P3_DATAO_REG_28_,
    P3_DATAO_REG_29_, P3_DATAO_REG_30_, P3_DATAO_REG_31_, P3_B_REG,
    P3_REG3_REG_15_, P3_REG3_REG_26_, P3_REG3_REG_6_, P3_REG3_REG_18_,
    P3_REG3_REG_2_, P3_REG3_REG_11_, P3_REG3_REG_22_, P3_REG3_REG_13_,
    P3_REG3_REG_20_, P3_REG3_REG_0_, P3_REG3_REG_9_, P3_REG3_REG_4_,
    P3_REG3_REG_24_, P3_REG3_REG_17_, P3_REG3_REG_5_, P3_REG3_REG_16_,
    P3_REG3_REG_25_, P3_REG3_REG_12_, P3_REG3_REG_21_, P3_REG3_REG_1_,
    P3_REG3_REG_8_, P3_REG3_REG_28_, P3_REG3_REG_19_, P3_REG3_REG_3_,
    P3_REG3_REG_10_, P3_REG3_REG_23_, P3_REG3_REG_14_, P3_REG3_REG_27_,
    P3_REG3_REG_7_, P3_STATE_REG, P3_RD_REG, P3_WR_REG, P4_IR_REG_0_,
    P4_IR_REG_1_, P4_IR_REG_2_, P4_IR_REG_3_, P4_IR_REG_4_, P4_IR_REG_5_,
    P4_IR_REG_6_, P4_IR_REG_7_, P4_IR_REG_8_, P4_IR_REG_9_, P4_IR_REG_10_,
    P4_IR_REG_11_, P4_IR_REG_12_, P4_IR_REG_13_, P4_IR_REG_14_,
    P4_IR_REG_15_, P4_IR_REG_16_, P4_IR_REG_17_, P4_IR_REG_18_,
    P4_IR_REG_19_, P4_IR_REG_20_, P4_IR_REG_21_, P4_IR_REG_22_,
    P4_IR_REG_23_, P4_IR_REG_24_, P4_IR_REG_25_, P4_IR_REG_26_,
    P4_IR_REG_27_, P4_IR_REG_28_, P4_IR_REG_29_, P4_IR_REG_30_,
    P4_IR_REG_31_, P4_D_REG_0_, P4_D_REG_1_, P4_D_REG_2_, P4_D_REG_3_,
    P4_D_REG_4_, P4_D_REG_5_, P4_D_REG_6_, P4_D_REG_7_, P4_D_REG_8_,
    P4_D_REG_9_, P4_D_REG_10_, P4_D_REG_11_, P4_D_REG_12_, P4_D_REG_13_,
    P4_D_REG_14_, P4_D_REG_15_, P4_D_REG_16_, P4_D_REG_17_, P4_D_REG_18_,
    P4_D_REG_19_, P4_D_REG_20_, P4_D_REG_21_, P4_D_REG_22_, P4_D_REG_23_,
    P4_D_REG_24_, P4_D_REG_25_, P4_D_REG_26_, P4_D_REG_27_, P4_D_REG_28_,
    P4_D_REG_29_, P4_D_REG_30_, P4_D_REG_31_, P4_REG0_REG_0_,
    P4_REG0_REG_1_, P4_REG0_REG_2_, P4_REG0_REG_3_, P4_REG0_REG_4_,
    P4_REG0_REG_5_, P4_REG0_REG_6_, P4_REG0_REG_7_, P4_REG0_REG_8_,
    P4_REG0_REG_9_, P4_REG0_REG_10_, P4_REG0_REG_11_, P4_REG0_REG_12_,
    P4_REG0_REG_13_, P4_REG0_REG_14_, P4_REG0_REG_15_, P4_REG0_REG_16_,
    P4_REG0_REG_17_, P4_REG0_REG_18_, P4_REG0_REG_19_, P4_REG0_REG_20_,
    P4_REG0_REG_21_, P4_REG0_REG_22_, P4_REG0_REG_23_, P4_REG0_REG_24_,
    P4_REG0_REG_25_, P4_REG0_REG_26_, P4_REG0_REG_27_, P4_REG0_REG_28_,
    P4_REG0_REG_29_, P4_REG0_REG_30_, P4_REG0_REG_31_, P4_REG1_REG_0_,
    P4_REG1_REG_1_, P4_REG1_REG_2_, P4_REG1_REG_3_, P4_REG1_REG_4_,
    P4_REG1_REG_5_, P4_REG1_REG_6_, P4_REG1_REG_7_, P4_REG1_REG_8_,
    P4_REG1_REG_9_, P4_REG1_REG_10_, P4_REG1_REG_11_, P4_REG1_REG_12_,
    P4_REG1_REG_13_, P4_REG1_REG_14_, P4_REG1_REG_15_, P4_REG1_REG_16_,
    P4_REG1_REG_17_, P4_REG1_REG_18_, P4_REG1_REG_19_, P4_REG1_REG_20_,
    P4_REG1_REG_21_, P4_REG1_REG_22_, P4_REG1_REG_23_, P4_REG1_REG_24_,
    P4_REG1_REG_25_, P4_REG1_REG_26_, P4_REG1_REG_27_, P4_REG1_REG_28_,
    P4_REG1_REG_29_, P4_REG1_REG_30_, P4_REG1_REG_31_, P4_REG2_REG_0_,
    P4_REG2_REG_1_, P4_REG2_REG_2_, P4_REG2_REG_3_, P4_REG2_REG_4_,
    P4_REG2_REG_5_, P4_REG2_REG_6_, P4_REG2_REG_7_, P4_REG2_REG_8_,
    P4_REG2_REG_9_, P4_REG2_REG_10_, P4_REG2_REG_11_, P4_REG2_REG_12_,
    P4_REG2_REG_13_, P4_REG2_REG_14_, P4_REG2_REG_15_, P4_REG2_REG_16_,
    P4_REG2_REG_17_, P4_REG2_REG_18_, P4_REG2_REG_19_, P4_REG2_REG_20_,
    P4_REG2_REG_21_, P4_REG2_REG_22_, P4_REG2_REG_23_, P4_REG2_REG_24_,
    P4_REG2_REG_25_, P4_REG2_REG_26_, P4_REG2_REG_27_, P4_REG2_REG_28_,
    P4_REG2_REG_29_, P4_REG2_REG_30_, P4_REG2_REG_31_, P4_ADDR_REG_19_,
    P4_ADDR_REG_18_, P4_ADDR_REG_17_, P4_ADDR_REG_16_, P4_ADDR_REG_15_,
    P4_ADDR_REG_14_, P4_ADDR_REG_13_, P4_ADDR_REG_12_, P4_ADDR_REG_11_,
    P4_ADDR_REG_10_, P4_ADDR_REG_9_, P4_ADDR_REG_8_, P4_ADDR_REG_7_,
    P4_ADDR_REG_6_, P4_ADDR_REG_5_, P4_ADDR_REG_4_, P4_ADDR_REG_3_,
    P4_ADDR_REG_2_, P4_ADDR_REG_1_, P4_ADDR_REG_0_, P4_DATAO_REG_0_,
    P4_DATAO_REG_1_, P4_DATAO_REG_2_, P4_DATAO_REG_3_, P4_DATAO_REG_4_,
    P4_DATAO_REG_5_, P4_DATAO_REG_6_, P4_DATAO_REG_7_, P4_DATAO_REG_8_,
    P4_DATAO_REG_9_, P4_DATAO_REG_10_, P4_DATAO_REG_11_, P4_DATAO_REG_12_,
    P4_DATAO_REG_13_, P4_DATAO_REG_14_, P4_DATAO_REG_15_, P4_DATAO_REG_16_,
    P4_DATAO_REG_17_, P4_DATAO_REG_18_, P4_DATAO_REG_19_, P4_DATAO_REG_20_,
    P4_DATAO_REG_21_, P4_DATAO_REG_22_, P4_DATAO_REG_23_, P4_DATAO_REG_24_,
    P4_DATAO_REG_25_, P4_DATAO_REG_26_, P4_DATAO_REG_27_, P4_DATAO_REG_28_,
    P4_DATAO_REG_29_, P4_DATAO_REG_30_, P4_DATAO_REG_31_, P4_B_REG,
    P4_REG3_REG_15_, P4_REG3_REG_26_, P4_REG3_REG_6_, P4_REG3_REG_18_,
    P4_REG3_REG_2_, P4_REG3_REG_11_, P4_REG3_REG_22_, P4_REG3_REG_13_,
    P4_REG3_REG_20_, P4_REG3_REG_0_, P4_REG3_REG_9_, P4_REG3_REG_4_,
    P4_REG3_REG_24_, P4_REG3_REG_17_, P4_REG3_REG_5_, P4_REG3_REG_16_,
    P4_REG3_REG_25_, P4_REG3_REG_12_, P4_REG3_REG_21_, P4_REG3_REG_1_,
    P4_REG3_REG_8_, P4_REG3_REG_28_, P4_REG3_REG_19_, P4_REG3_REG_3_,
    P4_REG3_REG_10_, P4_REG3_REG_23_, P4_REG3_REG_14_, P4_REG3_REG_27_,
    P4_REG3_REG_7_, P4_STATE_REG, P4_RD_REG, P4_WR_REG, P1_P3_BE_N_REG_3_,
    P1_P3_BE_N_REG_2_, P1_P3_BE_N_REG_1_, P1_P3_BE_N_REG_0_,
    P1_P3_ADDRESS_REG_29_, P1_P3_ADDRESS_REG_28_, P1_P3_ADDRESS_REG_27_,
    P1_P3_ADDRESS_REG_26_, P1_P3_ADDRESS_REG_25_, P1_P3_ADDRESS_REG_24_,
    P1_P3_ADDRESS_REG_23_, P1_P3_ADDRESS_REG_22_, P1_P3_ADDRESS_REG_21_,
    P1_P3_ADDRESS_REG_20_, P1_P3_ADDRESS_REG_19_, P1_P3_ADDRESS_REG_18_,
    P1_P3_ADDRESS_REG_17_, P1_P3_ADDRESS_REG_16_, P1_P3_ADDRESS_REG_15_,
    P1_P3_ADDRESS_REG_14_, P1_P3_ADDRESS_REG_13_, P1_P3_ADDRESS_REG_12_,
    P1_P3_ADDRESS_REG_11_, P1_P3_ADDRESS_REG_10_, P1_P3_ADDRESS_REG_9_,
    P1_P3_ADDRESS_REG_8_, P1_P3_ADDRESS_REG_7_, P1_P3_ADDRESS_REG_6_,
    P1_P3_ADDRESS_REG_5_, P1_P3_ADDRESS_REG_4_, P1_P3_ADDRESS_REG_3_,
    P1_P3_ADDRESS_REG_2_, P1_P3_ADDRESS_REG_1_, P1_P3_ADDRESS_REG_0_,
    P1_P3_STATE_REG_2_, P1_P3_STATE_REG_1_, P1_P3_STATE_REG_0_,
    P1_P3_DATAWIDTH_REG_0_, P1_P3_DATAWIDTH_REG_1_, P1_P3_DATAWIDTH_REG_2_,
    P1_P3_DATAWIDTH_REG_3_, P1_P3_DATAWIDTH_REG_4_, P1_P3_DATAWIDTH_REG_5_,
    P1_P3_DATAWIDTH_REG_6_, P1_P3_DATAWIDTH_REG_7_, P1_P3_DATAWIDTH_REG_8_,
    P1_P3_DATAWIDTH_REG_9_, P1_P3_DATAWIDTH_REG_10_,
    P1_P3_DATAWIDTH_REG_11_, P1_P3_DATAWIDTH_REG_12_,
    P1_P3_DATAWIDTH_REG_13_, P1_P3_DATAWIDTH_REG_14_,
    P1_P3_DATAWIDTH_REG_15_, P1_P3_DATAWIDTH_REG_16_,
    P1_P3_DATAWIDTH_REG_17_, P1_P3_DATAWIDTH_REG_18_,
    P1_P3_DATAWIDTH_REG_19_, P1_P3_DATAWIDTH_REG_20_,
    P1_P3_DATAWIDTH_REG_21_, P1_P3_DATAWIDTH_REG_22_,
    P1_P3_DATAWIDTH_REG_23_, P1_P3_DATAWIDTH_REG_24_,
    P1_P3_DATAWIDTH_REG_25_, P1_P3_DATAWIDTH_REG_26_,
    P1_P3_DATAWIDTH_REG_27_, P1_P3_DATAWIDTH_REG_28_,
    P1_P3_DATAWIDTH_REG_29_, P1_P3_DATAWIDTH_REG_30_,
    P1_P3_DATAWIDTH_REG_31_, P1_P3_STATE2_REG_3_, P1_P3_STATE2_REG_2_,
    P1_P3_STATE2_REG_1_, P1_P3_STATE2_REG_0_, P1_P3_INSTQUEUE_REG_15__7_,
    P1_P3_INSTQUEUE_REG_15__6_, P1_P3_INSTQUEUE_REG_15__5_,
    P1_P3_INSTQUEUE_REG_15__4_, P1_P3_INSTQUEUE_REG_15__3_,
    P1_P3_INSTQUEUE_REG_15__2_, P1_P3_INSTQUEUE_REG_15__1_,
    P1_P3_INSTQUEUE_REG_15__0_, P1_P3_INSTQUEUE_REG_14__7_,
    P1_P3_INSTQUEUE_REG_14__6_, P1_P3_INSTQUEUE_REG_14__5_,
    P1_P3_INSTQUEUE_REG_14__4_, P1_P3_INSTQUEUE_REG_14__3_,
    P1_P3_INSTQUEUE_REG_14__2_, P1_P3_INSTQUEUE_REG_14__1_,
    P1_P3_INSTQUEUE_REG_14__0_, P1_P3_INSTQUEUE_REG_13__7_,
    P1_P3_INSTQUEUE_REG_13__6_, P1_P3_INSTQUEUE_REG_13__5_,
    P1_P3_INSTQUEUE_REG_13__4_, P1_P3_INSTQUEUE_REG_13__3_,
    P1_P3_INSTQUEUE_REG_13__2_, P1_P3_INSTQUEUE_REG_13__1_,
    P1_P3_INSTQUEUE_REG_13__0_, P1_P3_INSTQUEUE_REG_12__7_,
    P1_P3_INSTQUEUE_REG_12__6_, P1_P3_INSTQUEUE_REG_12__5_,
    P1_P3_INSTQUEUE_REG_12__4_, P1_P3_INSTQUEUE_REG_12__3_,
    P1_P3_INSTQUEUE_REG_12__2_, P1_P3_INSTQUEUE_REG_12__1_,
    P1_P3_INSTQUEUE_REG_12__0_, P1_P3_INSTQUEUE_REG_11__7_,
    P1_P3_INSTQUEUE_REG_11__6_, P1_P3_INSTQUEUE_REG_11__5_,
    P1_P3_INSTQUEUE_REG_11__4_, P1_P3_INSTQUEUE_REG_11__3_,
    P1_P3_INSTQUEUE_REG_11__2_, P1_P3_INSTQUEUE_REG_11__1_,
    P1_P3_INSTQUEUE_REG_11__0_, P1_P3_INSTQUEUE_REG_10__7_,
    P1_P3_INSTQUEUE_REG_10__6_, P1_P3_INSTQUEUE_REG_10__5_,
    P1_P3_INSTQUEUE_REG_10__4_, P1_P3_INSTQUEUE_REG_10__3_,
    P1_P3_INSTQUEUE_REG_10__2_, P1_P3_INSTQUEUE_REG_10__1_,
    P1_P3_INSTQUEUE_REG_10__0_, P1_P3_INSTQUEUE_REG_9__7_,
    P1_P3_INSTQUEUE_REG_9__6_, P1_P3_INSTQUEUE_REG_9__5_,
    P1_P3_INSTQUEUE_REG_9__4_, P1_P3_INSTQUEUE_REG_9__3_,
    P1_P3_INSTQUEUE_REG_9__2_, P1_P3_INSTQUEUE_REG_9__1_,
    P1_P3_INSTQUEUE_REG_9__0_, P1_P3_INSTQUEUE_REG_8__7_,
    P1_P3_INSTQUEUE_REG_8__6_, P1_P3_INSTQUEUE_REG_8__5_,
    P1_P3_INSTQUEUE_REG_8__4_, P1_P3_INSTQUEUE_REG_8__3_,
    P1_P3_INSTQUEUE_REG_8__2_, P1_P3_INSTQUEUE_REG_8__1_,
    P1_P3_INSTQUEUE_REG_8__0_, P1_P3_INSTQUEUE_REG_7__7_,
    P1_P3_INSTQUEUE_REG_7__6_, P1_P3_INSTQUEUE_REG_7__5_,
    P1_P3_INSTQUEUE_REG_7__4_, P1_P3_INSTQUEUE_REG_7__3_,
    P1_P3_INSTQUEUE_REG_7__2_, P1_P3_INSTQUEUE_REG_7__1_,
    P1_P3_INSTQUEUE_REG_7__0_, P1_P3_INSTQUEUE_REG_6__7_,
    P1_P3_INSTQUEUE_REG_6__6_, P1_P3_INSTQUEUE_REG_6__5_,
    P1_P3_INSTQUEUE_REG_6__4_, P1_P3_INSTQUEUE_REG_6__3_,
    P1_P3_INSTQUEUE_REG_6__2_, P1_P3_INSTQUEUE_REG_6__1_,
    P1_P3_INSTQUEUE_REG_6__0_, P1_P3_INSTQUEUE_REG_5__7_,
    P1_P3_INSTQUEUE_REG_5__6_, P1_P3_INSTQUEUE_REG_5__5_,
    P1_P3_INSTQUEUE_REG_5__4_, P1_P3_INSTQUEUE_REG_5__3_,
    P1_P3_INSTQUEUE_REG_5__2_, P1_P3_INSTQUEUE_REG_5__1_,
    P1_P3_INSTQUEUE_REG_5__0_, P1_P3_INSTQUEUE_REG_4__7_,
    P1_P3_INSTQUEUE_REG_4__6_, P1_P3_INSTQUEUE_REG_4__5_,
    P1_P3_INSTQUEUE_REG_4__4_, P1_P3_INSTQUEUE_REG_4__3_,
    P1_P3_INSTQUEUE_REG_4__2_, P1_P3_INSTQUEUE_REG_4__1_,
    P1_P3_INSTQUEUE_REG_4__0_, P1_P3_INSTQUEUE_REG_3__7_,
    P1_P3_INSTQUEUE_REG_3__6_, P1_P3_INSTQUEUE_REG_3__5_,
    P1_P3_INSTQUEUE_REG_3__4_, P1_P3_INSTQUEUE_REG_3__3_,
    P1_P3_INSTQUEUE_REG_3__2_, P1_P3_INSTQUEUE_REG_3__1_,
    P1_P3_INSTQUEUE_REG_3__0_, P1_P3_INSTQUEUE_REG_2__7_,
    P1_P3_INSTQUEUE_REG_2__6_, P1_P3_INSTQUEUE_REG_2__5_,
    P1_P3_INSTQUEUE_REG_2__4_, P1_P3_INSTQUEUE_REG_2__3_,
    P1_P3_INSTQUEUE_REG_2__2_, P1_P3_INSTQUEUE_REG_2__1_,
    P1_P3_INSTQUEUE_REG_2__0_, P1_P3_INSTQUEUE_REG_1__7_,
    P1_P3_INSTQUEUE_REG_1__6_, P1_P3_INSTQUEUE_REG_1__5_,
    P1_P3_INSTQUEUE_REG_1__4_, P1_P3_INSTQUEUE_REG_1__3_,
    P1_P3_INSTQUEUE_REG_1__2_, P1_P3_INSTQUEUE_REG_1__1_,
    P1_P3_INSTQUEUE_REG_1__0_, P1_P3_INSTQUEUE_REG_0__7_,
    P1_P3_INSTQUEUE_REG_0__6_, P1_P3_INSTQUEUE_REG_0__5_,
    P1_P3_INSTQUEUE_REG_0__4_, P1_P3_INSTQUEUE_REG_0__3_,
    P1_P3_INSTQUEUE_REG_0__2_, P1_P3_INSTQUEUE_REG_0__1_,
    P1_P3_INSTQUEUE_REG_0__0_, P1_P3_INSTQUEUERD_ADDR_REG_4_,
    P1_P3_INSTQUEUERD_ADDR_REG_3_, P1_P3_INSTQUEUERD_ADDR_REG_2_,
    P1_P3_INSTQUEUERD_ADDR_REG_1_, P1_P3_INSTQUEUERD_ADDR_REG_0_,
    P1_P3_INSTQUEUEWR_ADDR_REG_4_, P1_P3_INSTQUEUEWR_ADDR_REG_3_,
    P1_P3_INSTQUEUEWR_ADDR_REG_2_, P1_P3_INSTQUEUEWR_ADDR_REG_1_,
    P1_P3_INSTQUEUEWR_ADDR_REG_0_, P1_P3_INSTADDRPOINTER_REG_0_,
    P1_P3_INSTADDRPOINTER_REG_1_, P1_P3_INSTADDRPOINTER_REG_2_,
    P1_P3_INSTADDRPOINTER_REG_3_, P1_P3_INSTADDRPOINTER_REG_4_,
    P1_P3_INSTADDRPOINTER_REG_5_, P1_P3_INSTADDRPOINTER_REG_6_,
    P1_P3_INSTADDRPOINTER_REG_7_, P1_P3_INSTADDRPOINTER_REG_8_,
    P1_P3_INSTADDRPOINTER_REG_9_, P1_P3_INSTADDRPOINTER_REG_10_,
    P1_P3_INSTADDRPOINTER_REG_11_, P1_P3_INSTADDRPOINTER_REG_12_,
    P1_P3_INSTADDRPOINTER_REG_13_, P1_P3_INSTADDRPOINTER_REG_14_,
    P1_P3_INSTADDRPOINTER_REG_15_, P1_P3_INSTADDRPOINTER_REG_16_,
    P1_P3_INSTADDRPOINTER_REG_17_, P1_P3_INSTADDRPOINTER_REG_18_,
    P1_P3_INSTADDRPOINTER_REG_19_, P1_P3_INSTADDRPOINTER_REG_20_,
    P1_P3_INSTADDRPOINTER_REG_21_, P1_P3_INSTADDRPOINTER_REG_22_,
    P1_P3_INSTADDRPOINTER_REG_23_, P1_P3_INSTADDRPOINTER_REG_24_,
    P1_P3_INSTADDRPOINTER_REG_25_, P1_P3_INSTADDRPOINTER_REG_26_,
    P1_P3_INSTADDRPOINTER_REG_27_, P1_P3_INSTADDRPOINTER_REG_28_,
    P1_P3_INSTADDRPOINTER_REG_29_, P1_P3_INSTADDRPOINTER_REG_30_,
    P1_P3_INSTADDRPOINTER_REG_31_, P1_P3_PHYADDRPOINTER_REG_0_,
    P1_P3_PHYADDRPOINTER_REG_1_, P1_P3_PHYADDRPOINTER_REG_2_,
    P1_P3_PHYADDRPOINTER_REG_3_, P1_P3_PHYADDRPOINTER_REG_4_,
    P1_P3_PHYADDRPOINTER_REG_5_, P1_P3_PHYADDRPOINTER_REG_6_,
    P1_P3_PHYADDRPOINTER_REG_7_, P1_P3_PHYADDRPOINTER_REG_8_,
    P1_P3_PHYADDRPOINTER_REG_9_, P1_P3_PHYADDRPOINTER_REG_10_,
    P1_P3_PHYADDRPOINTER_REG_11_, P1_P3_PHYADDRPOINTER_REG_12_,
    P1_P3_PHYADDRPOINTER_REG_13_, P1_P3_PHYADDRPOINTER_REG_14_,
    P1_P3_PHYADDRPOINTER_REG_15_, P1_P3_PHYADDRPOINTER_REG_16_,
    P1_P3_PHYADDRPOINTER_REG_17_, P1_P3_PHYADDRPOINTER_REG_18_,
    P1_P3_PHYADDRPOINTER_REG_19_, P1_P3_PHYADDRPOINTER_REG_20_,
    P1_P3_PHYADDRPOINTER_REG_21_, P1_P3_PHYADDRPOINTER_REG_22_,
    P1_P3_PHYADDRPOINTER_REG_23_, P1_P3_PHYADDRPOINTER_REG_24_,
    P1_P3_PHYADDRPOINTER_REG_25_, P1_P3_PHYADDRPOINTER_REG_26_,
    P1_P3_PHYADDRPOINTER_REG_27_, P1_P3_PHYADDRPOINTER_REG_28_,
    P1_P3_PHYADDRPOINTER_REG_29_, P1_P3_PHYADDRPOINTER_REG_30_,
    P1_P3_PHYADDRPOINTER_REG_31_, P1_P3_LWORD_REG_15_, P1_P3_LWORD_REG_14_,
    P1_P3_LWORD_REG_13_, P1_P3_LWORD_REG_12_, P1_P3_LWORD_REG_11_,
    P1_P3_LWORD_REG_10_, P1_P3_LWORD_REG_9_, P1_P3_LWORD_REG_8_,
    P1_P3_LWORD_REG_7_, P1_P3_LWORD_REG_6_, P1_P3_LWORD_REG_5_,
    P1_P3_LWORD_REG_4_, P1_P3_LWORD_REG_3_, P1_P3_LWORD_REG_2_,
    P1_P3_LWORD_REG_1_, P1_P3_LWORD_REG_0_, P1_P3_UWORD_REG_14_,
    P1_P3_UWORD_REG_13_, P1_P3_UWORD_REG_12_, P1_P3_UWORD_REG_11_,
    P1_P3_UWORD_REG_10_, P1_P3_UWORD_REG_9_, P1_P3_UWORD_REG_8_,
    P1_P3_UWORD_REG_7_, P1_P3_UWORD_REG_6_, P1_P3_UWORD_REG_5_,
    P1_P3_UWORD_REG_4_, P1_P3_UWORD_REG_3_, P1_P3_UWORD_REG_2_,
    P1_P3_UWORD_REG_1_, P1_P3_UWORD_REG_0_, P1_P3_DATAO_REG_0_,
    P1_P3_DATAO_REG_1_, P1_P3_DATAO_REG_2_, P1_P3_DATAO_REG_3_,
    P1_P3_DATAO_REG_4_, P1_P3_DATAO_REG_5_, P1_P3_DATAO_REG_6_,
    P1_P3_DATAO_REG_7_, P1_P3_DATAO_REG_8_, P1_P3_DATAO_REG_9_,
    P1_P3_DATAO_REG_10_, P1_P3_DATAO_REG_11_, P1_P3_DATAO_REG_12_,
    P1_P3_DATAO_REG_13_, P1_P3_DATAO_REG_14_, P1_P3_DATAO_REG_15_,
    P1_P3_DATAO_REG_16_, P1_P3_DATAO_REG_17_, P1_P3_DATAO_REG_18_,
    P1_P3_DATAO_REG_19_, P1_P3_DATAO_REG_20_, P1_P3_DATAO_REG_21_,
    P1_P3_DATAO_REG_22_, P1_P3_DATAO_REG_23_, P1_P3_DATAO_REG_24_,
    P1_P3_DATAO_REG_25_, P1_P3_DATAO_REG_26_, P1_P3_DATAO_REG_27_,
    P1_P3_DATAO_REG_28_, P1_P3_DATAO_REG_29_, P1_P3_DATAO_REG_30_,
    P1_P3_DATAO_REG_31_, P1_P3_EAX_REG_0_, P1_P3_EAX_REG_1_,
    P1_P3_EAX_REG_2_, P1_P3_EAX_REG_3_, P1_P3_EAX_REG_4_, P1_P3_EAX_REG_5_,
    P1_P3_EAX_REG_6_, P1_P3_EAX_REG_7_, P1_P3_EAX_REG_8_, P1_P3_EAX_REG_9_,
    P1_P3_EAX_REG_10_, P1_P3_EAX_REG_11_, P1_P3_EAX_REG_12_,
    P1_P3_EAX_REG_13_, P1_P3_EAX_REG_14_, P1_P3_EAX_REG_15_,
    P1_P3_EAX_REG_16_, P1_P3_EAX_REG_17_, P1_P3_EAX_REG_18_,
    P1_P3_EAX_REG_19_, P1_P3_EAX_REG_20_, P1_P3_EAX_REG_21_,
    P1_P3_EAX_REG_22_, P1_P3_EAX_REG_23_, P1_P3_EAX_REG_24_,
    P1_P3_EAX_REG_25_, P1_P3_EAX_REG_26_, P1_P3_EAX_REG_27_,
    P1_P3_EAX_REG_28_, P1_P3_EAX_REG_29_, P1_P3_EAX_REG_30_,
    P1_P3_EAX_REG_31_, P1_P3_EBX_REG_0_, P1_P3_EBX_REG_1_,
    P1_P3_EBX_REG_2_, P1_P3_EBX_REG_3_, P1_P3_EBX_REG_4_, P1_P3_EBX_REG_5_,
    P1_P3_EBX_REG_6_, P1_P3_EBX_REG_7_, P1_P3_EBX_REG_8_, P1_P3_EBX_REG_9_,
    P1_P3_EBX_REG_10_, P1_P3_EBX_REG_11_, P1_P3_EBX_REG_12_,
    P1_P3_EBX_REG_13_, P1_P3_EBX_REG_14_, P1_P3_EBX_REG_15_,
    P1_P3_EBX_REG_16_, P1_P3_EBX_REG_17_, P1_P3_EBX_REG_18_,
    P1_P3_EBX_REG_19_, P1_P3_EBX_REG_20_, P1_P3_EBX_REG_21_,
    P1_P3_EBX_REG_22_, P1_P3_EBX_REG_23_, P1_P3_EBX_REG_24_,
    P1_P3_EBX_REG_25_, P1_P3_EBX_REG_26_, P1_P3_EBX_REG_27_,
    P1_P3_EBX_REG_28_, P1_P3_EBX_REG_29_, P1_P3_EBX_REG_30_,
    P1_P3_EBX_REG_31_, P1_P3_REIP_REG_0_, P1_P3_REIP_REG_1_,
    P1_P3_REIP_REG_2_, P1_P3_REIP_REG_3_, P1_P3_REIP_REG_4_,
    P1_P3_REIP_REG_5_, P1_P3_REIP_REG_6_, P1_P3_REIP_REG_7_,
    P1_P3_REIP_REG_8_, P1_P3_REIP_REG_9_, P1_P3_REIP_REG_10_,
    P1_P3_REIP_REG_11_, P1_P3_REIP_REG_12_, P1_P3_REIP_REG_13_,
    P1_P3_REIP_REG_14_, P1_P3_REIP_REG_15_, P1_P3_REIP_REG_16_,
    P1_P3_REIP_REG_17_, P1_P3_REIP_REG_18_, P1_P3_REIP_REG_19_,
    P1_P3_REIP_REG_20_, P1_P3_REIP_REG_21_, P1_P3_REIP_REG_22_,
    P1_P3_REIP_REG_23_, P1_P3_REIP_REG_24_, P1_P3_REIP_REG_25_,
    P1_P3_REIP_REG_26_, P1_P3_REIP_REG_27_, P1_P3_REIP_REG_28_,
    P1_P3_REIP_REG_29_, P1_P3_REIP_REG_30_, P1_P3_REIP_REG_31_,
    P1_P3_BYTEENABLE_REG_3_, P1_P3_BYTEENABLE_REG_2_,
    P1_P3_BYTEENABLE_REG_1_, P1_P3_BYTEENABLE_REG_0_, P1_P3_W_R_N_REG,
    P1_P3_FLUSH_REG, P1_P3_MORE_REG, P1_P3_STATEBS16_REG,
    P1_P3_REQUESTPENDING_REG, P1_P3_D_C_N_REG, P1_P3_M_IO_N_REG,
    P1_P3_CODEFETCH_REG, P1_P3_ADS_N_REG, P1_P3_READREQUEST_REG,
    P1_P3_MEMORYFETCH_REG, P1_P2_BE_N_REG_3_, P1_P2_BE_N_REG_2_,
    P1_P2_BE_N_REG_1_, P1_P2_BE_N_REG_0_, P1_P2_ADDRESS_REG_29_,
    P1_P2_ADDRESS_REG_28_, P1_P2_ADDRESS_REG_27_, P1_P2_ADDRESS_REG_26_,
    P1_P2_ADDRESS_REG_25_, P1_P2_ADDRESS_REG_24_, P1_P2_ADDRESS_REG_23_,
    P1_P2_ADDRESS_REG_22_, P1_P2_ADDRESS_REG_21_, P1_P2_ADDRESS_REG_20_,
    P1_P2_ADDRESS_REG_19_, P1_P2_ADDRESS_REG_18_, P1_P2_ADDRESS_REG_17_,
    P1_P2_ADDRESS_REG_16_, P1_P2_ADDRESS_REG_15_, P1_P2_ADDRESS_REG_14_,
    P1_P2_ADDRESS_REG_13_, P1_P2_ADDRESS_REG_12_, P1_P2_ADDRESS_REG_11_,
    P1_P2_ADDRESS_REG_10_, P1_P2_ADDRESS_REG_9_, P1_P2_ADDRESS_REG_8_,
    P1_P2_ADDRESS_REG_7_, P1_P2_ADDRESS_REG_6_, P1_P2_ADDRESS_REG_5_,
    P1_P2_ADDRESS_REG_4_, P1_P2_ADDRESS_REG_3_, P1_P2_ADDRESS_REG_2_,
    P1_P2_ADDRESS_REG_1_, P1_P2_ADDRESS_REG_0_, P1_P2_STATE_REG_2_,
    P1_P2_STATE_REG_1_, P1_P2_STATE_REG_0_, P1_P2_DATAWIDTH_REG_0_,
    P1_P2_DATAWIDTH_REG_1_, P1_P2_DATAWIDTH_REG_2_, P1_P2_DATAWIDTH_REG_3_,
    P1_P2_DATAWIDTH_REG_4_, P1_P2_DATAWIDTH_REG_5_, P1_P2_DATAWIDTH_REG_6_,
    P1_P2_DATAWIDTH_REG_7_, P1_P2_DATAWIDTH_REG_8_, P1_P2_DATAWIDTH_REG_9_,
    P1_P2_DATAWIDTH_REG_10_, P1_P2_DATAWIDTH_REG_11_,
    P1_P2_DATAWIDTH_REG_12_, P1_P2_DATAWIDTH_REG_13_,
    P1_P2_DATAWIDTH_REG_14_, P1_P2_DATAWIDTH_REG_15_,
    P1_P2_DATAWIDTH_REG_16_, P1_P2_DATAWIDTH_REG_17_,
    P1_P2_DATAWIDTH_REG_18_, P1_P2_DATAWIDTH_REG_19_,
    P1_P2_DATAWIDTH_REG_20_, P1_P2_DATAWIDTH_REG_21_,
    P1_P2_DATAWIDTH_REG_22_, P1_P2_DATAWIDTH_REG_23_,
    P1_P2_DATAWIDTH_REG_24_, P1_P2_DATAWIDTH_REG_25_,
    P1_P2_DATAWIDTH_REG_26_, P1_P2_DATAWIDTH_REG_27_,
    P1_P2_DATAWIDTH_REG_28_, P1_P2_DATAWIDTH_REG_29_,
    P1_P2_DATAWIDTH_REG_30_, P1_P2_DATAWIDTH_REG_31_, P1_P2_STATE2_REG_3_,
    P1_P2_STATE2_REG_2_, P1_P2_STATE2_REG_1_, P1_P2_STATE2_REG_0_,
    P1_P2_INSTQUEUE_REG_15__7_, P1_P2_INSTQUEUE_REG_15__6_,
    P1_P2_INSTQUEUE_REG_15__5_, P1_P2_INSTQUEUE_REG_15__4_,
    P1_P2_INSTQUEUE_REG_15__3_, P1_P2_INSTQUEUE_REG_15__2_,
    P1_P2_INSTQUEUE_REG_15__1_, P1_P2_INSTQUEUE_REG_15__0_,
    P1_P2_INSTQUEUE_REG_14__7_, P1_P2_INSTQUEUE_REG_14__6_,
    P1_P2_INSTQUEUE_REG_14__5_, P1_P2_INSTQUEUE_REG_14__4_,
    P1_P2_INSTQUEUE_REG_14__3_, P1_P2_INSTQUEUE_REG_14__2_,
    P1_P2_INSTQUEUE_REG_14__1_, P1_P2_INSTQUEUE_REG_14__0_,
    P1_P2_INSTQUEUE_REG_13__7_, P1_P2_INSTQUEUE_REG_13__6_,
    P1_P2_INSTQUEUE_REG_13__5_, P1_P2_INSTQUEUE_REG_13__4_,
    P1_P2_INSTQUEUE_REG_13__3_, P1_P2_INSTQUEUE_REG_13__2_,
    P1_P2_INSTQUEUE_REG_13__1_, P1_P2_INSTQUEUE_REG_13__0_,
    P1_P2_INSTQUEUE_REG_12__7_, P1_P2_INSTQUEUE_REG_12__6_,
    P1_P2_INSTQUEUE_REG_12__5_, P1_P2_INSTQUEUE_REG_12__4_,
    P1_P2_INSTQUEUE_REG_12__3_, P1_P2_INSTQUEUE_REG_12__2_,
    P1_P2_INSTQUEUE_REG_12__1_, P1_P2_INSTQUEUE_REG_12__0_,
    P1_P2_INSTQUEUE_REG_11__7_, P1_P2_INSTQUEUE_REG_11__6_,
    P1_P2_INSTQUEUE_REG_11__5_, P1_P2_INSTQUEUE_REG_11__4_,
    P1_P2_INSTQUEUE_REG_11__3_, P1_P2_INSTQUEUE_REG_11__2_,
    P1_P2_INSTQUEUE_REG_11__1_, P1_P2_INSTQUEUE_REG_11__0_,
    P1_P2_INSTQUEUE_REG_10__7_, P1_P2_INSTQUEUE_REG_10__6_,
    P1_P2_INSTQUEUE_REG_10__5_, P1_P2_INSTQUEUE_REG_10__4_,
    P1_P2_INSTQUEUE_REG_10__3_, P1_P2_INSTQUEUE_REG_10__2_,
    P1_P2_INSTQUEUE_REG_10__1_, P1_P2_INSTQUEUE_REG_10__0_,
    P1_P2_INSTQUEUE_REG_9__7_, P1_P2_INSTQUEUE_REG_9__6_,
    P1_P2_INSTQUEUE_REG_9__5_, P1_P2_INSTQUEUE_REG_9__4_,
    P1_P2_INSTQUEUE_REG_9__3_, P1_P2_INSTQUEUE_REG_9__2_,
    P1_P2_INSTQUEUE_REG_9__1_, P1_P2_INSTQUEUE_REG_9__0_,
    P1_P2_INSTQUEUE_REG_8__7_, P1_P2_INSTQUEUE_REG_8__6_,
    P1_P2_INSTQUEUE_REG_8__5_, P1_P2_INSTQUEUE_REG_8__4_,
    P1_P2_INSTQUEUE_REG_8__3_, P1_P2_INSTQUEUE_REG_8__2_,
    P1_P2_INSTQUEUE_REG_8__1_, P1_P2_INSTQUEUE_REG_8__0_,
    P1_P2_INSTQUEUE_REG_7__7_, P1_P2_INSTQUEUE_REG_7__6_,
    P1_P2_INSTQUEUE_REG_7__5_, P1_P2_INSTQUEUE_REG_7__4_,
    P1_P2_INSTQUEUE_REG_7__3_, P1_P2_INSTQUEUE_REG_7__2_,
    P1_P2_INSTQUEUE_REG_7__1_, P1_P2_INSTQUEUE_REG_7__0_,
    P1_P2_INSTQUEUE_REG_6__7_, P1_P2_INSTQUEUE_REG_6__6_,
    P1_P2_INSTQUEUE_REG_6__5_, P1_P2_INSTQUEUE_REG_6__4_,
    P1_P2_INSTQUEUE_REG_6__3_, P1_P2_INSTQUEUE_REG_6__2_,
    P1_P2_INSTQUEUE_REG_6__1_, P1_P2_INSTQUEUE_REG_6__0_,
    P1_P2_INSTQUEUE_REG_5__7_, P1_P2_INSTQUEUE_REG_5__6_,
    P1_P2_INSTQUEUE_REG_5__5_, P1_P2_INSTQUEUE_REG_5__4_,
    P1_P2_INSTQUEUE_REG_5__3_, P1_P2_INSTQUEUE_REG_5__2_,
    P1_P2_INSTQUEUE_REG_5__1_, P1_P2_INSTQUEUE_REG_5__0_,
    P1_P2_INSTQUEUE_REG_4__7_, P1_P2_INSTQUEUE_REG_4__6_,
    P1_P2_INSTQUEUE_REG_4__5_, P1_P2_INSTQUEUE_REG_4__4_,
    P1_P2_INSTQUEUE_REG_4__3_, P1_P2_INSTQUEUE_REG_4__2_,
    P1_P2_INSTQUEUE_REG_4__1_, P1_P2_INSTQUEUE_REG_4__0_,
    P1_P2_INSTQUEUE_REG_3__7_, P1_P2_INSTQUEUE_REG_3__6_,
    P1_P2_INSTQUEUE_REG_3__5_, P1_P2_INSTQUEUE_REG_3__4_,
    P1_P2_INSTQUEUE_REG_3__3_, P1_P2_INSTQUEUE_REG_3__2_,
    P1_P2_INSTQUEUE_REG_3__1_, P1_P2_INSTQUEUE_REG_3__0_,
    P1_P2_INSTQUEUE_REG_2__7_, P1_P2_INSTQUEUE_REG_2__6_,
    P1_P2_INSTQUEUE_REG_2__5_, P1_P2_INSTQUEUE_REG_2__4_,
    P1_P2_INSTQUEUE_REG_2__3_, P1_P2_INSTQUEUE_REG_2__2_,
    P1_P2_INSTQUEUE_REG_2__1_, P1_P2_INSTQUEUE_REG_2__0_,
    P1_P2_INSTQUEUE_REG_1__7_, P1_P2_INSTQUEUE_REG_1__6_,
    P1_P2_INSTQUEUE_REG_1__5_, P1_P2_INSTQUEUE_REG_1__4_,
    P1_P2_INSTQUEUE_REG_1__3_, P1_P2_INSTQUEUE_REG_1__2_,
    P1_P2_INSTQUEUE_REG_1__1_, P1_P2_INSTQUEUE_REG_1__0_,
    P1_P2_INSTQUEUE_REG_0__7_, P1_P2_INSTQUEUE_REG_0__6_,
    P1_P2_INSTQUEUE_REG_0__5_, P1_P2_INSTQUEUE_REG_0__4_,
    P1_P2_INSTQUEUE_REG_0__3_, P1_P2_INSTQUEUE_REG_0__2_,
    P1_P2_INSTQUEUE_REG_0__1_, P1_P2_INSTQUEUE_REG_0__0_,
    P1_P2_INSTQUEUERD_ADDR_REG_4_, P1_P2_INSTQUEUERD_ADDR_REG_3_,
    P1_P2_INSTQUEUERD_ADDR_REG_2_, P1_P2_INSTQUEUERD_ADDR_REG_1_,
    P1_P2_INSTQUEUERD_ADDR_REG_0_, P1_P2_INSTQUEUEWR_ADDR_REG_4_,
    P1_P2_INSTQUEUEWR_ADDR_REG_3_, P1_P2_INSTQUEUEWR_ADDR_REG_2_,
    P1_P2_INSTQUEUEWR_ADDR_REG_1_, P1_P2_INSTQUEUEWR_ADDR_REG_0_,
    P1_P2_INSTADDRPOINTER_REG_0_, P1_P2_INSTADDRPOINTER_REG_1_,
    P1_P2_INSTADDRPOINTER_REG_2_, P1_P2_INSTADDRPOINTER_REG_3_,
    P1_P2_INSTADDRPOINTER_REG_4_, P1_P2_INSTADDRPOINTER_REG_5_,
    P1_P2_INSTADDRPOINTER_REG_6_, P1_P2_INSTADDRPOINTER_REG_7_,
    P1_P2_INSTADDRPOINTER_REG_8_, P1_P2_INSTADDRPOINTER_REG_9_,
    P1_P2_INSTADDRPOINTER_REG_10_, P1_P2_INSTADDRPOINTER_REG_11_,
    P1_P2_INSTADDRPOINTER_REG_12_, P1_P2_INSTADDRPOINTER_REG_13_,
    P1_P2_INSTADDRPOINTER_REG_14_, P1_P2_INSTADDRPOINTER_REG_15_,
    P1_P2_INSTADDRPOINTER_REG_16_, P1_P2_INSTADDRPOINTER_REG_17_,
    P1_P2_INSTADDRPOINTER_REG_18_, P1_P2_INSTADDRPOINTER_REG_19_,
    P1_P2_INSTADDRPOINTER_REG_20_, P1_P2_INSTADDRPOINTER_REG_21_,
    P1_P2_INSTADDRPOINTER_REG_22_, P1_P2_INSTADDRPOINTER_REG_23_,
    P1_P2_INSTADDRPOINTER_REG_24_, P1_P2_INSTADDRPOINTER_REG_25_,
    P1_P2_INSTADDRPOINTER_REG_26_, P1_P2_INSTADDRPOINTER_REG_27_,
    P1_P2_INSTADDRPOINTER_REG_28_, P1_P2_INSTADDRPOINTER_REG_29_,
    P1_P2_INSTADDRPOINTER_REG_30_, P1_P2_INSTADDRPOINTER_REG_31_,
    P1_P2_PHYADDRPOINTER_REG_0_, P1_P2_PHYADDRPOINTER_REG_1_,
    P1_P2_PHYADDRPOINTER_REG_2_, P1_P2_PHYADDRPOINTER_REG_3_,
    P1_P2_PHYADDRPOINTER_REG_4_, P1_P2_PHYADDRPOINTER_REG_5_,
    P1_P2_PHYADDRPOINTER_REG_6_, P1_P2_PHYADDRPOINTER_REG_7_,
    P1_P2_PHYADDRPOINTER_REG_8_, P1_P2_PHYADDRPOINTER_REG_9_,
    P1_P2_PHYADDRPOINTER_REG_10_, P1_P2_PHYADDRPOINTER_REG_11_,
    P1_P2_PHYADDRPOINTER_REG_12_, P1_P2_PHYADDRPOINTER_REG_13_,
    P1_P2_PHYADDRPOINTER_REG_14_, P1_P2_PHYADDRPOINTER_REG_15_,
    P1_P2_PHYADDRPOINTER_REG_16_, P1_P2_PHYADDRPOINTER_REG_17_,
    P1_P2_PHYADDRPOINTER_REG_18_, P1_P2_PHYADDRPOINTER_REG_19_,
    P1_P2_PHYADDRPOINTER_REG_20_, P1_P2_PHYADDRPOINTER_REG_21_,
    P1_P2_PHYADDRPOINTER_REG_22_, P1_P2_PHYADDRPOINTER_REG_23_,
    P1_P2_PHYADDRPOINTER_REG_24_, P1_P2_PHYADDRPOINTER_REG_25_,
    P1_P2_PHYADDRPOINTER_REG_26_, P1_P2_PHYADDRPOINTER_REG_27_,
    P1_P2_PHYADDRPOINTER_REG_28_, P1_P2_PHYADDRPOINTER_REG_29_,
    P1_P2_PHYADDRPOINTER_REG_30_, P1_P2_PHYADDRPOINTER_REG_31_,
    P1_P2_LWORD_REG_15_, P1_P2_LWORD_REG_14_, P1_P2_LWORD_REG_13_,
    P1_P2_LWORD_REG_12_, P1_P2_LWORD_REG_11_, P1_P2_LWORD_REG_10_,
    P1_P2_LWORD_REG_9_, P1_P2_LWORD_REG_8_, P1_P2_LWORD_REG_7_,
    P1_P2_LWORD_REG_6_, P1_P2_LWORD_REG_5_, P1_P2_LWORD_REG_4_,
    P1_P2_LWORD_REG_3_, P1_P2_LWORD_REG_2_, P1_P2_LWORD_REG_1_,
    P1_P2_LWORD_REG_0_, P1_P2_UWORD_REG_14_, P1_P2_UWORD_REG_13_,
    P1_P2_UWORD_REG_12_, P1_P2_UWORD_REG_11_, P1_P2_UWORD_REG_10_,
    P1_P2_UWORD_REG_9_, P1_P2_UWORD_REG_8_, P1_P2_UWORD_REG_7_,
    P1_P2_UWORD_REG_6_, P1_P2_UWORD_REG_5_, P1_P2_UWORD_REG_4_,
    P1_P2_UWORD_REG_3_, P1_P2_UWORD_REG_2_, P1_P2_UWORD_REG_1_,
    P1_P2_UWORD_REG_0_, P1_P2_DATAO_REG_0_, P1_P2_DATAO_REG_1_,
    P1_P2_DATAO_REG_2_, P1_P2_DATAO_REG_3_, P1_P2_DATAO_REG_4_,
    P1_P2_DATAO_REG_5_, P1_P2_DATAO_REG_6_, P1_P2_DATAO_REG_7_,
    P1_P2_DATAO_REG_8_, P1_P2_DATAO_REG_9_, P1_P2_DATAO_REG_10_,
    P1_P2_DATAO_REG_11_, P1_P2_DATAO_REG_12_, P1_P2_DATAO_REG_13_,
    P1_P2_DATAO_REG_14_, P1_P2_DATAO_REG_15_, P1_P2_DATAO_REG_16_,
    P1_P2_DATAO_REG_17_, P1_P2_DATAO_REG_18_, P1_P2_DATAO_REG_19_,
    P1_P2_DATAO_REG_20_, P1_P2_DATAO_REG_21_, P1_P2_DATAO_REG_22_,
    P1_P2_DATAO_REG_23_, P1_P2_DATAO_REG_24_, P1_P2_DATAO_REG_25_,
    P1_P2_DATAO_REG_26_, P1_P2_DATAO_REG_27_, P1_P2_DATAO_REG_28_,
    P1_P2_DATAO_REG_29_, P1_P2_DATAO_REG_30_, P1_P2_DATAO_REG_31_,
    P1_P2_EAX_REG_0_, P1_P2_EAX_REG_1_, P1_P2_EAX_REG_2_, P1_P2_EAX_REG_3_,
    P1_P2_EAX_REG_4_, P1_P2_EAX_REG_5_, P1_P2_EAX_REG_6_, P1_P2_EAX_REG_7_,
    P1_P2_EAX_REG_8_, P1_P2_EAX_REG_9_, P1_P2_EAX_REG_10_,
    P1_P2_EAX_REG_11_, P1_P2_EAX_REG_12_, P1_P2_EAX_REG_13_,
    P1_P2_EAX_REG_14_, P1_P2_EAX_REG_15_, P1_P2_EAX_REG_16_,
    P1_P2_EAX_REG_17_, P1_P2_EAX_REG_18_, P1_P2_EAX_REG_19_,
    P1_P2_EAX_REG_20_, P1_P2_EAX_REG_21_, P1_P2_EAX_REG_22_,
    P1_P2_EAX_REG_23_, P1_P2_EAX_REG_24_, P1_P2_EAX_REG_25_,
    P1_P2_EAX_REG_26_, P1_P2_EAX_REG_27_, P1_P2_EAX_REG_28_,
    P1_P2_EAX_REG_29_, P1_P2_EAX_REG_30_, P1_P2_EAX_REG_31_,
    P1_P2_EBX_REG_0_, P1_P2_EBX_REG_1_, P1_P2_EBX_REG_2_, P1_P2_EBX_REG_3_,
    P1_P2_EBX_REG_4_, P1_P2_EBX_REG_5_, P1_P2_EBX_REG_6_, P1_P2_EBX_REG_7_,
    P1_P2_EBX_REG_8_, P1_P2_EBX_REG_9_, P1_P2_EBX_REG_10_,
    P1_P2_EBX_REG_11_, P1_P2_EBX_REG_12_, P1_P2_EBX_REG_13_,
    P1_P2_EBX_REG_14_, P1_P2_EBX_REG_15_, P1_P2_EBX_REG_16_,
    P1_P2_EBX_REG_17_, P1_P2_EBX_REG_18_, P1_P2_EBX_REG_19_,
    P1_P2_EBX_REG_20_, P1_P2_EBX_REG_21_, P1_P2_EBX_REG_22_,
    P1_P2_EBX_REG_23_, P1_P2_EBX_REG_24_, P1_P2_EBX_REG_25_,
    P1_P2_EBX_REG_26_, P1_P2_EBX_REG_27_, P1_P2_EBX_REG_28_,
    P1_P2_EBX_REG_29_, P1_P2_EBX_REG_30_, P1_P2_EBX_REG_31_,
    P1_P2_REIP_REG_0_, P1_P2_REIP_REG_1_, P1_P2_REIP_REG_2_,
    P1_P2_REIP_REG_3_, P1_P2_REIP_REG_4_, P1_P2_REIP_REG_5_,
    P1_P2_REIP_REG_6_, P1_P2_REIP_REG_7_, P1_P2_REIP_REG_8_,
    P1_P2_REIP_REG_9_, P1_P2_REIP_REG_10_, P1_P2_REIP_REG_11_,
    P1_P2_REIP_REG_12_, P1_P2_REIP_REG_13_, P1_P2_REIP_REG_14_,
    P1_P2_REIP_REG_15_, P1_P2_REIP_REG_16_, P1_P2_REIP_REG_17_,
    P1_P2_REIP_REG_18_, P1_P2_REIP_REG_19_, P1_P2_REIP_REG_20_,
    P1_P2_REIP_REG_21_, P1_P2_REIP_REG_22_, P1_P2_REIP_REG_23_,
    P1_P2_REIP_REG_24_, P1_P2_REIP_REG_25_, P1_P2_REIP_REG_26_,
    P1_P2_REIP_REG_27_, P1_P2_REIP_REG_28_, P1_P2_REIP_REG_29_,
    P1_P2_REIP_REG_30_, P1_P2_REIP_REG_31_, P1_P2_BYTEENABLE_REG_3_,
    P1_P2_BYTEENABLE_REG_2_, P1_P2_BYTEENABLE_REG_1_,
    P1_P2_BYTEENABLE_REG_0_, P1_P2_W_R_N_REG, P1_P2_FLUSH_REG,
    P1_P2_MORE_REG, P1_P2_STATEBS16_REG, P1_P2_REQUESTPENDING_REG,
    P1_P2_D_C_N_REG, P1_P2_M_IO_N_REG, P1_P2_CODEFETCH_REG,
    P1_P2_ADS_N_REG, P1_P2_READREQUEST_REG, P1_P2_MEMORYFETCH_REG,
    P1_P1_BE_N_REG_3_, P1_P1_BE_N_REG_2_, P1_P1_BE_N_REG_1_,
    P1_P1_BE_N_REG_0_, P1_P1_ADDRESS_REG_29_, P1_P1_ADDRESS_REG_28_,
    P1_P1_ADDRESS_REG_27_, P1_P1_ADDRESS_REG_26_, P1_P1_ADDRESS_REG_25_,
    P1_P1_ADDRESS_REG_24_, P1_P1_ADDRESS_REG_23_, P1_P1_ADDRESS_REG_22_,
    P1_P1_ADDRESS_REG_21_, P1_P1_ADDRESS_REG_20_, P1_P1_ADDRESS_REG_19_,
    P1_P1_ADDRESS_REG_18_, P1_P1_ADDRESS_REG_17_, P1_P1_ADDRESS_REG_16_,
    P1_P1_ADDRESS_REG_15_, P1_P1_ADDRESS_REG_14_, P1_P1_ADDRESS_REG_13_,
    P1_P1_ADDRESS_REG_12_, P1_P1_ADDRESS_REG_11_, P1_P1_ADDRESS_REG_10_,
    P1_P1_ADDRESS_REG_9_, P1_P1_ADDRESS_REG_8_, P1_P1_ADDRESS_REG_7_,
    P1_P1_ADDRESS_REG_6_, P1_P1_ADDRESS_REG_5_, P1_P1_ADDRESS_REG_4_,
    P1_P1_ADDRESS_REG_3_, P1_P1_ADDRESS_REG_2_, P1_P1_ADDRESS_REG_1_,
    P1_P1_ADDRESS_REG_0_, P1_P1_STATE_REG_2_, P1_P1_STATE_REG_1_,
    P1_P1_STATE_REG_0_, P1_P1_DATAWIDTH_REG_0_, P1_P1_DATAWIDTH_REG_1_,
    P1_P1_DATAWIDTH_REG_2_, P1_P1_DATAWIDTH_REG_3_, P1_P1_DATAWIDTH_REG_4_,
    P1_P1_DATAWIDTH_REG_5_, P1_P1_DATAWIDTH_REG_6_, P1_P1_DATAWIDTH_REG_7_,
    P1_P1_DATAWIDTH_REG_8_, P1_P1_DATAWIDTH_REG_9_,
    P1_P1_DATAWIDTH_REG_10_, P1_P1_DATAWIDTH_REG_11_,
    P1_P1_DATAWIDTH_REG_12_, P1_P1_DATAWIDTH_REG_13_,
    P1_P1_DATAWIDTH_REG_14_, P1_P1_DATAWIDTH_REG_15_,
    P1_P1_DATAWIDTH_REG_16_, P1_P1_DATAWIDTH_REG_17_,
    P1_P1_DATAWIDTH_REG_18_, P1_P1_DATAWIDTH_REG_19_,
    P1_P1_DATAWIDTH_REG_20_, P1_P1_DATAWIDTH_REG_21_,
    P1_P1_DATAWIDTH_REG_22_, P1_P1_DATAWIDTH_REG_23_,
    P1_P1_DATAWIDTH_REG_24_, P1_P1_DATAWIDTH_REG_25_,
    P1_P1_DATAWIDTH_REG_26_, P1_P1_DATAWIDTH_REG_27_,
    P1_P1_DATAWIDTH_REG_28_, P1_P1_DATAWIDTH_REG_29_,
    P1_P1_DATAWIDTH_REG_30_, P1_P1_DATAWIDTH_REG_31_, P1_P1_STATE2_REG_3_,
    P1_P1_STATE2_REG_2_, P1_P1_STATE2_REG_1_, P1_P1_STATE2_REG_0_,
    P1_P1_INSTQUEUE_REG_15__7_, P1_P1_INSTQUEUE_REG_15__6_,
    P1_P1_INSTQUEUE_REG_15__5_, P1_P1_INSTQUEUE_REG_15__4_,
    P1_P1_INSTQUEUE_REG_15__3_, P1_P1_INSTQUEUE_REG_15__2_,
    P1_P1_INSTQUEUE_REG_15__1_, P1_P1_INSTQUEUE_REG_15__0_,
    P1_P1_INSTQUEUE_REG_14__7_, P1_P1_INSTQUEUE_REG_14__6_,
    P1_P1_INSTQUEUE_REG_14__5_, P1_P1_INSTQUEUE_REG_14__4_,
    P1_P1_INSTQUEUE_REG_14__3_, P1_P1_INSTQUEUE_REG_14__2_,
    P1_P1_INSTQUEUE_REG_14__1_, P1_P1_INSTQUEUE_REG_14__0_,
    P1_P1_INSTQUEUE_REG_13__7_, P1_P1_INSTQUEUE_REG_13__6_,
    P1_P1_INSTQUEUE_REG_13__5_, P1_P1_INSTQUEUE_REG_13__4_,
    P1_P1_INSTQUEUE_REG_13__3_, P1_P1_INSTQUEUE_REG_13__2_,
    P1_P1_INSTQUEUE_REG_13__1_, P1_P1_INSTQUEUE_REG_13__0_,
    P1_P1_INSTQUEUE_REG_12__7_, P1_P1_INSTQUEUE_REG_12__6_,
    P1_P1_INSTQUEUE_REG_12__5_, P1_P1_INSTQUEUE_REG_12__4_,
    P1_P1_INSTQUEUE_REG_12__3_, P1_P1_INSTQUEUE_REG_12__2_,
    P1_P1_INSTQUEUE_REG_12__1_, P1_P1_INSTQUEUE_REG_12__0_,
    P1_P1_INSTQUEUE_REG_11__7_, P1_P1_INSTQUEUE_REG_11__6_,
    P1_P1_INSTQUEUE_REG_11__5_, P1_P1_INSTQUEUE_REG_11__4_,
    P1_P1_INSTQUEUE_REG_11__3_, P1_P1_INSTQUEUE_REG_11__2_,
    P1_P1_INSTQUEUE_REG_11__1_, P1_P1_INSTQUEUE_REG_11__0_,
    P1_P1_INSTQUEUE_REG_10__7_, P1_P1_INSTQUEUE_REG_10__6_,
    P1_P1_INSTQUEUE_REG_10__5_, P1_P1_INSTQUEUE_REG_10__4_,
    P1_P1_INSTQUEUE_REG_10__3_, P1_P1_INSTQUEUE_REG_10__2_,
    P1_P1_INSTQUEUE_REG_10__1_, P1_P1_INSTQUEUE_REG_10__0_,
    P1_P1_INSTQUEUE_REG_9__7_, P1_P1_INSTQUEUE_REG_9__6_,
    P1_P1_INSTQUEUE_REG_9__5_, P1_P1_INSTQUEUE_REG_9__4_,
    P1_P1_INSTQUEUE_REG_9__3_, P1_P1_INSTQUEUE_REG_9__2_,
    P1_P1_INSTQUEUE_REG_9__1_, P1_P1_INSTQUEUE_REG_9__0_,
    P1_P1_INSTQUEUE_REG_8__7_, P1_P1_INSTQUEUE_REG_8__6_,
    P1_P1_INSTQUEUE_REG_8__5_, P1_P1_INSTQUEUE_REG_8__4_,
    P1_P1_INSTQUEUE_REG_8__3_, P1_P1_INSTQUEUE_REG_8__2_,
    P1_P1_INSTQUEUE_REG_8__1_, P1_P1_INSTQUEUE_REG_8__0_,
    P1_P1_INSTQUEUE_REG_7__7_, P1_P1_INSTQUEUE_REG_7__6_,
    P1_P1_INSTQUEUE_REG_7__5_, P1_P1_INSTQUEUE_REG_7__4_,
    P1_P1_INSTQUEUE_REG_7__3_, P1_P1_INSTQUEUE_REG_7__2_,
    P1_P1_INSTQUEUE_REG_7__1_, P1_P1_INSTQUEUE_REG_7__0_,
    P1_P1_INSTQUEUE_REG_6__7_, P1_P1_INSTQUEUE_REG_6__6_,
    P1_P1_INSTQUEUE_REG_6__5_, P1_P1_INSTQUEUE_REG_6__4_,
    P1_P1_INSTQUEUE_REG_6__3_, P1_P1_INSTQUEUE_REG_6__2_,
    P1_P1_INSTQUEUE_REG_6__1_, P1_P1_INSTQUEUE_REG_6__0_,
    P1_P1_INSTQUEUE_REG_5__7_, P1_P1_INSTQUEUE_REG_5__6_,
    P1_P1_INSTQUEUE_REG_5__5_, P1_P1_INSTQUEUE_REG_5__4_,
    P1_P1_INSTQUEUE_REG_5__3_, P1_P1_INSTQUEUE_REG_5__2_,
    P1_P1_INSTQUEUE_REG_5__1_, P1_P1_INSTQUEUE_REG_5__0_,
    P1_P1_INSTQUEUE_REG_4__7_, P1_P1_INSTQUEUE_REG_4__6_,
    P1_P1_INSTQUEUE_REG_4__5_, P1_P1_INSTQUEUE_REG_4__4_,
    P1_P1_INSTQUEUE_REG_4__3_, P1_P1_INSTQUEUE_REG_4__2_,
    P1_P1_INSTQUEUE_REG_4__1_, P1_P1_INSTQUEUE_REG_4__0_,
    P1_P1_INSTQUEUE_REG_3__7_, P1_P1_INSTQUEUE_REG_3__6_,
    P1_P1_INSTQUEUE_REG_3__5_, P1_P1_INSTQUEUE_REG_3__4_,
    P1_P1_INSTQUEUE_REG_3__3_, P1_P1_INSTQUEUE_REG_3__2_,
    P1_P1_INSTQUEUE_REG_3__1_, P1_P1_INSTQUEUE_REG_3__0_,
    P1_P1_INSTQUEUE_REG_2__7_, P1_P1_INSTQUEUE_REG_2__6_,
    P1_P1_INSTQUEUE_REG_2__5_, P1_P1_INSTQUEUE_REG_2__4_,
    P1_P1_INSTQUEUE_REG_2__3_, P1_P1_INSTQUEUE_REG_2__2_,
    P1_P1_INSTQUEUE_REG_2__1_, P1_P1_INSTQUEUE_REG_2__0_,
    P1_P1_INSTQUEUE_REG_1__7_, P1_P1_INSTQUEUE_REG_1__6_,
    P1_P1_INSTQUEUE_REG_1__5_, P1_P1_INSTQUEUE_REG_1__4_,
    P1_P1_INSTQUEUE_REG_1__3_, P1_P1_INSTQUEUE_REG_1__2_,
    P1_P1_INSTQUEUE_REG_1__1_, P1_P1_INSTQUEUE_REG_1__0_,
    P1_P1_INSTQUEUE_REG_0__7_, P1_P1_INSTQUEUE_REG_0__6_,
    P1_P1_INSTQUEUE_REG_0__5_, P1_P1_INSTQUEUE_REG_0__4_,
    P1_P1_INSTQUEUE_REG_0__3_, P1_P1_INSTQUEUE_REG_0__2_,
    P1_P1_INSTQUEUE_REG_0__1_, P1_P1_INSTQUEUE_REG_0__0_,
    P1_P1_INSTQUEUERD_ADDR_REG_4_, P1_P1_INSTQUEUERD_ADDR_REG_3_,
    P1_P1_INSTQUEUERD_ADDR_REG_2_, P1_P1_INSTQUEUERD_ADDR_REG_1_,
    P1_P1_INSTQUEUERD_ADDR_REG_0_, P1_P1_INSTQUEUEWR_ADDR_REG_4_,
    P1_P1_INSTQUEUEWR_ADDR_REG_3_, P1_P1_INSTQUEUEWR_ADDR_REG_2_,
    P1_P1_INSTQUEUEWR_ADDR_REG_1_, P1_P1_INSTQUEUEWR_ADDR_REG_0_,
    P1_P1_INSTADDRPOINTER_REG_0_, P1_P1_INSTADDRPOINTER_REG_1_,
    P1_P1_INSTADDRPOINTER_REG_2_, P1_P1_INSTADDRPOINTER_REG_3_,
    P1_P1_INSTADDRPOINTER_REG_4_, P1_P1_INSTADDRPOINTER_REG_5_,
    P1_P1_INSTADDRPOINTER_REG_6_, P1_P1_INSTADDRPOINTER_REG_7_,
    P1_P1_INSTADDRPOINTER_REG_8_, P1_P1_INSTADDRPOINTER_REG_9_,
    P1_P1_INSTADDRPOINTER_REG_10_, P1_P1_INSTADDRPOINTER_REG_11_,
    P1_P1_INSTADDRPOINTER_REG_12_, P1_P1_INSTADDRPOINTER_REG_13_,
    P1_P1_INSTADDRPOINTER_REG_14_, P1_P1_INSTADDRPOINTER_REG_15_,
    P1_P1_INSTADDRPOINTER_REG_16_, P1_P1_INSTADDRPOINTER_REG_17_,
    P1_P1_INSTADDRPOINTER_REG_18_, P1_P1_INSTADDRPOINTER_REG_19_,
    P1_P1_INSTADDRPOINTER_REG_20_, P1_P1_INSTADDRPOINTER_REG_21_,
    P1_P1_INSTADDRPOINTER_REG_22_, P1_P1_INSTADDRPOINTER_REG_23_,
    P1_P1_INSTADDRPOINTER_REG_24_, P1_P1_INSTADDRPOINTER_REG_25_,
    P1_P1_INSTADDRPOINTER_REG_26_, P1_P1_INSTADDRPOINTER_REG_27_,
    P1_P1_INSTADDRPOINTER_REG_28_, P1_P1_INSTADDRPOINTER_REG_29_,
    P1_P1_INSTADDRPOINTER_REG_30_, P1_P1_INSTADDRPOINTER_REG_31_,
    P1_P1_PHYADDRPOINTER_REG_0_, P1_P1_PHYADDRPOINTER_REG_1_,
    P1_P1_PHYADDRPOINTER_REG_2_, P1_P1_PHYADDRPOINTER_REG_3_,
    P1_P1_PHYADDRPOINTER_REG_4_, P1_P1_PHYADDRPOINTER_REG_5_,
    P1_P1_PHYADDRPOINTER_REG_6_, P1_P1_PHYADDRPOINTER_REG_7_,
    P1_P1_PHYADDRPOINTER_REG_8_, P1_P1_PHYADDRPOINTER_REG_9_,
    P1_P1_PHYADDRPOINTER_REG_10_, P1_P1_PHYADDRPOINTER_REG_11_,
    P1_P1_PHYADDRPOINTER_REG_12_, P1_P1_PHYADDRPOINTER_REG_13_,
    P1_P1_PHYADDRPOINTER_REG_14_, P1_P1_PHYADDRPOINTER_REG_15_,
    P1_P1_PHYADDRPOINTER_REG_16_, P1_P1_PHYADDRPOINTER_REG_17_,
    P1_P1_PHYADDRPOINTER_REG_18_, P1_P1_PHYADDRPOINTER_REG_19_,
    P1_P1_PHYADDRPOINTER_REG_20_, P1_P1_PHYADDRPOINTER_REG_21_,
    P1_P1_PHYADDRPOINTER_REG_22_, P1_P1_PHYADDRPOINTER_REG_23_,
    P1_P1_PHYADDRPOINTER_REG_24_, P1_P1_PHYADDRPOINTER_REG_25_,
    P1_P1_PHYADDRPOINTER_REG_26_, P1_P1_PHYADDRPOINTER_REG_27_,
    P1_P1_PHYADDRPOINTER_REG_28_, P1_P1_PHYADDRPOINTER_REG_29_,
    P1_P1_PHYADDRPOINTER_REG_30_, P1_P1_PHYADDRPOINTER_REG_31_,
    P1_P1_LWORD_REG_15_, P1_P1_LWORD_REG_14_, P1_P1_LWORD_REG_13_,
    P1_P1_LWORD_REG_12_, P1_P1_LWORD_REG_11_, P1_P1_LWORD_REG_10_,
    P1_P1_LWORD_REG_9_, P1_P1_LWORD_REG_8_, P1_P1_LWORD_REG_7_,
    P1_P1_LWORD_REG_6_, P1_P1_LWORD_REG_5_, P1_P1_LWORD_REG_4_,
    P1_P1_LWORD_REG_3_, P1_P1_LWORD_REG_2_, P1_P1_LWORD_REG_1_,
    P1_P1_LWORD_REG_0_, P1_P1_UWORD_REG_14_, P1_P1_UWORD_REG_13_,
    P1_P1_UWORD_REG_12_, P1_P1_UWORD_REG_11_, P1_P1_UWORD_REG_10_,
    P1_P1_UWORD_REG_9_, P1_P1_UWORD_REG_8_, P1_P1_UWORD_REG_7_,
    P1_P1_UWORD_REG_6_, P1_P1_UWORD_REG_5_, P1_P1_UWORD_REG_4_,
    P1_P1_UWORD_REG_3_, P1_P1_UWORD_REG_2_, P1_P1_UWORD_REG_1_,
    P1_P1_UWORD_REG_0_, P1_P1_DATAO_REG_0_, P1_P1_DATAO_REG_1_,
    P1_P1_DATAO_REG_2_, P1_P1_DATAO_REG_3_, P1_P1_DATAO_REG_4_,
    P1_P1_DATAO_REG_5_, P1_P1_DATAO_REG_6_, P1_P1_DATAO_REG_7_,
    P1_P1_DATAO_REG_8_, P1_P1_DATAO_REG_9_, P1_P1_DATAO_REG_10_,
    P1_P1_DATAO_REG_11_, P1_P1_DATAO_REG_12_, P1_P1_DATAO_REG_13_,
    P1_P1_DATAO_REG_14_, P1_P1_DATAO_REG_15_, P1_P1_DATAO_REG_16_,
    P1_P1_DATAO_REG_17_, P1_P1_DATAO_REG_18_, P1_P1_DATAO_REG_19_,
    P1_P1_DATAO_REG_20_, P1_P1_DATAO_REG_21_, P1_P1_DATAO_REG_22_,
    P1_P1_DATAO_REG_23_, P1_P1_DATAO_REG_24_, P1_P1_DATAO_REG_25_,
    P1_P1_DATAO_REG_26_, P1_P1_DATAO_REG_27_, P1_P1_DATAO_REG_28_,
    P1_P1_DATAO_REG_29_, P1_P1_DATAO_REG_30_, P1_P1_DATAO_REG_31_,
    P1_P1_EAX_REG_0_, P1_P1_EAX_REG_1_, P1_P1_EAX_REG_2_, P1_P1_EAX_REG_3_,
    P1_P1_EAX_REG_4_, P1_P1_EAX_REG_5_, P1_P1_EAX_REG_6_, P1_P1_EAX_REG_7_,
    P1_P1_EAX_REG_8_, P1_P1_EAX_REG_9_, P1_P1_EAX_REG_10_,
    P1_P1_EAX_REG_11_, P1_P1_EAX_REG_12_, P1_P1_EAX_REG_13_,
    P1_P1_EAX_REG_14_, P1_P1_EAX_REG_15_, P1_P1_EAX_REG_16_,
    P1_P1_EAX_REG_17_, P1_P1_EAX_REG_18_, P1_P1_EAX_REG_19_,
    P1_P1_EAX_REG_20_, P1_P1_EAX_REG_21_, P1_P1_EAX_REG_22_,
    P1_P1_EAX_REG_23_, P1_P1_EAX_REG_24_, P1_P1_EAX_REG_25_,
    P1_P1_EAX_REG_26_, P1_P1_EAX_REG_27_, P1_P1_EAX_REG_28_,
    P1_P1_EAX_REG_29_, P1_P1_EAX_REG_30_, P1_P1_EAX_REG_31_,
    P1_P1_EBX_REG_0_, P1_P1_EBX_REG_1_, P1_P1_EBX_REG_2_, P1_P1_EBX_REG_3_,
    P1_P1_EBX_REG_4_, P1_P1_EBX_REG_5_, P1_P1_EBX_REG_6_, P1_P1_EBX_REG_7_,
    P1_P1_EBX_REG_8_, P1_P1_EBX_REG_9_, P1_P1_EBX_REG_10_,
    P1_P1_EBX_REG_11_, P1_P1_EBX_REG_12_, P1_P1_EBX_REG_13_,
    P1_P1_EBX_REG_14_, P1_P1_EBX_REG_15_, P1_P1_EBX_REG_16_,
    P1_P1_EBX_REG_17_, P1_P1_EBX_REG_18_, P1_P1_EBX_REG_19_,
    P1_P1_EBX_REG_20_, P1_P1_EBX_REG_21_, P1_P1_EBX_REG_22_,
    P1_P1_EBX_REG_23_, P1_P1_EBX_REG_24_, P1_P1_EBX_REG_25_,
    P1_P1_EBX_REG_26_, P1_P1_EBX_REG_27_, P1_P1_EBX_REG_28_,
    P1_P1_EBX_REG_29_, P1_P1_EBX_REG_30_, P1_P1_EBX_REG_31_,
    P1_P1_REIP_REG_0_, P1_P1_REIP_REG_1_, P1_P1_REIP_REG_2_,
    P1_P1_REIP_REG_3_, P1_P1_REIP_REG_4_, P1_P1_REIP_REG_5_,
    P1_P1_REIP_REG_6_, P1_P1_REIP_REG_7_, P1_P1_REIP_REG_8_,
    P1_P1_REIP_REG_9_, P1_P1_REIP_REG_10_, P1_P1_REIP_REG_11_,
    P1_P1_REIP_REG_12_, P1_P1_REIP_REG_13_, P1_P1_REIP_REG_14_,
    P1_P1_REIP_REG_15_, P1_P1_REIP_REG_16_, P1_P1_REIP_REG_17_,
    P1_P1_REIP_REG_18_, P1_P1_REIP_REG_19_, P1_P1_REIP_REG_20_,
    P1_P1_REIP_REG_21_, P1_P1_REIP_REG_22_, P1_P1_REIP_REG_23_,
    P1_P1_REIP_REG_24_, P1_P1_REIP_REG_25_, P1_P1_REIP_REG_26_,
    P1_P1_REIP_REG_27_, P1_P1_REIP_REG_28_, P1_P1_REIP_REG_29_,
    P1_P1_REIP_REG_30_, P1_P1_REIP_REG_31_, P1_P1_BYTEENABLE_REG_3_,
    P1_P1_BYTEENABLE_REG_2_, P1_P1_BYTEENABLE_REG_1_,
    P1_P1_BYTEENABLE_REG_0_, P1_P1_W_R_N_REG, P1_P1_FLUSH_REG,
    P1_P1_MORE_REG, P1_P1_STATEBS16_REG, P1_P1_REQUESTPENDING_REG,
    P1_P1_D_C_N_REG, P1_P1_M_IO_N_REG, P1_P1_CODEFETCH_REG,
    P1_P1_ADS_N_REG, P1_P1_READREQUEST_REG, P1_P1_MEMORYFETCH_REG,
    P2_P3_BE_N_REG_3_, P2_P3_BE_N_REG_2_, P2_P3_BE_N_REG_1_,
    P2_P3_BE_N_REG_0_, P2_P3_ADDRESS_REG_29_, P2_P3_ADDRESS_REG_28_,
    P2_P3_ADDRESS_REG_27_, P2_P3_ADDRESS_REG_26_, P2_P3_ADDRESS_REG_25_,
    P2_P3_ADDRESS_REG_24_, P2_P3_ADDRESS_REG_23_, P2_P3_ADDRESS_REG_22_,
    P2_P3_ADDRESS_REG_21_, P2_P3_ADDRESS_REG_20_, P2_P3_ADDRESS_REG_19_,
    P2_P3_ADDRESS_REG_18_, P2_P3_ADDRESS_REG_17_, P2_P3_ADDRESS_REG_16_,
    P2_P3_ADDRESS_REG_15_, P2_P3_ADDRESS_REG_14_, P2_P3_ADDRESS_REG_13_,
    P2_P3_ADDRESS_REG_12_, P2_P3_ADDRESS_REG_11_, P2_P3_ADDRESS_REG_10_,
    P2_P3_ADDRESS_REG_9_, P2_P3_ADDRESS_REG_8_, P2_P3_ADDRESS_REG_7_,
    P2_P3_ADDRESS_REG_6_, P2_P3_ADDRESS_REG_5_, P2_P3_ADDRESS_REG_4_,
    P2_P3_ADDRESS_REG_3_, P2_P3_ADDRESS_REG_2_, P2_P3_ADDRESS_REG_1_,
    P2_P3_ADDRESS_REG_0_, P2_P3_STATE_REG_2_, P2_P3_STATE_REG_1_,
    P2_P3_STATE_REG_0_, P2_P3_DATAWIDTH_REG_0_, P2_P3_DATAWIDTH_REG_1_,
    P2_P3_DATAWIDTH_REG_2_, P2_P3_DATAWIDTH_REG_3_, P2_P3_DATAWIDTH_REG_4_,
    P2_P3_DATAWIDTH_REG_5_, P2_P3_DATAWIDTH_REG_6_, P2_P3_DATAWIDTH_REG_7_,
    P2_P3_DATAWIDTH_REG_8_, P2_P3_DATAWIDTH_REG_9_,
    P2_P3_DATAWIDTH_REG_10_, P2_P3_DATAWIDTH_REG_11_,
    P2_P3_DATAWIDTH_REG_12_, P2_P3_DATAWIDTH_REG_13_,
    P2_P3_DATAWIDTH_REG_14_, P2_P3_DATAWIDTH_REG_15_,
    P2_P3_DATAWIDTH_REG_16_, P2_P3_DATAWIDTH_REG_17_,
    P2_P3_DATAWIDTH_REG_18_, P2_P3_DATAWIDTH_REG_19_,
    P2_P3_DATAWIDTH_REG_20_, P2_P3_DATAWIDTH_REG_21_,
    P2_P3_DATAWIDTH_REG_22_, P2_P3_DATAWIDTH_REG_23_,
    P2_P3_DATAWIDTH_REG_24_, P2_P3_DATAWIDTH_REG_25_,
    P2_P3_DATAWIDTH_REG_26_, P2_P3_DATAWIDTH_REG_27_,
    P2_P3_DATAWIDTH_REG_28_, P2_P3_DATAWIDTH_REG_29_,
    P2_P3_DATAWIDTH_REG_30_, P2_P3_DATAWIDTH_REG_31_, P2_P3_STATE2_REG_3_,
    P2_P3_STATE2_REG_2_, P2_P3_STATE2_REG_1_, P2_P3_STATE2_REG_0_,
    P2_P3_INSTQUEUE_REG_15__7_, P2_P3_INSTQUEUE_REG_15__6_,
    P2_P3_INSTQUEUE_REG_15__5_, P2_P3_INSTQUEUE_REG_15__4_,
    P2_P3_INSTQUEUE_REG_15__3_, P2_P3_INSTQUEUE_REG_15__2_,
    P2_P3_INSTQUEUE_REG_15__1_, P2_P3_INSTQUEUE_REG_15__0_,
    P2_P3_INSTQUEUE_REG_14__7_, P2_P3_INSTQUEUE_REG_14__6_,
    P2_P3_INSTQUEUE_REG_14__5_, P2_P3_INSTQUEUE_REG_14__4_,
    P2_P3_INSTQUEUE_REG_14__3_, P2_P3_INSTQUEUE_REG_14__2_,
    P2_P3_INSTQUEUE_REG_14__1_, P2_P3_INSTQUEUE_REG_14__0_,
    P2_P3_INSTQUEUE_REG_13__7_, P2_P3_INSTQUEUE_REG_13__6_,
    P2_P3_INSTQUEUE_REG_13__5_, P2_P3_INSTQUEUE_REG_13__4_,
    P2_P3_INSTQUEUE_REG_13__3_, P2_P3_INSTQUEUE_REG_13__2_,
    P2_P3_INSTQUEUE_REG_13__1_, P2_P3_INSTQUEUE_REG_13__0_,
    P2_P3_INSTQUEUE_REG_12__7_, P2_P3_INSTQUEUE_REG_12__6_,
    P2_P3_INSTQUEUE_REG_12__5_, P2_P3_INSTQUEUE_REG_12__4_,
    P2_P3_INSTQUEUE_REG_12__3_, P2_P3_INSTQUEUE_REG_12__2_,
    P2_P3_INSTQUEUE_REG_12__1_, P2_P3_INSTQUEUE_REG_12__0_,
    P2_P3_INSTQUEUE_REG_11__7_, P2_P3_INSTQUEUE_REG_11__6_,
    P2_P3_INSTQUEUE_REG_11__5_, P2_P3_INSTQUEUE_REG_11__4_,
    P2_P3_INSTQUEUE_REG_11__3_, P2_P3_INSTQUEUE_REG_11__2_,
    P2_P3_INSTQUEUE_REG_11__1_, P2_P3_INSTQUEUE_REG_11__0_,
    P2_P3_INSTQUEUE_REG_10__7_, P2_P3_INSTQUEUE_REG_10__6_,
    P2_P3_INSTQUEUE_REG_10__5_, P2_P3_INSTQUEUE_REG_10__4_,
    P2_P3_INSTQUEUE_REG_10__3_, P2_P3_INSTQUEUE_REG_10__2_,
    P2_P3_INSTQUEUE_REG_10__1_, P2_P3_INSTQUEUE_REG_10__0_,
    P2_P3_INSTQUEUE_REG_9__7_, P2_P3_INSTQUEUE_REG_9__6_,
    P2_P3_INSTQUEUE_REG_9__5_, P2_P3_INSTQUEUE_REG_9__4_,
    P2_P3_INSTQUEUE_REG_9__3_, P2_P3_INSTQUEUE_REG_9__2_,
    P2_P3_INSTQUEUE_REG_9__1_, P2_P3_INSTQUEUE_REG_9__0_,
    P2_P3_INSTQUEUE_REG_8__7_, P2_P3_INSTQUEUE_REG_8__6_,
    P2_P3_INSTQUEUE_REG_8__5_, P2_P3_INSTQUEUE_REG_8__4_,
    P2_P3_INSTQUEUE_REG_8__3_, P2_P3_INSTQUEUE_REG_8__2_,
    P2_P3_INSTQUEUE_REG_8__1_, P2_P3_INSTQUEUE_REG_8__0_,
    P2_P3_INSTQUEUE_REG_7__7_, P2_P3_INSTQUEUE_REG_7__6_,
    P2_P3_INSTQUEUE_REG_7__5_, P2_P3_INSTQUEUE_REG_7__4_,
    P2_P3_INSTQUEUE_REG_7__3_, P2_P3_INSTQUEUE_REG_7__2_,
    P2_P3_INSTQUEUE_REG_7__1_, P2_P3_INSTQUEUE_REG_7__0_,
    P2_P3_INSTQUEUE_REG_6__7_, P2_P3_INSTQUEUE_REG_6__6_,
    P2_P3_INSTQUEUE_REG_6__5_, P2_P3_INSTQUEUE_REG_6__4_,
    P2_P3_INSTQUEUE_REG_6__3_, P2_P3_INSTQUEUE_REG_6__2_,
    P2_P3_INSTQUEUE_REG_6__1_, P2_P3_INSTQUEUE_REG_6__0_,
    P2_P3_INSTQUEUE_REG_5__7_, P2_P3_INSTQUEUE_REG_5__6_,
    P2_P3_INSTQUEUE_REG_5__5_, P2_P3_INSTQUEUE_REG_5__4_,
    P2_P3_INSTQUEUE_REG_5__3_, P2_P3_INSTQUEUE_REG_5__2_,
    P2_P3_INSTQUEUE_REG_5__1_, P2_P3_INSTQUEUE_REG_5__0_,
    P2_P3_INSTQUEUE_REG_4__7_, P2_P3_INSTQUEUE_REG_4__6_,
    P2_P3_INSTQUEUE_REG_4__5_, P2_P3_INSTQUEUE_REG_4__4_,
    P2_P3_INSTQUEUE_REG_4__3_, P2_P3_INSTQUEUE_REG_4__2_,
    P2_P3_INSTQUEUE_REG_4__1_, P2_P3_INSTQUEUE_REG_4__0_,
    P2_P3_INSTQUEUE_REG_3__7_, P2_P3_INSTQUEUE_REG_3__6_,
    P2_P3_INSTQUEUE_REG_3__5_, P2_P3_INSTQUEUE_REG_3__4_,
    P2_P3_INSTQUEUE_REG_3__3_, P2_P3_INSTQUEUE_REG_3__2_,
    P2_P3_INSTQUEUE_REG_3__1_, P2_P3_INSTQUEUE_REG_3__0_,
    P2_P3_INSTQUEUE_REG_2__7_, P2_P3_INSTQUEUE_REG_2__6_,
    P2_P3_INSTQUEUE_REG_2__5_, P2_P3_INSTQUEUE_REG_2__4_,
    P2_P3_INSTQUEUE_REG_2__3_, P2_P3_INSTQUEUE_REG_2__2_,
    P2_P3_INSTQUEUE_REG_2__1_, P2_P3_INSTQUEUE_REG_2__0_,
    P2_P3_INSTQUEUE_REG_1__7_, P2_P3_INSTQUEUE_REG_1__6_,
    P2_P3_INSTQUEUE_REG_1__5_, P2_P3_INSTQUEUE_REG_1__4_,
    P2_P3_INSTQUEUE_REG_1__3_, P2_P3_INSTQUEUE_REG_1__2_,
    P2_P3_INSTQUEUE_REG_1__1_, P2_P3_INSTQUEUE_REG_1__0_,
    P2_P3_INSTQUEUE_REG_0__7_, P2_P3_INSTQUEUE_REG_0__6_,
    P2_P3_INSTQUEUE_REG_0__5_, P2_P3_INSTQUEUE_REG_0__4_,
    P2_P3_INSTQUEUE_REG_0__3_, P2_P3_INSTQUEUE_REG_0__2_,
    P2_P3_INSTQUEUE_REG_0__1_, P2_P3_INSTQUEUE_REG_0__0_,
    P2_P3_INSTQUEUERD_ADDR_REG_4_, P2_P3_INSTQUEUERD_ADDR_REG_3_,
    P2_P3_INSTQUEUERD_ADDR_REG_2_, P2_P3_INSTQUEUERD_ADDR_REG_1_,
    P2_P3_INSTQUEUERD_ADDR_REG_0_, P2_P3_INSTQUEUEWR_ADDR_REG_4_,
    P2_P3_INSTQUEUEWR_ADDR_REG_3_, P2_P3_INSTQUEUEWR_ADDR_REG_2_,
    P2_P3_INSTQUEUEWR_ADDR_REG_1_, P2_P3_INSTQUEUEWR_ADDR_REG_0_,
    P2_P3_INSTADDRPOINTER_REG_0_, P2_P3_INSTADDRPOINTER_REG_1_,
    P2_P3_INSTADDRPOINTER_REG_2_, P2_P3_INSTADDRPOINTER_REG_3_,
    P2_P3_INSTADDRPOINTER_REG_4_, P2_P3_INSTADDRPOINTER_REG_5_,
    P2_P3_INSTADDRPOINTER_REG_6_, P2_P3_INSTADDRPOINTER_REG_7_,
    P2_P3_INSTADDRPOINTER_REG_8_, P2_P3_INSTADDRPOINTER_REG_9_,
    P2_P3_INSTADDRPOINTER_REG_10_, P2_P3_INSTADDRPOINTER_REG_11_,
    P2_P3_INSTADDRPOINTER_REG_12_, P2_P3_INSTADDRPOINTER_REG_13_,
    P2_P3_INSTADDRPOINTER_REG_14_, P2_P3_INSTADDRPOINTER_REG_15_,
    P2_P3_INSTADDRPOINTER_REG_16_, P2_P3_INSTADDRPOINTER_REG_17_,
    P2_P3_INSTADDRPOINTER_REG_18_, P2_P3_INSTADDRPOINTER_REG_19_,
    P2_P3_INSTADDRPOINTER_REG_20_, P2_P3_INSTADDRPOINTER_REG_21_,
    P2_P3_INSTADDRPOINTER_REG_22_, P2_P3_INSTADDRPOINTER_REG_23_,
    P2_P3_INSTADDRPOINTER_REG_24_, P2_P3_INSTADDRPOINTER_REG_25_,
    P2_P3_INSTADDRPOINTER_REG_26_, P2_P3_INSTADDRPOINTER_REG_27_,
    P2_P3_INSTADDRPOINTER_REG_28_, P2_P3_INSTADDRPOINTER_REG_29_,
    P2_P3_INSTADDRPOINTER_REG_30_, P2_P3_INSTADDRPOINTER_REG_31_,
    P2_P3_PHYADDRPOINTER_REG_0_, P2_P3_PHYADDRPOINTER_REG_1_,
    P2_P3_PHYADDRPOINTER_REG_2_, P2_P3_PHYADDRPOINTER_REG_3_,
    P2_P3_PHYADDRPOINTER_REG_4_, P2_P3_PHYADDRPOINTER_REG_5_,
    P2_P3_PHYADDRPOINTER_REG_6_, P2_P3_PHYADDRPOINTER_REG_7_,
    P2_P3_PHYADDRPOINTER_REG_8_, P2_P3_PHYADDRPOINTER_REG_9_,
    P2_P3_PHYADDRPOINTER_REG_10_, P2_P3_PHYADDRPOINTER_REG_11_,
    P2_P3_PHYADDRPOINTER_REG_12_, P2_P3_PHYADDRPOINTER_REG_13_,
    P2_P3_PHYADDRPOINTER_REG_14_, P2_P3_PHYADDRPOINTER_REG_15_,
    P2_P3_PHYADDRPOINTER_REG_16_, P2_P3_PHYADDRPOINTER_REG_17_,
    P2_P3_PHYADDRPOINTER_REG_18_, P2_P3_PHYADDRPOINTER_REG_19_,
    P2_P3_PHYADDRPOINTER_REG_20_, P2_P3_PHYADDRPOINTER_REG_21_,
    P2_P3_PHYADDRPOINTER_REG_22_, P2_P3_PHYADDRPOINTER_REG_23_,
    P2_P3_PHYADDRPOINTER_REG_24_, P2_P3_PHYADDRPOINTER_REG_25_,
    P2_P3_PHYADDRPOINTER_REG_26_, P2_P3_PHYADDRPOINTER_REG_27_,
    P2_P3_PHYADDRPOINTER_REG_28_, P2_P3_PHYADDRPOINTER_REG_29_,
    P2_P3_PHYADDRPOINTER_REG_30_, P2_P3_PHYADDRPOINTER_REG_31_,
    P2_P3_LWORD_REG_15_, P2_P3_LWORD_REG_14_, P2_P3_LWORD_REG_13_,
    P2_P3_LWORD_REG_12_, P2_P3_LWORD_REG_11_, P2_P3_LWORD_REG_10_,
    P2_P3_LWORD_REG_9_, P2_P3_LWORD_REG_8_, P2_P3_LWORD_REG_7_,
    P2_P3_LWORD_REG_6_, P2_P3_LWORD_REG_5_, P2_P3_LWORD_REG_4_,
    P2_P3_LWORD_REG_3_, P2_P3_LWORD_REG_2_, P2_P3_LWORD_REG_1_,
    P2_P3_LWORD_REG_0_, P2_P3_UWORD_REG_14_, P2_P3_UWORD_REG_13_,
    P2_P3_UWORD_REG_12_, P2_P3_UWORD_REG_11_, P2_P3_UWORD_REG_10_,
    P2_P3_UWORD_REG_9_, P2_P3_UWORD_REG_8_, P2_P3_UWORD_REG_7_,
    P2_P3_UWORD_REG_6_, P2_P3_UWORD_REG_5_, P2_P3_UWORD_REG_4_,
    P2_P3_UWORD_REG_3_, P2_P3_UWORD_REG_2_, P2_P3_UWORD_REG_1_,
    P2_P3_UWORD_REG_0_, P2_P3_DATAO_REG_0_, P2_P3_DATAO_REG_1_,
    P2_P3_DATAO_REG_2_, P2_P3_DATAO_REG_3_, P2_P3_DATAO_REG_4_,
    P2_P3_DATAO_REG_5_, P2_P3_DATAO_REG_6_, P2_P3_DATAO_REG_7_,
    P2_P3_DATAO_REG_8_, P2_P3_DATAO_REG_9_, P2_P3_DATAO_REG_10_,
    P2_P3_DATAO_REG_11_, P2_P3_DATAO_REG_12_, P2_P3_DATAO_REG_13_,
    P2_P3_DATAO_REG_14_, P2_P3_DATAO_REG_15_, P2_P3_DATAO_REG_16_,
    P2_P3_DATAO_REG_17_, P2_P3_DATAO_REG_18_, P2_P3_DATAO_REG_19_,
    P2_P3_DATAO_REG_20_, P2_P3_DATAO_REG_21_, P2_P3_DATAO_REG_22_,
    P2_P3_DATAO_REG_23_, P2_P3_DATAO_REG_24_, P2_P3_DATAO_REG_25_,
    P2_P3_DATAO_REG_26_, P2_P3_DATAO_REG_27_, P2_P3_DATAO_REG_28_,
    P2_P3_DATAO_REG_29_, P2_P3_DATAO_REG_30_, P2_P3_DATAO_REG_31_,
    P2_P3_EAX_REG_0_, P2_P3_EAX_REG_1_, P2_P3_EAX_REG_2_, P2_P3_EAX_REG_3_,
    P2_P3_EAX_REG_4_, P2_P3_EAX_REG_5_, P2_P3_EAX_REG_6_, P2_P3_EAX_REG_7_,
    P2_P3_EAX_REG_8_, P2_P3_EAX_REG_9_, P2_P3_EAX_REG_10_,
    P2_P3_EAX_REG_11_, P2_P3_EAX_REG_12_, P2_P3_EAX_REG_13_,
    P2_P3_EAX_REG_14_, P2_P3_EAX_REG_15_, P2_P3_EAX_REG_16_,
    P2_P3_EAX_REG_17_, P2_P3_EAX_REG_18_, P2_P3_EAX_REG_19_,
    P2_P3_EAX_REG_20_, P2_P3_EAX_REG_21_, P2_P3_EAX_REG_22_,
    P2_P3_EAX_REG_23_, P2_P3_EAX_REG_24_, P2_P3_EAX_REG_25_,
    P2_P3_EAX_REG_26_, P2_P3_EAX_REG_27_, P2_P3_EAX_REG_28_,
    P2_P3_EAX_REG_29_, P2_P3_EAX_REG_30_, P2_P3_EAX_REG_31_,
    P2_P3_EBX_REG_0_, P2_P3_EBX_REG_1_, P2_P3_EBX_REG_2_, P2_P3_EBX_REG_3_,
    P2_P3_EBX_REG_4_, P2_P3_EBX_REG_5_, P2_P3_EBX_REG_6_, P2_P3_EBX_REG_7_,
    P2_P3_EBX_REG_8_, P2_P3_EBX_REG_9_, P2_P3_EBX_REG_10_,
    P2_P3_EBX_REG_11_, P2_P3_EBX_REG_12_, P2_P3_EBX_REG_13_,
    P2_P3_EBX_REG_14_, P2_P3_EBX_REG_15_, P2_P3_EBX_REG_16_,
    P2_P3_EBX_REG_17_, P2_P3_EBX_REG_18_, P2_P3_EBX_REG_19_,
    P2_P3_EBX_REG_20_, P2_P3_EBX_REG_21_, P2_P3_EBX_REG_22_,
    P2_P3_EBX_REG_23_, P2_P3_EBX_REG_24_, P2_P3_EBX_REG_25_,
    P2_P3_EBX_REG_26_, P2_P3_EBX_REG_27_, P2_P3_EBX_REG_28_,
    P2_P3_EBX_REG_29_, P2_P3_EBX_REG_30_, P2_P3_EBX_REG_31_,
    P2_P3_REIP_REG_0_, P2_P3_REIP_REG_1_, P2_P3_REIP_REG_2_,
    P2_P3_REIP_REG_3_, P2_P3_REIP_REG_4_, P2_P3_REIP_REG_5_,
    P2_P3_REIP_REG_6_, P2_P3_REIP_REG_7_, P2_P3_REIP_REG_8_,
    P2_P3_REIP_REG_9_, P2_P3_REIP_REG_10_, P2_P3_REIP_REG_11_,
    P2_P3_REIP_REG_12_, P2_P3_REIP_REG_13_, P2_P3_REIP_REG_14_,
    P2_P3_REIP_REG_15_, P2_P3_REIP_REG_16_, P2_P3_REIP_REG_17_,
    P2_P3_REIP_REG_18_, P2_P3_REIP_REG_19_, P2_P3_REIP_REG_20_,
    P2_P3_REIP_REG_21_, P2_P3_REIP_REG_22_, P2_P3_REIP_REG_23_,
    P2_P3_REIP_REG_24_, P2_P3_REIP_REG_25_, P2_P3_REIP_REG_26_,
    P2_P3_REIP_REG_27_, P2_P3_REIP_REG_28_, P2_P3_REIP_REG_29_,
    P2_P3_REIP_REG_30_, P2_P3_REIP_REG_31_, P2_P3_BYTEENABLE_REG_3_,
    P2_P3_BYTEENABLE_REG_2_, P2_P3_BYTEENABLE_REG_1_,
    P2_P3_BYTEENABLE_REG_0_, P2_P3_W_R_N_REG, P2_P3_FLUSH_REG,
    P2_P3_MORE_REG, P2_P3_STATEBS16_REG, P2_P3_REQUESTPENDING_REG,
    P2_P3_D_C_N_REG, P2_P3_M_IO_N_REG, P2_P3_CODEFETCH_REG,
    P2_P3_ADS_N_REG, P2_P3_READREQUEST_REG, P2_P3_MEMORYFETCH_REG,
    P2_P2_BE_N_REG_3_, P2_P2_BE_N_REG_2_, P2_P2_BE_N_REG_1_,
    P2_P2_BE_N_REG_0_, P2_P2_ADDRESS_REG_29_, P2_P2_ADDRESS_REG_28_,
    P2_P2_ADDRESS_REG_27_, P2_P2_ADDRESS_REG_26_, P2_P2_ADDRESS_REG_25_,
    P2_P2_ADDRESS_REG_24_, P2_P2_ADDRESS_REG_23_, P2_P2_ADDRESS_REG_22_,
    P2_P2_ADDRESS_REG_21_, P2_P2_ADDRESS_REG_20_, P2_P2_ADDRESS_REG_19_,
    P2_P2_ADDRESS_REG_18_, P2_P2_ADDRESS_REG_17_, P2_P2_ADDRESS_REG_16_,
    P2_P2_ADDRESS_REG_15_, P2_P2_ADDRESS_REG_14_, P2_P2_ADDRESS_REG_13_,
    P2_P2_ADDRESS_REG_12_, P2_P2_ADDRESS_REG_11_, P2_P2_ADDRESS_REG_10_,
    P2_P2_ADDRESS_REG_9_, P2_P2_ADDRESS_REG_8_, P2_P2_ADDRESS_REG_7_,
    P2_P2_ADDRESS_REG_6_, P2_P2_ADDRESS_REG_5_, P2_P2_ADDRESS_REG_4_,
    P2_P2_ADDRESS_REG_3_, P2_P2_ADDRESS_REG_2_, P2_P2_ADDRESS_REG_1_,
    P2_P2_ADDRESS_REG_0_, P2_P2_STATE_REG_2_, P2_P2_STATE_REG_1_,
    P2_P2_STATE_REG_0_, P2_P2_DATAWIDTH_REG_0_, P2_P2_DATAWIDTH_REG_1_,
    P2_P2_DATAWIDTH_REG_2_, P2_P2_DATAWIDTH_REG_3_, P2_P2_DATAWIDTH_REG_4_,
    P2_P2_DATAWIDTH_REG_5_, P2_P2_DATAWIDTH_REG_6_, P2_P2_DATAWIDTH_REG_7_,
    P2_P2_DATAWIDTH_REG_8_, P2_P2_DATAWIDTH_REG_9_,
    P2_P2_DATAWIDTH_REG_10_, P2_P2_DATAWIDTH_REG_11_,
    P2_P2_DATAWIDTH_REG_12_, P2_P2_DATAWIDTH_REG_13_,
    P2_P2_DATAWIDTH_REG_14_, P2_P2_DATAWIDTH_REG_15_,
    P2_P2_DATAWIDTH_REG_16_, P2_P2_DATAWIDTH_REG_17_,
    P2_P2_DATAWIDTH_REG_18_, P2_P2_DATAWIDTH_REG_19_,
    P2_P2_DATAWIDTH_REG_20_, P2_P2_DATAWIDTH_REG_21_,
    P2_P2_DATAWIDTH_REG_22_, P2_P2_DATAWIDTH_REG_23_,
    P2_P2_DATAWIDTH_REG_24_, P2_P2_DATAWIDTH_REG_25_,
    P2_P2_DATAWIDTH_REG_26_, P2_P2_DATAWIDTH_REG_27_,
    P2_P2_DATAWIDTH_REG_28_, P2_P2_DATAWIDTH_REG_29_,
    P2_P2_DATAWIDTH_REG_30_, P2_P2_DATAWIDTH_REG_31_, P2_P2_STATE2_REG_3_,
    P2_P2_STATE2_REG_2_, P2_P2_STATE2_REG_1_, P2_P2_STATE2_REG_0_,
    P2_P2_INSTQUEUE_REG_15__7_, P2_P2_INSTQUEUE_REG_15__6_,
    P2_P2_INSTQUEUE_REG_15__5_, P2_P2_INSTQUEUE_REG_15__4_,
    P2_P2_INSTQUEUE_REG_15__3_, P2_P2_INSTQUEUE_REG_15__2_,
    P2_P2_INSTQUEUE_REG_15__1_, P2_P2_INSTQUEUE_REG_15__0_,
    P2_P2_INSTQUEUE_REG_14__7_, P2_P2_INSTQUEUE_REG_14__6_,
    P2_P2_INSTQUEUE_REG_14__5_, P2_P2_INSTQUEUE_REG_14__4_,
    P2_P2_INSTQUEUE_REG_14__3_, P2_P2_INSTQUEUE_REG_14__2_,
    P2_P2_INSTQUEUE_REG_14__1_, P2_P2_INSTQUEUE_REG_14__0_,
    P2_P2_INSTQUEUE_REG_13__7_, P2_P2_INSTQUEUE_REG_13__6_,
    P2_P2_INSTQUEUE_REG_13__5_, P2_P2_INSTQUEUE_REG_13__4_,
    P2_P2_INSTQUEUE_REG_13__3_, P2_P2_INSTQUEUE_REG_13__2_,
    P2_P2_INSTQUEUE_REG_13__1_, P2_P2_INSTQUEUE_REG_13__0_,
    P2_P2_INSTQUEUE_REG_12__7_, P2_P2_INSTQUEUE_REG_12__6_,
    P2_P2_INSTQUEUE_REG_12__5_, P2_P2_INSTQUEUE_REG_12__4_,
    P2_P2_INSTQUEUE_REG_12__3_, P2_P2_INSTQUEUE_REG_12__2_,
    P2_P2_INSTQUEUE_REG_12__1_, P2_P2_INSTQUEUE_REG_12__0_,
    P2_P2_INSTQUEUE_REG_11__7_, P2_P2_INSTQUEUE_REG_11__6_,
    P2_P2_INSTQUEUE_REG_11__5_, P2_P2_INSTQUEUE_REG_11__4_,
    P2_P2_INSTQUEUE_REG_11__3_, P2_P2_INSTQUEUE_REG_11__2_,
    P2_P2_INSTQUEUE_REG_11__1_, P2_P2_INSTQUEUE_REG_11__0_,
    P2_P2_INSTQUEUE_REG_10__7_, P2_P2_INSTQUEUE_REG_10__6_,
    P2_P2_INSTQUEUE_REG_10__5_, P2_P2_INSTQUEUE_REG_10__4_,
    P2_P2_INSTQUEUE_REG_10__3_, P2_P2_INSTQUEUE_REG_10__2_,
    P2_P2_INSTQUEUE_REG_10__1_, P2_P2_INSTQUEUE_REG_10__0_,
    P2_P2_INSTQUEUE_REG_9__7_, P2_P2_INSTQUEUE_REG_9__6_,
    P2_P2_INSTQUEUE_REG_9__5_, P2_P2_INSTQUEUE_REG_9__4_,
    P2_P2_INSTQUEUE_REG_9__3_, P2_P2_INSTQUEUE_REG_9__2_,
    P2_P2_INSTQUEUE_REG_9__1_, P2_P2_INSTQUEUE_REG_9__0_,
    P2_P2_INSTQUEUE_REG_8__7_, P2_P2_INSTQUEUE_REG_8__6_,
    P2_P2_INSTQUEUE_REG_8__5_, P2_P2_INSTQUEUE_REG_8__4_,
    P2_P2_INSTQUEUE_REG_8__3_, P2_P2_INSTQUEUE_REG_8__2_,
    P2_P2_INSTQUEUE_REG_8__1_, P2_P2_INSTQUEUE_REG_8__0_,
    P2_P2_INSTQUEUE_REG_7__7_, P2_P2_INSTQUEUE_REG_7__6_,
    P2_P2_INSTQUEUE_REG_7__5_, P2_P2_INSTQUEUE_REG_7__4_,
    P2_P2_INSTQUEUE_REG_7__3_, P2_P2_INSTQUEUE_REG_7__2_,
    P2_P2_INSTQUEUE_REG_7__1_, P2_P2_INSTQUEUE_REG_7__0_,
    P2_P2_INSTQUEUE_REG_6__7_, P2_P2_INSTQUEUE_REG_6__6_,
    P2_P2_INSTQUEUE_REG_6__5_, P2_P2_INSTQUEUE_REG_6__4_,
    P2_P2_INSTQUEUE_REG_6__3_, P2_P2_INSTQUEUE_REG_6__2_,
    P2_P2_INSTQUEUE_REG_6__1_, P2_P2_INSTQUEUE_REG_6__0_,
    P2_P2_INSTQUEUE_REG_5__7_, P2_P2_INSTQUEUE_REG_5__6_,
    P2_P2_INSTQUEUE_REG_5__5_, P2_P2_INSTQUEUE_REG_5__4_,
    P2_P2_INSTQUEUE_REG_5__3_, P2_P2_INSTQUEUE_REG_5__2_,
    P2_P2_INSTQUEUE_REG_5__1_, P2_P2_INSTQUEUE_REG_5__0_,
    P2_P2_INSTQUEUE_REG_4__7_, P2_P2_INSTQUEUE_REG_4__6_,
    P2_P2_INSTQUEUE_REG_4__5_, P2_P2_INSTQUEUE_REG_4__4_,
    P2_P2_INSTQUEUE_REG_4__3_, P2_P2_INSTQUEUE_REG_4__2_,
    P2_P2_INSTQUEUE_REG_4__1_, P2_P2_INSTQUEUE_REG_4__0_,
    P2_P2_INSTQUEUE_REG_3__7_, P2_P2_INSTQUEUE_REG_3__6_,
    P2_P2_INSTQUEUE_REG_3__5_, P2_P2_INSTQUEUE_REG_3__4_,
    P2_P2_INSTQUEUE_REG_3__3_, P2_P2_INSTQUEUE_REG_3__2_,
    P2_P2_INSTQUEUE_REG_3__1_, P2_P2_INSTQUEUE_REG_3__0_,
    P2_P2_INSTQUEUE_REG_2__7_, P2_P2_INSTQUEUE_REG_2__6_,
    P2_P2_INSTQUEUE_REG_2__5_, P2_P2_INSTQUEUE_REG_2__4_,
    P2_P2_INSTQUEUE_REG_2__3_, P2_P2_INSTQUEUE_REG_2__2_,
    P2_P2_INSTQUEUE_REG_2__1_, P2_P2_INSTQUEUE_REG_2__0_,
    P2_P2_INSTQUEUE_REG_1__7_, P2_P2_INSTQUEUE_REG_1__6_,
    P2_P2_INSTQUEUE_REG_1__5_, P2_P2_INSTQUEUE_REG_1__4_,
    P2_P2_INSTQUEUE_REG_1__3_, P2_P2_INSTQUEUE_REG_1__2_,
    P2_P2_INSTQUEUE_REG_1__1_, P2_P2_INSTQUEUE_REG_1__0_,
    P2_P2_INSTQUEUE_REG_0__7_, P2_P2_INSTQUEUE_REG_0__6_,
    P2_P2_INSTQUEUE_REG_0__5_, P2_P2_INSTQUEUE_REG_0__4_,
    P2_P2_INSTQUEUE_REG_0__3_, P2_P2_INSTQUEUE_REG_0__2_,
    P2_P2_INSTQUEUE_REG_0__1_, P2_P2_INSTQUEUE_REG_0__0_,
    P2_P2_INSTQUEUERD_ADDR_REG_4_, P2_P2_INSTQUEUERD_ADDR_REG_3_,
    P2_P2_INSTQUEUERD_ADDR_REG_2_, P2_P2_INSTQUEUERD_ADDR_REG_1_,
    P2_P2_INSTQUEUERD_ADDR_REG_0_, P2_P2_INSTQUEUEWR_ADDR_REG_4_,
    P2_P2_INSTQUEUEWR_ADDR_REG_3_, P2_P2_INSTQUEUEWR_ADDR_REG_2_,
    P2_P2_INSTQUEUEWR_ADDR_REG_1_, P2_P2_INSTQUEUEWR_ADDR_REG_0_,
    P2_P2_INSTADDRPOINTER_REG_0_, P2_P2_INSTADDRPOINTER_REG_1_,
    P2_P2_INSTADDRPOINTER_REG_2_, P2_P2_INSTADDRPOINTER_REG_3_,
    P2_P2_INSTADDRPOINTER_REG_4_, P2_P2_INSTADDRPOINTER_REG_5_,
    P2_P2_INSTADDRPOINTER_REG_6_, P2_P2_INSTADDRPOINTER_REG_7_,
    P2_P2_INSTADDRPOINTER_REG_8_, P2_P2_INSTADDRPOINTER_REG_9_,
    P2_P2_INSTADDRPOINTER_REG_10_, P2_P2_INSTADDRPOINTER_REG_11_,
    P2_P2_INSTADDRPOINTER_REG_12_, P2_P2_INSTADDRPOINTER_REG_13_,
    P2_P2_INSTADDRPOINTER_REG_14_, P2_P2_INSTADDRPOINTER_REG_15_,
    P2_P2_INSTADDRPOINTER_REG_16_, P2_P2_INSTADDRPOINTER_REG_17_,
    P2_P2_INSTADDRPOINTER_REG_18_, P2_P2_INSTADDRPOINTER_REG_19_,
    P2_P2_INSTADDRPOINTER_REG_20_, P2_P2_INSTADDRPOINTER_REG_21_,
    P2_P2_INSTADDRPOINTER_REG_22_, P2_P2_INSTADDRPOINTER_REG_23_,
    P2_P2_INSTADDRPOINTER_REG_24_, P2_P2_INSTADDRPOINTER_REG_25_,
    P2_P2_INSTADDRPOINTER_REG_26_, P2_P2_INSTADDRPOINTER_REG_27_,
    P2_P2_INSTADDRPOINTER_REG_28_, P2_P2_INSTADDRPOINTER_REG_29_,
    P2_P2_INSTADDRPOINTER_REG_30_, P2_P2_INSTADDRPOINTER_REG_31_,
    P2_P2_PHYADDRPOINTER_REG_0_, P2_P2_PHYADDRPOINTER_REG_1_,
    P2_P2_PHYADDRPOINTER_REG_2_, P2_P2_PHYADDRPOINTER_REG_3_,
    P2_P2_PHYADDRPOINTER_REG_4_, P2_P2_PHYADDRPOINTER_REG_5_,
    P2_P2_PHYADDRPOINTER_REG_6_, P2_P2_PHYADDRPOINTER_REG_7_,
    P2_P2_PHYADDRPOINTER_REG_8_, P2_P2_PHYADDRPOINTER_REG_9_,
    P2_P2_PHYADDRPOINTER_REG_10_, P2_P2_PHYADDRPOINTER_REG_11_,
    P2_P2_PHYADDRPOINTER_REG_12_, P2_P2_PHYADDRPOINTER_REG_13_,
    P2_P2_PHYADDRPOINTER_REG_14_, P2_P2_PHYADDRPOINTER_REG_15_,
    P2_P2_PHYADDRPOINTER_REG_16_, P2_P2_PHYADDRPOINTER_REG_17_,
    P2_P2_PHYADDRPOINTER_REG_18_, P2_P2_PHYADDRPOINTER_REG_19_,
    P2_P2_PHYADDRPOINTER_REG_20_, P2_P2_PHYADDRPOINTER_REG_21_,
    P2_P2_PHYADDRPOINTER_REG_22_, P2_P2_PHYADDRPOINTER_REG_23_,
    P2_P2_PHYADDRPOINTER_REG_24_, P2_P2_PHYADDRPOINTER_REG_25_,
    P2_P2_PHYADDRPOINTER_REG_26_, P2_P2_PHYADDRPOINTER_REG_27_,
    P2_P2_PHYADDRPOINTER_REG_28_, P2_P2_PHYADDRPOINTER_REG_29_,
    P2_P2_PHYADDRPOINTER_REG_30_, P2_P2_PHYADDRPOINTER_REG_31_,
    P2_P2_LWORD_REG_15_, P2_P2_LWORD_REG_14_, P2_P2_LWORD_REG_13_,
    P2_P2_LWORD_REG_12_, P2_P2_LWORD_REG_11_, P2_P2_LWORD_REG_10_,
    P2_P2_LWORD_REG_9_, P2_P2_LWORD_REG_8_, P2_P2_LWORD_REG_7_,
    P2_P2_LWORD_REG_6_, P2_P2_LWORD_REG_5_, P2_P2_LWORD_REG_4_,
    P2_P2_LWORD_REG_3_, P2_P2_LWORD_REG_2_, P2_P2_LWORD_REG_1_,
    P2_P2_LWORD_REG_0_, P2_P2_UWORD_REG_14_, P2_P2_UWORD_REG_13_,
    P2_P2_UWORD_REG_12_, P2_P2_UWORD_REG_11_, P2_P2_UWORD_REG_10_,
    P2_P2_UWORD_REG_9_, P2_P2_UWORD_REG_8_, P2_P2_UWORD_REG_7_,
    P2_P2_UWORD_REG_6_, P2_P2_UWORD_REG_5_, P2_P2_UWORD_REG_4_,
    P2_P2_UWORD_REG_3_, P2_P2_UWORD_REG_2_, P2_P2_UWORD_REG_1_,
    P2_P2_UWORD_REG_0_, P2_P2_DATAO_REG_0_, P2_P2_DATAO_REG_1_,
    P2_P2_DATAO_REG_2_, P2_P2_DATAO_REG_3_, P2_P2_DATAO_REG_4_,
    P2_P2_DATAO_REG_5_, P2_P2_DATAO_REG_6_, P2_P2_DATAO_REG_7_,
    P2_P2_DATAO_REG_8_, P2_P2_DATAO_REG_9_, P2_P2_DATAO_REG_10_,
    P2_P2_DATAO_REG_11_, P2_P2_DATAO_REG_12_, P2_P2_DATAO_REG_13_,
    P2_P2_DATAO_REG_14_, P2_P2_DATAO_REG_15_, P2_P2_DATAO_REG_16_,
    P2_P2_DATAO_REG_17_, P2_P2_DATAO_REG_18_, P2_P2_DATAO_REG_19_,
    P2_P2_DATAO_REG_20_, P2_P2_DATAO_REG_21_, P2_P2_DATAO_REG_22_,
    P2_P2_DATAO_REG_23_, P2_P2_DATAO_REG_24_, P2_P2_DATAO_REG_25_,
    P2_P2_DATAO_REG_26_, P2_P2_DATAO_REG_27_, P2_P2_DATAO_REG_28_,
    P2_P2_DATAO_REG_29_, P2_P2_DATAO_REG_30_, P2_P2_DATAO_REG_31_,
    P2_P2_EAX_REG_0_, P2_P2_EAX_REG_1_, P2_P2_EAX_REG_2_, P2_P2_EAX_REG_3_,
    P2_P2_EAX_REG_4_, P2_P2_EAX_REG_5_, P2_P2_EAX_REG_6_, P2_P2_EAX_REG_7_,
    P2_P2_EAX_REG_8_, P2_P2_EAX_REG_9_, P2_P2_EAX_REG_10_,
    P2_P2_EAX_REG_11_, P2_P2_EAX_REG_12_, P2_P2_EAX_REG_13_,
    P2_P2_EAX_REG_14_, P2_P2_EAX_REG_15_, P2_P2_EAX_REG_16_,
    P2_P2_EAX_REG_17_, P2_P2_EAX_REG_18_, P2_P2_EAX_REG_19_,
    P2_P2_EAX_REG_20_, P2_P2_EAX_REG_21_, P2_P2_EAX_REG_22_,
    P2_P2_EAX_REG_23_, P2_P2_EAX_REG_24_, P2_P2_EAX_REG_25_,
    P2_P2_EAX_REG_26_, P2_P2_EAX_REG_27_, P2_P2_EAX_REG_28_,
    P2_P2_EAX_REG_29_, P2_P2_EAX_REG_30_, P2_P2_EAX_REG_31_,
    P2_P2_EBX_REG_0_, P2_P2_EBX_REG_1_, P2_P2_EBX_REG_2_, P2_P2_EBX_REG_3_,
    P2_P2_EBX_REG_4_, P2_P2_EBX_REG_5_, P2_P2_EBX_REG_6_, P2_P2_EBX_REG_7_,
    P2_P2_EBX_REG_8_, P2_P2_EBX_REG_9_, P2_P2_EBX_REG_10_,
    P2_P2_EBX_REG_11_, P2_P2_EBX_REG_12_, P2_P2_EBX_REG_13_,
    P2_P2_EBX_REG_14_, P2_P2_EBX_REG_15_, P2_P2_EBX_REG_16_,
    P2_P2_EBX_REG_17_, P2_P2_EBX_REG_18_, P2_P2_EBX_REG_19_,
    P2_P2_EBX_REG_20_, P2_P2_EBX_REG_21_, P2_P2_EBX_REG_22_,
    P2_P2_EBX_REG_23_, P2_P2_EBX_REG_24_, P2_P2_EBX_REG_25_,
    P2_P2_EBX_REG_26_, P2_P2_EBX_REG_27_, P2_P2_EBX_REG_28_,
    P2_P2_EBX_REG_29_, P2_P2_EBX_REG_30_, P2_P2_EBX_REG_31_,
    P2_P2_REIP_REG_0_, P2_P2_REIP_REG_1_, P2_P2_REIP_REG_2_,
    P2_P2_REIP_REG_3_, P2_P2_REIP_REG_4_, P2_P2_REIP_REG_5_,
    P2_P2_REIP_REG_6_, P2_P2_REIP_REG_7_, P2_P2_REIP_REG_8_,
    P2_P2_REIP_REG_9_, P2_P2_REIP_REG_10_, P2_P2_REIP_REG_11_,
    P2_P2_REIP_REG_12_, P2_P2_REIP_REG_13_, P2_P2_REIP_REG_14_,
    P2_P2_REIP_REG_15_, P2_P2_REIP_REG_16_, P2_P2_REIP_REG_17_,
    P2_P2_REIP_REG_18_, P2_P2_REIP_REG_19_, P2_P2_REIP_REG_20_,
    P2_P2_REIP_REG_21_, P2_P2_REIP_REG_22_, P2_P2_REIP_REG_23_,
    P2_P2_REIP_REG_24_, P2_P2_REIP_REG_25_, P2_P2_REIP_REG_26_,
    P2_P2_REIP_REG_27_, P2_P2_REIP_REG_28_, P2_P2_REIP_REG_29_,
    P2_P2_REIP_REG_30_, P2_P2_REIP_REG_31_, P2_P2_BYTEENABLE_REG_3_,
    P2_P2_BYTEENABLE_REG_2_, P2_P2_BYTEENABLE_REG_1_,
    P2_P2_BYTEENABLE_REG_0_, P2_P2_W_R_N_REG, P2_P2_FLUSH_REG,
    P2_P2_MORE_REG, P2_P2_STATEBS16_REG, P2_P2_REQUESTPENDING_REG,
    P2_P2_D_C_N_REG, P2_P2_M_IO_N_REG, P2_P2_CODEFETCH_REG,
    P2_P2_ADS_N_REG, P2_P2_READREQUEST_REG, P2_P2_MEMORYFETCH_REG,
    P2_P1_BE_N_REG_3_, P2_P1_BE_N_REG_2_, P2_P1_BE_N_REG_1_,
    P2_P1_BE_N_REG_0_, P2_P1_ADDRESS_REG_29_, P2_P1_ADDRESS_REG_28_,
    P2_P1_ADDRESS_REG_27_, P2_P1_ADDRESS_REG_26_, P2_P1_ADDRESS_REG_25_,
    P2_P1_ADDRESS_REG_24_, P2_P1_ADDRESS_REG_23_, P2_P1_ADDRESS_REG_22_,
    P2_P1_ADDRESS_REG_21_, P2_P1_ADDRESS_REG_20_, P2_P1_ADDRESS_REG_19_,
    P2_P1_ADDRESS_REG_18_, P2_P1_ADDRESS_REG_17_, P2_P1_ADDRESS_REG_16_,
    P2_P1_ADDRESS_REG_15_, P2_P1_ADDRESS_REG_14_, P2_P1_ADDRESS_REG_13_,
    P2_P1_ADDRESS_REG_12_, P2_P1_ADDRESS_REG_11_, P2_P1_ADDRESS_REG_10_,
    P2_P1_ADDRESS_REG_9_, P2_P1_ADDRESS_REG_8_, P2_P1_ADDRESS_REG_7_,
    P2_P1_ADDRESS_REG_6_, P2_P1_ADDRESS_REG_5_, P2_P1_ADDRESS_REG_4_,
    P2_P1_ADDRESS_REG_3_, P2_P1_ADDRESS_REG_2_, P2_P1_ADDRESS_REG_1_,
    P2_P1_ADDRESS_REG_0_, P2_P1_STATE_REG_2_, P2_P1_STATE_REG_1_,
    P2_P1_STATE_REG_0_, P2_P1_DATAWIDTH_REG_0_, P2_P1_DATAWIDTH_REG_1_,
    P2_P1_DATAWIDTH_REG_2_, P2_P1_DATAWIDTH_REG_3_, P2_P1_DATAWIDTH_REG_4_,
    P2_P1_DATAWIDTH_REG_5_, P2_P1_DATAWIDTH_REG_6_, P2_P1_DATAWIDTH_REG_7_,
    P2_P1_DATAWIDTH_REG_8_, P2_P1_DATAWIDTH_REG_9_,
    P2_P1_DATAWIDTH_REG_10_, P2_P1_DATAWIDTH_REG_11_,
    P2_P1_DATAWIDTH_REG_12_, P2_P1_DATAWIDTH_REG_13_,
    P2_P1_DATAWIDTH_REG_14_, P2_P1_DATAWIDTH_REG_15_,
    P2_P1_DATAWIDTH_REG_16_, P2_P1_DATAWIDTH_REG_17_,
    P2_P1_DATAWIDTH_REG_18_, P2_P1_DATAWIDTH_REG_19_,
    P2_P1_DATAWIDTH_REG_20_, P2_P1_DATAWIDTH_REG_21_,
    P2_P1_DATAWIDTH_REG_22_, P2_P1_DATAWIDTH_REG_23_,
    P2_P1_DATAWIDTH_REG_24_, P2_P1_DATAWIDTH_REG_25_,
    P2_P1_DATAWIDTH_REG_26_, P2_P1_DATAWIDTH_REG_27_,
    P2_P1_DATAWIDTH_REG_28_, P2_P1_DATAWIDTH_REG_29_,
    P2_P1_DATAWIDTH_REG_30_, P2_P1_DATAWIDTH_REG_31_, P2_P1_STATE2_REG_3_,
    P2_P1_STATE2_REG_2_, P2_P1_STATE2_REG_1_, P2_P1_STATE2_REG_0_,
    P2_P1_INSTQUEUE_REG_15__7_, P2_P1_INSTQUEUE_REG_15__6_,
    P2_P1_INSTQUEUE_REG_15__5_, P2_P1_INSTQUEUE_REG_15__4_,
    P2_P1_INSTQUEUE_REG_15__3_, P2_P1_INSTQUEUE_REG_15__2_,
    P2_P1_INSTQUEUE_REG_15__1_, P2_P1_INSTQUEUE_REG_15__0_,
    P2_P1_INSTQUEUE_REG_14__7_, P2_P1_INSTQUEUE_REG_14__6_,
    P2_P1_INSTQUEUE_REG_14__5_, P2_P1_INSTQUEUE_REG_14__4_,
    P2_P1_INSTQUEUE_REG_14__3_, P2_P1_INSTQUEUE_REG_14__2_,
    P2_P1_INSTQUEUE_REG_14__1_, P2_P1_INSTQUEUE_REG_14__0_,
    P2_P1_INSTQUEUE_REG_13__7_, P2_P1_INSTQUEUE_REG_13__6_,
    P2_P1_INSTQUEUE_REG_13__5_, P2_P1_INSTQUEUE_REG_13__4_,
    P2_P1_INSTQUEUE_REG_13__3_, P2_P1_INSTQUEUE_REG_13__2_,
    P2_P1_INSTQUEUE_REG_13__1_, P2_P1_INSTQUEUE_REG_13__0_,
    P2_P1_INSTQUEUE_REG_12__7_, P2_P1_INSTQUEUE_REG_12__6_,
    P2_P1_INSTQUEUE_REG_12__5_, P2_P1_INSTQUEUE_REG_12__4_,
    P2_P1_INSTQUEUE_REG_12__3_, P2_P1_INSTQUEUE_REG_12__2_,
    P2_P1_INSTQUEUE_REG_12__1_, P2_P1_INSTQUEUE_REG_12__0_,
    P2_P1_INSTQUEUE_REG_11__7_, P2_P1_INSTQUEUE_REG_11__6_,
    P2_P1_INSTQUEUE_REG_11__5_, P2_P1_INSTQUEUE_REG_11__4_,
    P2_P1_INSTQUEUE_REG_11__3_, P2_P1_INSTQUEUE_REG_11__2_,
    P2_P1_INSTQUEUE_REG_11__1_, P2_P1_INSTQUEUE_REG_11__0_,
    P2_P1_INSTQUEUE_REG_10__7_, P2_P1_INSTQUEUE_REG_10__6_,
    P2_P1_INSTQUEUE_REG_10__5_, P2_P1_INSTQUEUE_REG_10__4_,
    P2_P1_INSTQUEUE_REG_10__3_, P2_P1_INSTQUEUE_REG_10__2_,
    P2_P1_INSTQUEUE_REG_10__1_, P2_P1_INSTQUEUE_REG_10__0_,
    P2_P1_INSTQUEUE_REG_9__7_, P2_P1_INSTQUEUE_REG_9__6_,
    P2_P1_INSTQUEUE_REG_9__5_, P2_P1_INSTQUEUE_REG_9__4_,
    P2_P1_INSTQUEUE_REG_9__3_, P2_P1_INSTQUEUE_REG_9__2_,
    P2_P1_INSTQUEUE_REG_9__1_, P2_P1_INSTQUEUE_REG_9__0_,
    P2_P1_INSTQUEUE_REG_8__7_, P2_P1_INSTQUEUE_REG_8__6_,
    P2_P1_INSTQUEUE_REG_8__5_, P2_P1_INSTQUEUE_REG_8__4_,
    P2_P1_INSTQUEUE_REG_8__3_, P2_P1_INSTQUEUE_REG_8__2_,
    P2_P1_INSTQUEUE_REG_8__1_, P2_P1_INSTQUEUE_REG_8__0_,
    P2_P1_INSTQUEUE_REG_7__7_, P2_P1_INSTQUEUE_REG_7__6_,
    P2_P1_INSTQUEUE_REG_7__5_, P2_P1_INSTQUEUE_REG_7__4_,
    P2_P1_INSTQUEUE_REG_7__3_, P2_P1_INSTQUEUE_REG_7__2_,
    P2_P1_INSTQUEUE_REG_7__1_, P2_P1_INSTQUEUE_REG_7__0_,
    P2_P1_INSTQUEUE_REG_6__7_, P2_P1_INSTQUEUE_REG_6__6_,
    P2_P1_INSTQUEUE_REG_6__5_, P2_P1_INSTQUEUE_REG_6__4_,
    P2_P1_INSTQUEUE_REG_6__3_, P2_P1_INSTQUEUE_REG_6__2_,
    P2_P1_INSTQUEUE_REG_6__1_, P2_P1_INSTQUEUE_REG_6__0_,
    P2_P1_INSTQUEUE_REG_5__7_, P2_P1_INSTQUEUE_REG_5__6_,
    P2_P1_INSTQUEUE_REG_5__5_, P2_P1_INSTQUEUE_REG_5__4_,
    P2_P1_INSTQUEUE_REG_5__3_, P2_P1_INSTQUEUE_REG_5__2_,
    P2_P1_INSTQUEUE_REG_5__1_, P2_P1_INSTQUEUE_REG_5__0_,
    P2_P1_INSTQUEUE_REG_4__7_, P2_P1_INSTQUEUE_REG_4__6_,
    P2_P1_INSTQUEUE_REG_4__5_, P2_P1_INSTQUEUE_REG_4__4_,
    P2_P1_INSTQUEUE_REG_4__3_, P2_P1_INSTQUEUE_REG_4__2_,
    P2_P1_INSTQUEUE_REG_4__1_, P2_P1_INSTQUEUE_REG_4__0_,
    P2_P1_INSTQUEUE_REG_3__7_, P2_P1_INSTQUEUE_REG_3__6_,
    P2_P1_INSTQUEUE_REG_3__5_, P2_P1_INSTQUEUE_REG_3__4_,
    P2_P1_INSTQUEUE_REG_3__3_, P2_P1_INSTQUEUE_REG_3__2_,
    P2_P1_INSTQUEUE_REG_3__1_, P2_P1_INSTQUEUE_REG_3__0_,
    P2_P1_INSTQUEUE_REG_2__7_, P2_P1_INSTQUEUE_REG_2__6_,
    P2_P1_INSTQUEUE_REG_2__5_, P2_P1_INSTQUEUE_REG_2__4_,
    P2_P1_INSTQUEUE_REG_2__3_, P2_P1_INSTQUEUE_REG_2__2_,
    P2_P1_INSTQUEUE_REG_2__1_, P2_P1_INSTQUEUE_REG_2__0_,
    P2_P1_INSTQUEUE_REG_1__7_, P2_P1_INSTQUEUE_REG_1__6_,
    P2_P1_INSTQUEUE_REG_1__5_, P2_P1_INSTQUEUE_REG_1__4_,
    P2_P1_INSTQUEUE_REG_1__3_, P2_P1_INSTQUEUE_REG_1__2_,
    P2_P1_INSTQUEUE_REG_1__1_, P2_P1_INSTQUEUE_REG_1__0_,
    P2_P1_INSTQUEUE_REG_0__7_, P2_P1_INSTQUEUE_REG_0__6_,
    P2_P1_INSTQUEUE_REG_0__5_, P2_P1_INSTQUEUE_REG_0__4_,
    P2_P1_INSTQUEUE_REG_0__3_, P2_P1_INSTQUEUE_REG_0__2_,
    P2_P1_INSTQUEUE_REG_0__1_, P2_P1_INSTQUEUE_REG_0__0_,
    P2_P1_INSTQUEUERD_ADDR_REG_4_, P2_P1_INSTQUEUERD_ADDR_REG_3_,
    P2_P1_INSTQUEUERD_ADDR_REG_2_, P2_P1_INSTQUEUERD_ADDR_REG_1_,
    P2_P1_INSTQUEUERD_ADDR_REG_0_, P2_P1_INSTQUEUEWR_ADDR_REG_4_,
    P2_P1_INSTQUEUEWR_ADDR_REG_3_, P2_P1_INSTQUEUEWR_ADDR_REG_2_,
    P2_P1_INSTQUEUEWR_ADDR_REG_1_, P2_P1_INSTQUEUEWR_ADDR_REG_0_,
    P2_P1_INSTADDRPOINTER_REG_0_, P2_P1_INSTADDRPOINTER_REG_1_,
    P2_P1_INSTADDRPOINTER_REG_2_, P2_P1_INSTADDRPOINTER_REG_3_,
    P2_P1_INSTADDRPOINTER_REG_4_, P2_P1_INSTADDRPOINTER_REG_5_,
    P2_P1_INSTADDRPOINTER_REG_6_, P2_P1_INSTADDRPOINTER_REG_7_,
    P2_P1_INSTADDRPOINTER_REG_8_, P2_P1_INSTADDRPOINTER_REG_9_,
    P2_P1_INSTADDRPOINTER_REG_10_, P2_P1_INSTADDRPOINTER_REG_11_,
    P2_P1_INSTADDRPOINTER_REG_12_, P2_P1_INSTADDRPOINTER_REG_13_,
    P2_P1_INSTADDRPOINTER_REG_14_, P2_P1_INSTADDRPOINTER_REG_15_,
    P2_P1_INSTADDRPOINTER_REG_16_, P2_P1_INSTADDRPOINTER_REG_17_,
    P2_P1_INSTADDRPOINTER_REG_18_, P2_P1_INSTADDRPOINTER_REG_19_,
    P2_P1_INSTADDRPOINTER_REG_20_, P2_P1_INSTADDRPOINTER_REG_21_,
    P2_P1_INSTADDRPOINTER_REG_22_, P2_P1_INSTADDRPOINTER_REG_23_,
    P2_P1_INSTADDRPOINTER_REG_24_, P2_P1_INSTADDRPOINTER_REG_25_,
    P2_P1_INSTADDRPOINTER_REG_26_, P2_P1_INSTADDRPOINTER_REG_27_,
    P2_P1_INSTADDRPOINTER_REG_28_, P2_P1_INSTADDRPOINTER_REG_29_,
    P2_P1_INSTADDRPOINTER_REG_30_, P2_P1_INSTADDRPOINTER_REG_31_,
    P2_P1_PHYADDRPOINTER_REG_0_, P2_P1_PHYADDRPOINTER_REG_1_,
    P2_P1_PHYADDRPOINTER_REG_2_, P2_P1_PHYADDRPOINTER_REG_3_,
    P2_P1_PHYADDRPOINTER_REG_4_, P2_P1_PHYADDRPOINTER_REG_5_,
    P2_P1_PHYADDRPOINTER_REG_6_, P2_P1_PHYADDRPOINTER_REG_7_,
    P2_P1_PHYADDRPOINTER_REG_8_, P2_P1_PHYADDRPOINTER_REG_9_,
    P2_P1_PHYADDRPOINTER_REG_10_, P2_P1_PHYADDRPOINTER_REG_11_,
    P2_P1_PHYADDRPOINTER_REG_12_, P2_P1_PHYADDRPOINTER_REG_13_,
    P2_P1_PHYADDRPOINTER_REG_14_, P2_P1_PHYADDRPOINTER_REG_15_,
    P2_P1_PHYADDRPOINTER_REG_16_, P2_P1_PHYADDRPOINTER_REG_17_,
    P2_P1_PHYADDRPOINTER_REG_18_, P2_P1_PHYADDRPOINTER_REG_19_,
    P2_P1_PHYADDRPOINTER_REG_20_, P2_P1_PHYADDRPOINTER_REG_21_,
    P2_P1_PHYADDRPOINTER_REG_22_, P2_P1_PHYADDRPOINTER_REG_23_,
    P2_P1_PHYADDRPOINTER_REG_24_, P2_P1_PHYADDRPOINTER_REG_25_,
    P2_P1_PHYADDRPOINTER_REG_26_, P2_P1_PHYADDRPOINTER_REG_27_,
    P2_P1_PHYADDRPOINTER_REG_28_, P2_P1_PHYADDRPOINTER_REG_29_,
    P2_P1_PHYADDRPOINTER_REG_30_, P2_P1_PHYADDRPOINTER_REG_31_,
    P2_P1_LWORD_REG_15_, P2_P1_LWORD_REG_14_, P2_P1_LWORD_REG_13_,
    P2_P1_LWORD_REG_12_, P2_P1_LWORD_REG_11_, P2_P1_LWORD_REG_10_,
    P2_P1_LWORD_REG_9_, P2_P1_LWORD_REG_8_, P2_P1_LWORD_REG_7_,
    P2_P1_LWORD_REG_6_, P2_P1_LWORD_REG_5_, P2_P1_LWORD_REG_4_,
    P2_P1_LWORD_REG_3_, P2_P1_LWORD_REG_2_, P2_P1_LWORD_REG_1_,
    P2_P1_LWORD_REG_0_, P2_P1_UWORD_REG_14_, P2_P1_UWORD_REG_13_,
    P2_P1_UWORD_REG_12_, P2_P1_UWORD_REG_11_, P2_P1_UWORD_REG_10_,
    P2_P1_UWORD_REG_9_, P2_P1_UWORD_REG_8_, P2_P1_UWORD_REG_7_,
    P2_P1_UWORD_REG_6_, P2_P1_UWORD_REG_5_, P2_P1_UWORD_REG_4_,
    P2_P1_UWORD_REG_3_, P2_P1_UWORD_REG_2_, P2_P1_UWORD_REG_1_,
    P2_P1_UWORD_REG_0_, P2_P1_DATAO_REG_0_, P2_P1_DATAO_REG_1_,
    P2_P1_DATAO_REG_2_, P2_P1_DATAO_REG_3_, P2_P1_DATAO_REG_4_,
    P2_P1_DATAO_REG_5_, P2_P1_DATAO_REG_6_, P2_P1_DATAO_REG_7_,
    P2_P1_DATAO_REG_8_, P2_P1_DATAO_REG_9_, P2_P1_DATAO_REG_10_,
    P2_P1_DATAO_REG_11_, P2_P1_DATAO_REG_12_, P2_P1_DATAO_REG_13_,
    P2_P1_DATAO_REG_14_, P2_P1_DATAO_REG_15_, P2_P1_DATAO_REG_16_,
    P2_P1_DATAO_REG_17_, P2_P1_DATAO_REG_18_, P2_P1_DATAO_REG_19_,
    P2_P1_DATAO_REG_20_, P2_P1_DATAO_REG_21_, P2_P1_DATAO_REG_22_,
    P2_P1_DATAO_REG_23_, P2_P1_DATAO_REG_24_, P2_P1_DATAO_REG_25_,
    P2_P1_DATAO_REG_26_, P2_P1_DATAO_REG_27_, P2_P1_DATAO_REG_28_,
    P2_P1_DATAO_REG_29_, P2_P1_DATAO_REG_30_, P2_P1_DATAO_REG_31_,
    P2_P1_EAX_REG_0_, P2_P1_EAX_REG_1_, P2_P1_EAX_REG_2_, P2_P1_EAX_REG_3_,
    P2_P1_EAX_REG_4_, P2_P1_EAX_REG_5_, P2_P1_EAX_REG_6_, P2_P1_EAX_REG_7_,
    P2_P1_EAX_REG_8_, P2_P1_EAX_REG_9_, P2_P1_EAX_REG_10_,
    P2_P1_EAX_REG_11_, P2_P1_EAX_REG_12_, P2_P1_EAX_REG_13_,
    P2_P1_EAX_REG_14_, P2_P1_EAX_REG_15_, P2_P1_EAX_REG_16_,
    P2_P1_EAX_REG_17_, P2_P1_EAX_REG_18_, P2_P1_EAX_REG_19_,
    P2_P1_EAX_REG_20_, P2_P1_EAX_REG_21_, P2_P1_EAX_REG_22_,
    P2_P1_EAX_REG_23_, P2_P1_EAX_REG_24_, P2_P1_EAX_REG_25_,
    P2_P1_EAX_REG_26_, P2_P1_EAX_REG_27_, P2_P1_EAX_REG_28_,
    P2_P1_EAX_REG_29_, P2_P1_EAX_REG_30_, P2_P1_EAX_REG_31_,
    P2_P1_EBX_REG_0_, P2_P1_EBX_REG_1_, P2_P1_EBX_REG_2_, P2_P1_EBX_REG_3_,
    P2_P1_EBX_REG_4_, P2_P1_EBX_REG_5_, P2_P1_EBX_REG_6_, P2_P1_EBX_REG_7_,
    P2_P1_EBX_REG_8_, P2_P1_EBX_REG_9_, P2_P1_EBX_REG_10_,
    P2_P1_EBX_REG_11_, P2_P1_EBX_REG_12_, P2_P1_EBX_REG_13_,
    P2_P1_EBX_REG_14_, P2_P1_EBX_REG_15_, P2_P1_EBX_REG_16_,
    P2_P1_EBX_REG_17_, P2_P1_EBX_REG_18_, P2_P1_EBX_REG_19_,
    P2_P1_EBX_REG_20_, P2_P1_EBX_REG_21_, P2_P1_EBX_REG_22_,
    P2_P1_EBX_REG_23_, P2_P1_EBX_REG_24_, P2_P1_EBX_REG_25_,
    P2_P1_EBX_REG_26_, P2_P1_EBX_REG_27_, P2_P1_EBX_REG_28_,
    P2_P1_EBX_REG_29_, P2_P1_EBX_REG_30_, P2_P1_EBX_REG_31_,
    P2_P1_REIP_REG_0_, P2_P1_REIP_REG_1_, P2_P1_REIP_REG_2_,
    P2_P1_REIP_REG_3_, P2_P1_REIP_REG_4_, P2_P1_REIP_REG_5_,
    P2_P1_REIP_REG_6_, P2_P1_REIP_REG_7_, P2_P1_REIP_REG_8_,
    P2_P1_REIP_REG_9_, P2_P1_REIP_REG_10_, P2_P1_REIP_REG_11_,
    P2_P1_REIP_REG_12_, P2_P1_REIP_REG_13_, P2_P1_REIP_REG_14_,
    P2_P1_REIP_REG_15_, P2_P1_REIP_REG_16_, P2_P1_REIP_REG_17_,
    P2_P1_REIP_REG_18_, P2_P1_REIP_REG_19_, P2_P1_REIP_REG_20_,
    P2_P1_REIP_REG_21_, P2_P1_REIP_REG_22_, P2_P1_REIP_REG_23_,
    P2_P1_REIP_REG_24_, P2_P1_REIP_REG_25_, P2_P1_REIP_REG_26_,
    P2_P1_REIP_REG_27_, P2_P1_REIP_REG_28_, P2_P1_REIP_REG_29_,
    P2_P1_REIP_REG_30_, P2_P1_REIP_REG_31_, P2_P1_BYTEENABLE_REG_3_,
    P2_P1_BYTEENABLE_REG_2_, P2_P1_BYTEENABLE_REG_1_,
    P2_P1_BYTEENABLE_REG_0_, P2_P1_W_R_N_REG, P2_P1_FLUSH_REG,
    P2_P1_MORE_REG, P2_P1_STATEBS16_REG, P2_P1_REQUESTPENDING_REG,
    P2_P1_D_C_N_REG, P2_P1_M_IO_N_REG, P2_P1_CODEFETCH_REG,
    P2_P1_ADS_N_REG, P2_P1_READREQUEST_REG, P2_P1_MEMORYFETCH_REG;
  wire n10021_1, n10022, n10023, n10024, n10025, n10026_1, n10027, n10028,
    n10029, n10030, n10031_1, n10032, n10033, n10034, n10035, n10036_1,
    n10037, n10038, n10039, n10040, n10041_1, n10042, n10043, n10044,
    n10045, n10046_1, n10047, n10048, n10049, n10050, n10051_1, n10052,
    n10053, n10054, n10055, n10056_1, n10057, n10058, n10059, n10060,
    n10061_1, n10062, n10063, n10064, n10065, n10066_1, n10067, n10068,
    n10069, n10070, n10071_1, n10072, n10073, n10074, n10075, n10076_1,
    n10077, n10078, n10079, n10080, n10081_1, n10082, n10083, n10084,
    n10085, n10086_1, n10087, n10088, n10089, n10090, n10091_1, n10092,
    n10093, n10094, n10095, n10096_1, n10097, n10098, n10099, n10100,
    n10101_1, n10102, n10103, n10104, n10105, n10106_1, n10107, n10108,
    n10109, n10110, n10111_1, n10112, n10113, n10114, n10115, n10116_1,
    n10117, n10118, n10119, n10120, n10121_1, n10122, n10123, n10124,
    n10125, n10126_1, n10127, n10128, n10129, n10130, n10131_1, n10132,
    n10133, n10134, n10135, n10136_1, n10137, n10138, n10139, n10140,
    n10141_1, n10142, n10143, n10144, n10145, n10146_1, n10147, n10148,
    n10149, n10150, n10151_1, n10152, n10153, n10154, n10155, n10156_1,
    n10157, n10158, n10159, n10160, n10161_1, n10162, n10163, n10164,
    n10165, n10166_1, n10167, n10168, n10169, n10170, n10171_1, n10172,
    n10173, n10174, n10175, n10176_1, n10177, n10178, n10179, n10180,
    n10181_1, n10182, n10183, n10184, n10185, n10186_1, n10187, n10188,
    n10189, n10190, n10191_1, n10192, n10193, n10194, n10195, n10196_1,
    n10197, n10198, n10199, n10200, n10201_1, n10202, n10203, n10204,
    n10205, n10206_1, n10207, n10208, n10209, n10210, n10211_1, n10212,
    n10213, n10214, n10215, n10216_1, n10217, n10218, n10219, n10220,
    n10221_1, n10222, n10223, n10224, n10225, n10226_1, n10227, n10228,
    n10229, n10230, n10231_1, n10232, n10233, n10234, n10235, n10236_1,
    n10237, n10238, n10239, n10240, n10241_1, n10242, n10243, n10244,
    n10245, n10246_1, n10247, n10248, n10249, n10250, n10251_1, n10252,
    n10253, n10254, n10255, n10256_1, n10257, n10258, n10259, n10260,
    n10261_1, n10262, n10263, n10264, n10265, n10266_1, n10267, n10268,
    n10269, n10270, n10271_1, n10272, n10273, n10274, n10275, n10276_1,
    n10277, n10278, n10279, n10280, n10281_1, n10282, n10283, n10284,
    n10285, n10286_1, n10287, n10288, n10289, n10290, n10291_1, n10292,
    n10293, n10294, n10295, n10296_1, n10297, n10298, n10299, n10300,
    n10301_1, n10302, n10303, n10304, n10305, n10306_1, n10307, n10308,
    n10309, n10310, n10311_1, n10312, n10313, n10314, n10315, n10316_1,
    n10317, n10318, n10319, n10320, n10321_1, n10322, n10323, n10324,
    n10325, n10326_1, n10327, n10328, n10329, n10330, n10331_1, n10332,
    n10333, n10334, n10335, n10336_1, n10337, n10338, n10339, n10340,
    n10341_1, n10342, n10343, n10344, n10345, n10346_1, n10347, n10348,
    n10349, n10350, n10351_1, n10352, n10353, n10354, n10355, n10356_1,
    n10357, n10358, n10359, n10360, n10361_1, n10362, n10363, n10364,
    n10365, n10366_1, n10367, n10368, n10369, n10370, n10371_1, n10372,
    n10373, n10374, n10375, n10376_1, n10377, n10378, n10379, n10380,
    n10381_1, n10382, n10383, n10384, n10385, n10386_1, n10387, n10388,
    n10389, n10390, n10391_1, n10392, n10393, n10394, n10395, n10396_1,
    n10397, n10398, n10399, n10400, n10401_1, n10402, n10403, n10404,
    n10405, n10406_1, n10407, n10408, n10409, n10410, n10411_1, n10412,
    n10413, n10414, n10415, n10416_1, n10417, n10418, n10419, n10420,
    n10421_1, n10422, n10423, n10424, n10425, n10426_1, n10427, n10428,
    n10429, n10430, n10431_1, n10432, n10433, n10434, n10435, n10436_1,
    n10437, n10438, n10439, n10440, n10441_1, n10442, n10443, n10444,
    n10445, n10446_1, n10447, n10448, n10449, n10450, n10451_1, n10452,
    n10453, n10454, n10455, n10456_1, n10457, n10458, n10459, n10460,
    n10461_1, n10462, n10463, n10464, n10465, n10466_1, n10467, n10468,
    n10469, n10470, n10471_1, n10472, n10473, n10474, n10475, n10476_1,
    n10477, n10478, n10479, n10480, n10481_1, n10482, n10483, n10484,
    n10485, n10486_1, n10487, n10488, n10489, n10490, n10491_1, n10492,
    n10493, n10494, n10495, n10496_1, n10497, n10498, n10499, n10500,
    n10501_1, n10502, n10503, n10504, n10505, n10506_1, n10507, n10508,
    n10509, n10510, n10511_1, n10512, n10513, n10514, n10515, n10516_1,
    n10517, n10518, n10519, n10520, n10521_1, n10522, n10523, n10524,
    n10525, n10526_1, n10527, n10528, n10529, n10530, n10531_1, n10532,
    n10533, n10534, n10535, n10536_1, n10537, n10538, n10539, n10540,
    n10541_1, n10542, n10543, n10544, n10545, n10546_1, n10547, n10548,
    n10549, n10550, n10551_1, n10552, n10553, n10554, n10555, n10556_1,
    n10557, n10558, n10559, n10560, n10561_1, n10562, n10563, n10564,
    n10565, n10566_1, n10567, n10568, n10569, n10570, n10571_1, n10572,
    n10573, n10574, n10575, n10576_1, n10577, n10578, n10579, n10580,
    n10581_1, n10582, n10583, n10584, n10585, n10586_1, n10587, n10588,
    n10589, n10590, n10591_1, n10592, n10593, n10594, n10595, n10596_1,
    n10597, n10598, n10599, n10600, n10601_1, n10602, n10603, n10604,
    n10605, n10606_1, n10607, n10608, n10609, n10610, n10611_1, n10612,
    n10613, n10614, n10615, n10616_1, n10617, n10618, n10619, n10620,
    n10621_1, n10622, n10623, n10624, n10625, n10626_1, n10627, n10628,
    n10629, n10630, n10631_1, n10632, n10633, n10634, n10635, n10636_1,
    n10637, n10638, n10639, n10640, n10641_1, n10642, n10643, n10644,
    n10645, n10646_1, n10647, n10648, n10649, n10650, n10651_1, n10652,
    n10653, n10654, n10655, n10656_1, n10657, n10658, n10659, n10660,
    n10661_1, n10662, n10663, n10664, n10665, n10666_1, n10667, n10668,
    n10669, n10670, n10671_1, n10672, n10673, n10674, n10675, n10676_1,
    n10677, n10678, n10679, n10680, n10681_1, n10682, n10683, n10684,
    n10685, n10686_1, n10687, n10688, n10689, n10690, n10691_1, n10692,
    n10693, n10694, n10695, n10696_1, n10697, n10698, n10699, n10700,
    n10701_1, n10702, n10703, n10704, n10705, n10706_1, n10707, n10708,
    n10709, n10710, n10711_1, n10712, n10713, n10714, n10715, n10716_1,
    n10717, n10718, n10719, n10720, n10721_1, n10722, n10723, n10724,
    n10725, n10726_1, n10727, n10728, n10729, n10730, n10731_1, n10732,
    n10733, n10734, n10735, n10736_1, n10737, n10738, n10739, n10740,
    n10741_1, n10742, n10743, n10744, n10745, n10746_1, n10747, n10748,
    n10749, n10750, n10751_1, n10752, n10753, n10754, n10755, n10756_1,
    n10757, n10758, n10759, n10760, n10761_1, n10762, n10763, n10764,
    n10765, n10766_1, n10767, n10768, n10769, n10770, n10771_1, n10772,
    n10773, n10774, n10775, n10776_1, n10777, n10778, n10779, n10780,
    n10781_1, n10782, n10783, n10784, n10785, n10786_1, n10787, n10788,
    n10789, n10790, n10791_1, n10792, n10793, n10794, n10795, n10796_1,
    n10797, n10798, n10799, n10800, n10801_1, n10802, n10803, n10804,
    n10805, n10806_1, n10807, n10808, n10809, n10810, n10811_1, n10812,
    n10813, n10814, n10815, n10816_1, n10817, n10818, n10819, n10820,
    n10821_1, n10822, n10823, n10824, n10825, n10826_1, n10827, n10828,
    n10829, n10830, n10831_1, n10832, n10833, n10834, n10835, n10836_1,
    n10837, n10838, n10839, n10840, n10841_1, n10842, n10843, n10844,
    n10845, n10846_1, n10847, n10848, n10849, n10850, n10851_1, n10852,
    n10853, n10854, n10855, n10856_1, n10857, n10858, n10859, n10860,
    n10861_1, n10862, n10863, n10864, n10865, n10866_1, n10867, n10868,
    n10869, n10870, n10871_1, n10872, n10873, n10874, n10875, n10876_1,
    n10877, n10878, n10879, n10880, n10881_1, n10882, n10883, n10884,
    n10885, n10886_1, n10887, n10888, n10889, n10890, n10891_1, n10892,
    n10893, n10894, n10895, n10896_1, n10897, n10898, n10899, n10900,
    n10901_1, n10902, n10903, n10904, n10905, n10906_1, n10907, n10908,
    n10909, n10910, n10911_1, n10912, n10913, n10914, n10915, n10916_1,
    n10917, n10918, n10919, n10920, n10921_1, n10922, n10923, n10924,
    n10925, n10926_1, n10927, n10928, n10929, n10930, n10931_1, n10932,
    n10933, n10934, n10935, n10936_1, n10937, n10938, n10939, n10940,
    n10941_1, n10942, n10943, n10944, n10945, n10946_1, n10947, n10948,
    n10949, n10950, n10951_1, n10952, n10953, n10954, n10955, n10956_1,
    n10957, n10958, n10959, n10960, n10961_1, n10962, n10963, n10964,
    n10965, n10966_1, n10967, n10968, n10969, n10970, n10971_1, n10972,
    n10973, n10974, n10975, n10976_1, n10977, n10978, n10979, n10980,
    n10981_1, n10982, n10983, n10984, n10985, n10986_1, n10987, n10988,
    n10989, n10990, n10991_1, n10992, n10993, n10994, n10995, n10996_1,
    n10997, n10998, n10999, n11000, n11001_1, n11002, n11003, n11004,
    n11005, n11006_1, n11007, n11008, n11009, n11010, n11011_1, n11012,
    n11013, n11014, n11015, n11016_1, n11017, n11018, n11019, n11020,
    n11021_1, n11022, n11023, n11024, n11025, n11026_1, n11027, n11028,
    n11029, n11030, n11031_1, n11032, n11033, n11034, n11035, n11036_1,
    n11037, n11038, n11039, n11040, n11041_1, n11042, n11043, n11044,
    n11045, n11046_1, n11047, n11048, n11049, n11050, n11051_1, n11052,
    n11053, n11054, n11055, n11056_1, n11057, n11058, n11059, n11060,
    n11061_1, n11062, n11063, n11064, n11065, n11066_1, n11067, n11068,
    n11069, n11070, n11071_1, n11072, n11073, n11074, n11075, n11076_1,
    n11077, n11078, n11079, n11080, n11081_1, n11082, n11083, n11084,
    n11085, n11086_1, n11087, n11088, n11089, n11090, n11091_1, n11092,
    n11093, n11094, n11095, n11096_1, n11097, n11098, n11099, n11100,
    n11101_1, n11102, n11103, n11104, n11105, n11106_1, n11107, n11108,
    n11109, n11110, n11111_1, n11112, n11113, n11114, n11115, n11116_1,
    n11117, n11118, n11119, n11120, n11121_1, n11122, n11123, n11124,
    n11125, n11126_1, n11127, n11128, n11129, n11130, n11131_1, n11132,
    n11133, n11134, n11135, n11136_1, n11137, n11138, n11139, n11140,
    n11141_1, n11142, n11143, n11144, n11145, n11146_1, n11147, n11148,
    n11149, n11150, n11151_1, n11152, n11153, n11154, n11155, n11156_1,
    n11157, n11158, n11159, n11160, n11161_1, n11162, n11163, n11164,
    n11165, n11166_1, n11167, n11168, n11169, n11170, n11171_1, n11172,
    n11173, n11174, n11175, n11176_1, n11177, n11178, n11179, n11180,
    n11181_1, n11182, n11183, n11184, n11185, n11186_1, n11187, n11188,
    n11189, n11190, n11191_1, n11192, n11193, n11194, n11195, n11196_1,
    n11197, n11198, n11199, n11200, n11201_1, n11202, n11203, n11204,
    n11205, n11206_1, n11207, n11208, n11209, n11210, n11211_1, n11212,
    n11213, n11214, n11215, n11216_1, n11217, n11218, n11219, n11220,
    n11221_1, n11222, n11223, n11224, n11225, n11226_1, n11227, n11228,
    n11229, n11230, n11231_1, n11232, n11233, n11234, n11235, n11236_1,
    n11237, n11238, n11239, n11240, n11241_1, n11242, n11243, n11244,
    n11245, n11246_1, n11247, n11248, n11249, n11250, n11251_1, n11252,
    n11253, n11254, n11255, n11256_1, n11257, n11258, n11259, n11260,
    n11261_1, n11262, n11263, n11264, n11265, n11266_1, n11267, n11268,
    n11269, n11270, n11271_1, n11272, n11273, n11274, n11275, n11276_1,
    n11277, n11278, n11279, n11280, n11281_1, n11282, n11283, n11284,
    n11285, n11286_1, n11287, n11288, n11289, n11290, n11291_1, n11292,
    n11293, n11294, n11295, n11296_1, n11297, n11298, n11299, n11300,
    n11301_1, n11302, n11303, n11304, n11305, n11306_1, n11307, n11308,
    n11309, n11310, n11311_1, n11312, n11313, n11314, n11315, n11316_1,
    n11317, n11318, n11319, n11320, n11321_1, n11322, n11323, n11324,
    n11325, n11326_1, n11327, n11328, n11329, n11330, n11331_1, n11332,
    n11333, n11334, n11335, n11336_1, n11337, n11338, n11339, n11340,
    n11341_1, n11342, n11343, n11344, n11345, n11346_1, n11347, n11348,
    n11349, n11350, n11351_1, n11352, n11353, n11354, n11355, n11356_1,
    n11357, n11358, n11359, n11360, n11361_1, n11362, n11363, n11364,
    n11365, n11366_1, n11367, n11368, n11369, n11370, n11371_1, n11372,
    n11373, n11374, n11375, n11376_1, n11377, n11378, n11379, n11380,
    n11381_1, n11382, n11383, n11384, n11385, n11386_1, n11387, n11388,
    n11389, n11390, n11391_1, n11392, n11393, n11394, n11395, n11396_1,
    n11397, n11398, n11399, n11400, n11401_1, n11402, n11403, n11404,
    n11405, n11406_1, n11407, n11408, n11409, n11410, n11411_1, n11412,
    n11413, n11414, n11415, n11416_1, n11417, n11418, n11419, n11420,
    n11421_1, n11422, n11423, n11424, n11425, n11426_1, n11427, n11428,
    n11429, n11430, n11431_1, n11432, n11433, n11434, n11435, n11436_1,
    n11437, n11438, n11439, n11440, n11441_1, n11442, n11443, n11444,
    n11445, n11446_1, n11447, n11448, n11449, n11450, n11451_1, n11452,
    n11453, n11454, n11455, n11456_1, n11457, n11458, n11459, n11460,
    n11461_1, n11462, n11463, n11464, n11465, n11466_1, n11467, n11468,
    n11469, n11470, n11471_1, n11472, n11473, n11474, n11475, n11476_1,
    n11477, n11478, n11479, n11480, n11481_1, n11482, n11483, n11484,
    n11485, n11486_1, n11487, n11488, n11489, n11490, n11491_1, n11492,
    n11493, n11494, n11495, n11496_1, n11497, n11498, n11499, n11500,
    n11501_1, n11502, n11503, n11504, n11505, n11506_1, n11507, n11508,
    n11509, n11510, n11511_1, n11512, n11513, n11514, n11515, n11516_1,
    n11517, n11518, n11519, n11520, n11521_1, n11522, n11523, n11524,
    n11525, n11526_1, n11527, n11528, n11529, n11530, n11531_1, n11532,
    n11533, n11534, n11535, n11536_1, n11537, n11538, n11539, n11540,
    n11541_1, n11542, n11543, n11544, n11545, n11546_1, n11547, n11548,
    n11549, n11550, n11551_1, n11552, n11553, n11554, n11555, n11556_1,
    n11557, n11558, n11559, n11560, n11561_1, n11562, n11563, n11564,
    n11565, n11566_1, n11567, n11568, n11569, n11570, n11571_1, n11572,
    n11573, n11574, n11575, n11576_1, n11577, n11578, n11579, n11580,
    n11581_1, n11582, n11583, n11584, n11585, n11586_1, n11587, n11588,
    n11589, n11590, n11591_1, n11592, n11593, n11594, n11595, n11596_1,
    n11597, n11598, n11599, n11600, n11601_1, n11602, n11603, n11604,
    n11605, n11606_1, n11607, n11608, n11609, n11610, n11611_1, n11612,
    n11613, n11614, n11615, n11616_1, n11617, n11618, n11619, n11620,
    n11621_1, n11622, n11623, n11624, n11625, n11626_1, n11627, n11628,
    n11629, n11630, n11631_1, n11632, n11633, n11634, n11635, n11636_1,
    n11637, n11638, n11639, n11640, n11641_1, n11642, n11643, n11644,
    n11645, n11646_1, n11647, n11648, n11649, n11650, n11651_1, n11652,
    n11653, n11654, n11655, n11656_1, n11657, n11658, n11659, n11660,
    n11661_1, n11662, n11663, n11664, n11665, n11666_1, n11667, n11668,
    n11669, n11670, n11671_1, n11672, n11673, n11674, n11675, n11676_1,
    n11677, n11678, n11679, n11680, n11681_1, n11682, n11683, n11684,
    n11685, n11686_1, n11687, n11688, n11689, n11690, n11691_1, n11692,
    n11693, n11694, n11695, n11696_1, n11697, n11698, n11699, n11700,
    n11701_1, n11702, n11703, n11704, n11705, n11706_1, n11707, n11708,
    n11709, n11710, n11711_1, n11712, n11713, n11714, n11715, n11716_1,
    n11717, n11718, n11719, n11720, n11721_1, n11722, n11723, n11724,
    n11725, n11726_1, n11727, n11728, n11729, n11730, n11731_1, n11732,
    n11733, n11734, n11735, n11736_1, n11737, n11738, n11739, n11740,
    n11741_1, n11742, n11743, n11744, n11745, n11746_1, n11747, n11748,
    n11749, n11750, n11751_1, n11752, n11753, n11754, n11755, n11756_1,
    n11757, n11758, n11759, n11760, n11761_1, n11762, n11763, n11764,
    n11765, n11766_1, n11767, n11768, n11769, n11770, n11771_1, n11772,
    n11773, n11774, n11775, n11776_1, n11777, n11778, n11779, n11780,
    n11781_1, n11782, n11783, n11784, n11785, n11786_1, n11787, n11788,
    n11789, n11790, n11791_1, n11792, n11793, n11794, n11795, n11796_1,
    n11797, n11798, n11799, n11800, n11801_1, n11802, n11803, n11804,
    n11805, n11806_1, n11807, n11808, n11809, n11810, n11811_1, n11812,
    n11813, n11814, n11815, n11816_1, n11817, n11818, n11819, n11820,
    n11821_1, n11822, n11823, n11824, n11825, n11826_1, n11827, n11828,
    n11829, n11830, n11831_1, n11832, n11833, n11834, n11835, n11836_1,
    n11837, n11838, n11839, n11840, n11841_1, n11842, n11843, n11844,
    n11845, n11846_1, n11847, n11848, n11849, n11850, n11851_1, n11852,
    n11853, n11854, n11855, n11856_1, n11857, n11858, n11859, n11860,
    n11861_1, n11862, n11863, n11864, n11865, n11866_1, n11867, n11868,
    n11869, n11870, n11871_1, n11872, n11873, n11874, n11875, n11876_1,
    n11877, n11878, n11879, n11880, n11881_1, n11882, n11883, n11884,
    n11885, n11886_1, n11887, n11888, n11889, n11890, n11891_1, n11892,
    n11893, n11894, n11895, n11896_1, n11897, n11898, n11899, n11900,
    n11901_1, n11902, n11903, n11904, n11905, n11906_1, n11907, n11908,
    n11909, n11910, n11911_1, n11912, n11913, n11914, n11915, n11916_1,
    n11917, n11918, n11919, n11920, n11921_1, n11922, n11923, n11924,
    n11925, n11926_1, n11927, n11928, n11929, n11930, n11931_1, n11932,
    n11933, n11934, n11935, n11936_1, n11937, n11938, n11939, n11940,
    n11941_1, n11942, n11943, n11944, n11945, n11946_1, n11947, n11948,
    n11949, n11950, n11951_1, n11952, n11953, n11954, n11955, n11956_1,
    n11957, n11958, n11959, n11960, n11961_1, n11962, n11963, n11964,
    n11965, n11966_1, n11967, n11968, n11969, n11970, n11971_1, n11972,
    n11973, n11974, n11975, n11976_1, n11977, n11978, n11979, n11980,
    n11981_1, n11982, n11983, n11984, n11985, n11986_1, n11987, n11988,
    n11989, n11990, n11991_1, n11992, n11993, n11994, n11995, n11996_1,
    n11997, n11998, n11999, n12000, n12001_1, n12002, n12003, n12004,
    n12005, n12006_1, n12007, n12008, n12009, n12010, n12011_1, n12012,
    n12013, n12014, n12015, n12016_1, n12017, n12018, n12019, n12020,
    n12021_1, n12022, n12023, n12024, n12025, n12026_1, n12027, n12028,
    n12029, n12030, n12031_1, n12032, n12033, n12034, n12035, n12036_1,
    n12037, n12038, n12039, n12040, n12041_1, n12042, n12043, n12044,
    n12045, n12046_1, n12047, n12048, n12049, n12050, n12051_1, n12052,
    n12053, n12054, n12055, n12056_1, n12057, n12058, n12059, n12060,
    n12061_1, n12062, n12063, n12064, n12065, n12066_1, n12067, n12068,
    n12069, n12070, n12071_1, n12072, n12073, n12074, n12075, n12076_1,
    n12077, n12078, n12079, n12080, n12081_1, n12082, n12083, n12084,
    n12085, n12086_1, n12087, n12088, n12089, n12090, n12091_1, n12092,
    n12093, n12094, n12095, n12096_1, n12097, n12098, n12099, n12100,
    n12101_1, n12102, n12103, n12104, n12105, n12106_1, n12107, n12108,
    n12109, n12110, n12111_1, n12112, n12113, n12114, n12115, n12116_1,
    n12117, n12118, n12119, n12120, n12121_1, n12122, n12123, n12124,
    n12125, n12126_1, n12127, n12128, n12129, n12130, n12131_1, n12132,
    n12133, n12134, n12135, n12136_1, n12137, n12138, n12139, n12140,
    n12141_1, n12142, n12143, n12144, n12145, n12146_1, n12147, n12148,
    n12149, n12150, n12151_1, n12152, n12154, n12155, n12156_1, n12157,
    n12158, n12159, n12160, n12161_1, n12162, n12163, n12164, n12165,
    n12166_1, n12167, n12168, n12169, n12170, n12171_1, n12172, n12173,
    n12174, n12175, n12176_1, n12177, n12178, n12179, n12180, n12181_1,
    n12182, n12183, n12184, n12185, n12186_1, n12187, n12188, n12189,
    n12190, n12191_1, n12192, n12193, n12194, n12195, n12196_1, n12197,
    n12198, n12199, n12200, n12201_1, n12202, n12203, n12204, n12205,
    n12206_1, n12207, n12208, n12209, n12210, n12211_1, n12212, n12213,
    n12214, n12215, n12216_1, n12217, n12218, n12219, n12220, n12221_1,
    n12222, n12223, n12224, n12225, n12226_1, n12227, n12228, n12229,
    n12230, n12231_1, n12232, n12233, n12234, n12235, n12236_1, n12237,
    n12238, n12239, n12240, n12241_1, n12242, n12243, n12244, n12245,
    n12246_1, n12247, n12248, n12249, n12250, n12251_1, n12252, n12253,
    n12254, n12255, n12256_1, n12257, n12258, n12259, n12260, n12261_1,
    n12262, n12263, n12264, n12265, n12266_1, n12267, n12268, n12269,
    n12270, n12271_1, n12272, n12273, n12274, n12275, n12276_1, n12277,
    n12278, n12280, n12281_1, n12282, n12284, n12285, n12286_1, n12287,
    n12288, n12289, n12290, n12291_1, n12293, n12294, n12295, n12296_1,
    n12297, n12298, n12300, n12301_1, n12302, n12303, n12304, n12305,
    n12306_1, n12307, n12309, n12310, n12311_1, n12312, n12313, n12314,
    n12316_1, n12317, n12318, n12319, n12320, n12321_1, n12322, n12324,
    n12325, n12326_1, n12327, n12328, n12329, n12331_1, n12332, n12333,
    n12334, n12335, n12336_1, n12337, n12338, n12340, n12341_1, n12342,
    n12344, n12345, n12346_1, n12347, n12348, n12349, n12350, n12351_1,
    n12353, n12354, n12355, n12356_1, n12357, n12358, n12360, n12361_1,
    n12362, n12363, n12364, n12365, n12366_1, n12368, n12369, n12370,
    n12372, n12373, n12374, n12375, n12376_1, n12377, n12378, n12379,
    n12381_1, n12382, n12383, n12384, n12385, n12386_1, n12388, n12389,
    n12390, n12391_1, n12392, n12393, n12394, n12396_1, n12397, n12398,
    n12399, n12400, n12401_1, n12404, n12405, n12406_1, n12407, n12408,
    n12409, n12410, n12411_1, n12412, n12413, n12414, n12415, n12416_1,
    n12417, n12418, n12419, n12420, n12421_1, n12423, n12424, n12425,
    n12426_1, n12428, n12429, n12430, n12431_1, n12432, n12433, n12434,
    n12435, n12436_1, n12437, n12438, n12439, n12440, n12441_1, n12442,
    n12443, n12444, n12445, n12446_1, n12447, n12448, n12449, n12450,
    n12451_1, n12452, n12453, n12454, n12455, n12456_1, n12457, n12458,
    n12459, n12460, n12461_1, n12462, n12463, n12465, n12466_1, n12467,
    n12468, n12469, n12470, n12471_1, n12472, n12473, n12474, n12475,
    n12476_1, n12477, n12478, n12479, n12480, n12481_1, n12482, n12483,
    n12484, n12485, n12486_1, n12487, n12488, n12489, n12490, n12491_1,
    n12492, n12493, n12494, n12495, n12496_1, n12497, n12498, n12499,
    n12500, n12501_1, n12502, n12503, n12504, n12505, n12506_1, n12507,
    n12509, n12510, n12511_1, n12512, n12514, n12515, n12516_1, n12517,
    n12519, n12520, n12521_1, n12522, n12524, n12525, n12526_1, n12527,
    n12529, n12530, n12531_1, n12532, n12534, n12535, n12536_1, n12537,
    n12539, n12540, n12541_1, n12542, n12544, n12545, n12546_1, n12547,
    n12549, n12550, n12551_1, n12552, n12554, n12555, n12556_1, n12557,
    n12559, n12560, n12561_1, n12562, n12564, n12565, n12566_1, n12567,
    n12569, n12570, n12571_1, n12572, n12574, n12575, n12576_1, n12577,
    n12579, n12580, n12581_1, n12582, n12584, n12585, n12586_1, n12587,
    n12589, n12590, n12591_1, n12592, n12594, n12595, n12596_1, n12597,
    n12599, n12600, n12601_1, n12602, n12604, n12605, n12606_1, n12607,
    n12609, n12610, n12611_1, n12612, n12614, n12615, n12616_1, n12617,
    n12619, n12620, n12621_1, n12622, n12624, n12625, n12626_1, n12627,
    n12629, n12630, n12631_1, n12632, n12634, n12635, n12636_1, n12637,
    n12639, n12640, n12641_1, n12642, n12644, n12645, n12646_1, n12647,
    n12649, n12650, n12651_1, n12652, n12654, n12655, n12656_1, n12657,
    n12659, n12660, n12661_1, n12662, n12665, n12666_1, n12668, n12669,
    n12671_1, n12672, n12674, n12675, n12677, n12678, n12680, n12681_1,
    n12683, n12684, n12686_1, n12687, n12689, n12690, n12692, n12693,
    n12695, n12696_1, n12698, n12699, n12701_1, n12702, n12704, n12705,
    n12707, n12708, n12710, n12711_1, n12713, n12714, n12716_1, n12717,
    n12719, n12720, n12722, n12723, n12725, n12726_1, n12728, n12729,
    n12731_1, n12732, n12734, n12735, n12737, n12738, n12740, n12741_1,
    n12743, n12744, n12746_1, n12747, n12749, n12750, n12752, n12753,
    n12755, n12756_1, n12758, n12759, n12762, n12763, n12764, n12765,
    n12766_1, n12767, n12768, n12770, n12771_1, n12772, n12773, n12774,
    n12775, n12776_1, n12777, n12778, n12779, n12780, n12781_1, n12782,
    n12783, n12784, n12785, n12786_1, n12787, n12788, n12789, n12790,
    n12791_1, n12792, n12793, n12794, n12795, n12796_1, n12797, n12798,
    n12799, n12800, n12801_1, n12802, n12803, n12804, n12805, n12807,
    n12808, n12809, n12810, n12811_1, n12812, n12813, n12814, n12815,
    n12816_1, n12817, n12818, n12819, n12820, n12821_1, n12822, n12823,
    n12824, n12825, n12826_1, n12827, n12828, n12829, n12830, n12831_1,
    n12832, n12833, n12834, n12835, n12836_1, n12837, n12838, n12839,
    n12840, n12841_1, n12842, n12843, n12844, n12845, n12846_1, n12847,
    n12848, n12849, n12851_1, n12852, n12853, n12854, n12856_1, n12857,
    n12858, n12859, n12861_1, n12862, n12863, n12864, n12866_1, n12867,
    n12868, n12869, n12871_1, n12872, n12873, n12874, n12876_1, n12877,
    n12878, n12879, n12881_1, n12882, n12883, n12884, n12886_1, n12887,
    n12888, n12889, n12891_1, n12892, n12893, n12894, n12896_1, n12897,
    n12898, n12899, n12901_1, n12902, n12903, n12904, n12906_1, n12907,
    n12908, n12909, n12911_1, n12912, n12913, n12914, n12916_1, n12917,
    n12918, n12919, n12921_1, n12922, n12923, n12924, n12926_1, n12927,
    n12928, n12929, n12931_1, n12932, n12933, n12934, n12936_1, n12937,
    n12938, n12939, n12941_1, n12942, n12943, n12944, n12946_1, n12947,
    n12948, n12949, n12951_1, n12952, n12953, n12954, n12956_1, n12957,
    n12958, n12959, n12961_1, n12962, n12963, n12964, n12966_1, n12967,
    n12968, n12969, n12971_1, n12972, n12973, n12974, n12976_1, n12977,
    n12978, n12979, n12981_1, n12982, n12983, n12984, n12986_1, n12987,
    n12988, n12989, n12991_1, n12992, n12993, n12994, n12996_1, n12997,
    n12998, n12999, n13001_1, n13002, n13003, n13004, n13007, n13008,
    n13010, n13011_1, n13013, n13014, n13016_1, n13017, n13019, n13020,
    n13022, n13023, n13025, n13026_1, n13028, n13029, n13031_1, n13032,
    n13034, n13035, n13037, n13038, n13040, n13041_1, n13043, n13044,
    n13046_1, n13047, n13049, n13050, n13052, n13053, n13055, n13056_1,
    n13058, n13059, n13061_1, n13062, n13064, n13065, n13067, n13068,
    n13070, n13071_1, n13073, n13074, n13076_1, n13077, n13079, n13080,
    n13082, n13083, n13085, n13086_1, n13088, n13089, n13091_1, n13092,
    n13094, n13095, n13097, n13098, n13100, n13101_1, n13104, n13105,
    n13106_1, n13107, n13108, n13109, n13110, n13112, n13113, n13114,
    n13115, n13116_1, n13117, n13119, n13120, n13121_1, n13122, n13123,
    n13124, n13125, n13127, n13128, n13129, n13130, n13131_1, n13132,
    n13133, n13134, n13136_1, n13137, n13138, n13139, n13140, n13141_1,
    n13142, n13144, n13145, n13146_1, n13147, n13148, n13149, n13150,
    n13151_1, n13153, n13154, n13155, n13156_1, n13157, n13158, n13159,
    n13161_1, n13162, n13163, n13164, n13165, n13166_1, n13167, n13168,
    n13170, n13171_1, n13172, n13173, n13174, n13175, n13176_1, n13178,
    n13179, n13180, n13181_1, n13182, n13183, n13184, n13185, n13186_1,
    n13187, n13188, n13190, n13191_1, n13192, n13193, n13194, n13195,
    n13196_1, n13198, n13199, n13200, n13201_1, n13202, n13203, n13204,
    n13205, n13207, n13208, n13209, n13210, n13211_1, n13212, n13213,
    n13215, n13216_1, n13217, n13218, n13219, n13220, n13221_1, n13222,
    n13223, n13224, n13226_1, n13227, n13228, n13229, n13230, n13231_1,
    n13232, n13234, n13235, n13236_1, n13237, n13238, n13239, n13240,
    n13241_1, n13243, n13244, n13245, n13246_1, n13247, n13248, n13249,
    n13251_1, n13252, n13253, n13254, n13255, n13256_1, n13257, n13258,
    n13259, n13260, n13261_1, n13262, n13263, n13264, n13265, n13266_1,
    n13267, n13268, n13269, n13270, n13271_1, n13273, n13274, n13275,
    n13276_1, n13277, n13278, n13279, n13281_1, n13282, n13283, n13284,
    n13285, n13286_1, n13287, n13288, n13289, n13290, n13291_1, n13292,
    n13293, n13294, n13295, n13296_1, n13297, n13299, n13300, n13301_1,
    n13302, n13303, n13304, n13305, n13306_1, n13307, n13308, n13309,
    n13310, n13311_1, n13312, n13313, n13314, n13315, n13316_1, n13317,
    n13318, n13320, n13321_1, n13322, n13323, n13324, n13325, n13326_1,
    n13327, n13328, n13329, n13330, n13331_1, n13332, n13333, n13334,
    n13335, n13336_1, n13337, n13338, n13339, n13341_1, n13342, n13343,
    n13344, n13345, n13346_1, n13348, n13349, n13350, n13351_1, n13352,
    n13353, n13354, n13355, n13356_1, n13357, n13358, n13359, n13360,
    n13361_1, n13362, n13363, n13364, n13365, n13366_1, n13368, n13369,
    n13370, n13371_1, n13372, n13373, n13374, n13375, n13376_1, n13377,
    n13378, n13379, n13380, n13381_1, n13382, n13383, n13384, n13385,
    n13386_1, n13387, n13388, n13389, n13390, n13391_1, n13393, n13394,
    n13395, n13396_1, n13397, n13398, n13399, n13400, n13401_1, n13402,
    n13403, n13404, n13405, n13406_1, n13407, n13408, n13409, n13410,
    n13411_1, n13412, n13413, n13414, n13416_1, n13417, n13418, n13419,
    n13420, n13421_1, n13423, n13424, n13425, n13426_1, n13427, n13428,
    n13429, n13430, n13431_1, n13432, n13433, n13434, n13435, n13436_1,
    n13437, n13438, n13439, n13440, n13441_1, n13442, n13443, n13444,
    n13445, n13446_1, n13447, n13449, n13450, n13451_1, n13452, n13453,
    n13454, n13456_1, n13457, n13458, n13459, n13460, n13461_1, n13462,
    n13463, n13464, n13465, n13466_1, n13467, n13468, n13469, n13470,
    n13471_1, n13472, n13473, n13474, n13475, n13476_1, n13477, n13478,
    n13479, n13480, n13481_1, n13482, n13484, n13485, n13486_1, n13487,
    n13488, n13489, n13490, n13491_1, n13492, n13493, n13494, n13496_1,
    n13497, n13498, n13499, n13500, n13501_1, n13503, n13504, n13505,
    n13506_1, n13507, n13508, n13510, n13511_1, n13512, n13513, n13514,
    n13515, n13516_1, n13517, n13518, n13519, n13520, n13521_1, n13522,
    n13523, n13524, n13525, n13526_1, n13527, n13528, n13529, n13530,
    n13531_1, n13532, n13533, n13534, n13535, n13537, n13538, n13539,
    n13571_1, n13572, n13573, n13574, n13575, n13576_1, n13577, n13578,
    n13579, n13580, n13581_1, n13582, n13583, n13584, n13585, n13586_1,
    n13587, n13588, n13589, n13590, n13591_1, n13592, n13593, n13594,
    n13595, n13596_1, n13597, n13598, n13599, n13600, n13601_1, n13602,
    n13603, n13604, n13605, n13606_1, n13607, n13608, n13609, n13610,
    n13611_1, n13612, n13613, n13614, n13615, n13616_1, n13617, n13618,
    n13619, n13620, n13621_1, n13622, n13623, n13624, n13625, n13626_1,
    n13627, n13628, n13629, n13630, n13631_1, n13632, n13633, n13634,
    n13635, n13636_1, n13637, n13638, n13639, n13640, n13641_1, n13642,
    n13643, n13644, n13645, n13646_1, n13647, n13648, n13649, n13650,
    n13651_1, n13652, n13653, n13654, n13655, n13656_1, n13657, n13658,
    n13659, n13660, n13661_1, n13662, n13663, n13664, n13665, n13666_1,
    n13667, n13668, n13669, n13670, n13671_1, n13672, n13673, n13674,
    n13675, n13676_1, n13677, n13678, n13679, n13680, n13681_1, n13682,
    n13683, n13684, n13685, n13686_1, n13687, n13688, n13689, n13690,
    n13691_1, n13692, n13693, n13694, n13695, n13696_1, n13697, n13698,
    n13699, n13700, n13701_1, n13702, n13703, n13704, n13705, n13706_1,
    n13707, n13708, n13709, n13710, n13711_1, n13712, n13713, n13714,
    n13715, n13716_1, n13717, n13718, n13719, n13720, n13721_1, n13722,
    n13723, n13724, n13725, n13726_1, n13727, n13728, n13729, n13730,
    n13731_1, n13732, n13733, n13734, n13735, n13736_1, n13737, n13738,
    n13739, n13740, n13741_1, n13742, n13744, n13745, n13746_1, n13747,
    n13748, n13749, n13750, n13751_1, n13752, n13753, n13754, n13755,
    n13756_1, n13757, n13758, n13759, n13760, n13761_1, n13762, n13763,
    n13764, n13765, n13766_1, n13767, n13768, n13769, n13770, n13771_1,
    n13772, n13773, n13774, n13775, n13776_1, n13777, n13778, n13779,
    n13780, n13781_1, n13782, n13783, n13784, n13785, n13786_1, n13787,
    n13788, n13789, n13790, n13791_1, n13792, n13793, n13794, n13795,
    n13796_1, n13797, n13798, n13800, n13801_1, n13802, n13803, n13804,
    n13805, n13806_1, n13807, n13808, n13809, n13810, n13811_1, n13812,
    n13813, n13814, n13815, n13816_1, n13817, n13818, n13819, n13820,
    n13821_1, n13822, n13823, n13824, n13825, n13826_1, n13827, n13828,
    n13829, n13830, n13831_1, n13832, n13833, n13834, n13835, n13836_1,
    n13837, n13838, n13839, n13840, n13841_1, n13842, n13843, n13844,
    n13845, n13846_1, n13847, n13848, n13849, n13850, n13851_1, n13852,
    n13853, n13854, n13855, n13856_1, n13857, n13858, n13859, n13860,
    n13862, n13863, n13864, n13865, n13866_1, n13867, n13868, n13869,
    n13870, n13871_1, n13872, n13873, n13874, n13875, n13876_1, n13877,
    n13878, n13879, n13880, n13881_1, n13882, n13883, n13884, n13885,
    n13886_1, n13887, n13888, n13889, n13890, n13891_1, n13892, n13893,
    n13894, n13895, n13896_1, n13897, n13898, n13899, n13900, n13901_1,
    n13902, n13903, n13904, n13905, n13906_1, n13907, n13908, n13909,
    n13910, n13911_1, n13912, n13913, n13914, n13915, n13916_1, n13917,
    n13918, n13919, n13920, n13921_1, n13922, n13923, n13924, n13925,
    n13927, n13928, n13929, n13930, n13931_1, n13932, n13933, n13934,
    n13935, n13936_1, n13937, n13938, n13939, n13940, n13941_1, n13942,
    n13943, n13944, n13945, n13946_1, n13947, n13948, n13949, n13950,
    n13951_1, n13952, n13953, n13954, n13955, n13956_1, n13957, n13958,
    n13959, n13960, n13961_1, n13962, n13963, n13964, n13965, n13966_1,
    n13967, n13968, n13969, n13970, n13971_1, n13972, n13973, n13974,
    n13975, n13976_1, n13977, n13978, n13979, n13980, n13981_1, n13982,
    n13983, n13984, n13985, n13986_1, n13987, n13988, n13989, n13990,
    n13991_1, n13992, n13993, n13994, n13995, n13997, n13998, n13999,
    n14000, n14001_1, n14002, n14003, n14004, n14005, n14006_1, n14007,
    n14008, n14009, n14010, n14011_1, n14012, n14013, n14014, n14015,
    n14016_1, n14017, n14018, n14019, n14020, n14021_1, n14022, n14023,
    n14024, n14025, n14026_1, n14027, n14028, n14029, n14030, n14031_1,
    n14032, n14033, n14034, n14035, n14036_1, n14037, n14038, n14039,
    n14040, n14041_1, n14042, n14043, n14044, n14045, n14046_1, n14047,
    n14048, n14049, n14050, n14051_1, n14052, n14053, n14054, n14055,
    n14056_1, n14057, n14058, n14059, n14061_1, n14062, n14063, n14064,
    n14065, n14066_1, n14067, n14068, n14069, n14070, n14071_1, n14072,
    n14073, n14074, n14075, n14076_1, n14077, n14078, n14079, n14080,
    n14081_1, n14082, n14083, n14084, n14085, n14086_1, n14087, n14088,
    n14089, n14090, n14091_1, n14092, n14093, n14094, n14095, n14096_1,
    n14097, n14098, n14099, n14100, n14101_1, n14102, n14103, n14104,
    n14105, n14106_1, n14107, n14108, n14109, n14110, n14111_1, n14112,
    n14113, n14114, n14115, n14116_1, n14117, n14118, n14119, n14120,
    n14121_1, n14122, n14123, n14124, n14125, n14126_1, n14127, n14128,
    n14129, n14130, n14131_1, n14132, n14134, n14135, n14136_1, n14137,
    n14138, n14139, n14140, n14141_1, n14142, n14143, n14144, n14145,
    n14146_1, n14147, n14148, n14149, n14150, n14151_1, n14152, n14153,
    n14154, n14155, n14156_1, n14157, n14158, n14159, n14160, n14161_1,
    n14162, n14163, n14164, n14165, n14166_1, n14167, n14168, n14169,
    n14170, n14171_1, n14172, n14173, n14174, n14175, n14176_1, n14177,
    n14178, n14179, n14180, n14181_1, n14182, n14183, n14184, n14185,
    n14186_1, n14187, n14188, n14189, n14190, n14191_1, n14192, n14193,
    n14194, n14195, n14196_1, n14197, n14198, n14199, n14200, n14201_1,
    n14203, n14204, n14205, n14206_1, n14207, n14208, n14209, n14210,
    n14211_1, n14212, n14213, n14214, n14215, n14216_1, n14217, n14218,
    n14219, n14220, n14221_1, n14222, n14223, n14224, n14225, n14226_1,
    n14227, n14228, n14229, n14230, n14231_1, n14232, n14233, n14234,
    n14235, n14236_1, n14237, n14238, n14239, n14240, n14241_1, n14242,
    n14243, n14244, n14245, n14246_1, n14247, n14248, n14249, n14250,
    n14251_1, n14252, n14253, n14254, n14255, n14256_1, n14257, n14258,
    n14259, n14260, n14261_1, n14262, n14263, n14264, n14265, n14266_1,
    n14267, n14268, n14269, n14271_1, n14272, n14273, n14274, n14275,
    n14276_1, n14277, n14278, n14279, n14280, n14281_1, n14282, n14283,
    n14284, n14285, n14286_1, n14287, n14288, n14289, n14290, n14291_1,
    n14292, n14293, n14294, n14295, n14296_1, n14297, n14298, n14299,
    n14300, n14301_1, n14302, n14303, n14304, n14305, n14306_1, n14307,
    n14308, n14309, n14310, n14311_1, n14312, n14313, n14314, n14315,
    n14316_1, n14317, n14318, n14319, n14320, n14321_1, n14322, n14323,
    n14324, n14325, n14326_1, n14327, n14328, n14329, n14330, n14331_1,
    n14332, n14333, n14334, n14335, n14336_1, n14338, n14339, n14340,
    n14341_1, n14342, n14343, n14344, n14345, n14346_1, n14347, n14348,
    n14349, n14350, n14351_1, n14352, n14353, n14354, n14355, n14356_1,
    n14357, n14358, n14359, n14360, n14361_1, n14362, n14363, n14364,
    n14365, n14366_1, n14367, n14368, n14369, n14370, n14371_1, n14372,
    n14373, n14374, n14375, n14376_1, n14377, n14378, n14379, n14380,
    n14381_1, n14382, n14383, n14384, n14385, n14386_1, n14387, n14388,
    n14389, n14390, n14391_1, n14392, n14393, n14394, n14395, n14396_1,
    n14397, n14398, n14399, n14400, n14402, n14403, n14404, n14405,
    n14406_1, n14407, n14408, n14409, n14410, n14411_1, n14412, n14413,
    n14414, n14415, n14416_1, n14417, n14418, n14419, n14420, n14421_1,
    n14422, n14423, n14424, n14425, n14426_1, n14427, n14428, n14429,
    n14430, n14431_1, n14432, n14433, n14434, n14435, n14436_1, n14437,
    n14438, n14439, n14440, n14441_1, n14442, n14443, n14444, n14445,
    n14446_1, n14447, n14448, n14449, n14450, n14451_1, n14452, n14453,
    n14454, n14455, n14456_1, n14457, n14458, n14459, n14460, n14461_1,
    n14462, n14463, n14464, n14465, n14466_1, n14467, n14468, n14469,
    n14470, n14472, n14473, n14474, n14475, n14476_1, n14477, n14478,
    n14479, n14480, n14481_1, n14482, n14483, n14484, n14485, n14486_1,
    n14487, n14488, n14489, n14490, n14491_1, n14492, n14493, n14494,
    n14495, n14496_1, n14497, n14498, n14499, n14500, n14501_1, n14502,
    n14503, n14504, n14505, n14506_1, n14507, n14508, n14509, n14510,
    n14511_1, n14512, n14513, n14514, n14515, n14516_1, n14517, n14518,
    n14519, n14520, n14521_1, n14522, n14523, n14524, n14525, n14526_1,
    n14527, n14528, n14529, n14530, n14531_1, n14532, n14533, n14534,
    n14535, n14536_1, n14538, n14539, n14540, n14541_1, n14542, n14543,
    n14544, n14545, n14546_1, n14547, n14548, n14549, n14550, n14551_1,
    n14552, n14553, n14554, n14555, n14556_1, n14557, n14558, n14559,
    n14560, n14561_1, n14562, n14563, n14564, n14565, n14566_1, n14567,
    n14568, n14569, n14570, n14571_1, n14572, n14573, n14574, n14575,
    n14576_1, n14577, n14578, n14579, n14580, n14581_1, n14582, n14583,
    n14584, n14585, n14586_1, n14587, n14588, n14589, n14590, n14591_1,
    n14592, n14593, n14594, n14595, n14596_1, n14597, n14598, n14599,
    n14600, n14602, n14603, n14604, n14605, n14606_1, n14607, n14608,
    n14609, n14610, n14611_1, n14612, n14613, n14614, n14615, n14616_1,
    n14617, n14618, n14619, n14620, n14621_1, n14622, n14623, n14624,
    n14625, n14626_1, n14627, n14628, n14629, n14630, n14631_1, n14632,
    n14633, n14634, n14635, n14636_1, n14637, n14638, n14639, n14640,
    n14641_1, n14642, n14643, n14644, n14645, n14646_1, n14647, n14648,
    n14649, n14650, n14651_1, n14652, n14653, n14654, n14655, n14656_1,
    n14657, n14658, n14659, n14660, n14661_1, n14662, n14663, n14665,
    n14666_1, n14667, n14668, n14669, n14670, n14671_1, n14672, n14673,
    n14674, n14675, n14676_1, n14677, n14678, n14679, n14680, n14681_1,
    n14682, n14683, n14684, n14685, n14686_1, n14687, n14688, n14689,
    n14690, n14691_1, n14692, n14693, n14694, n14695, n14696_1, n14697,
    n14698, n14699, n14700, n14701_1, n14702, n14703, n14704, n14705,
    n14706_1, n14707, n14708, n14709, n14710, n14711_1, n14712, n14713,
    n14714, n14715, n14716_1, n14717, n14718, n14719, n14720, n14721_1,
    n14722, n14723, n14724, n14726_1, n14727, n14728, n14729, n14730,
    n14731_1, n14732, n14733, n14734, n14735, n14736_1, n14737, n14738,
    n14739, n14740, n14741_1, n14742, n14743, n14744, n14745, n14746_1,
    n14747, n14748, n14749, n14750, n14751_1, n14752, n14753, n14754,
    n14755, n14756_1, n14757, n14758, n14759, n14760, n14761_1, n14762,
    n14763, n14764, n14765, n14766_1, n14767, n14768, n14769, n14770,
    n14771_1, n14772, n14773, n14774, n14775, n14776_1, n14777, n14778,
    n14779, n14780, n14781_1, n14782, n14783, n14784, n14785, n14786_1,
    n14787, n14788, n14789, n14790, n14791_1, n14793, n14794, n14795,
    n14796_1, n14797, n14798, n14799, n14800, n14801_1, n14802, n14803,
    n14804, n14805, n14806_1, n14807, n14808, n14809, n14810, n14811_1,
    n14812, n14813, n14814, n14815, n14816_1, n14817, n14818, n14819,
    n14820, n14821_1, n14822, n14823, n14824, n14825, n14826_1, n14827,
    n14828, n14829, n14830, n14831_1, n14832, n14833, n14834, n14835,
    n14836_1, n14837, n14838, n14839, n14840, n14841_1, n14842, n14843,
    n14844, n14845, n14846_1, n14847, n14848, n14849, n14850, n14851_1,
    n14852, n14853, n14854, n14855, n14856_1, n14857, n14858, n14859,
    n14861_1, n14862, n14863, n14864, n14865, n14866_1, n14867, n14868,
    n14869, n14870, n14871_1, n14872, n14873, n14874, n14875, n14876_1,
    n14877, n14878, n14879, n14880, n14881_1, n14882, n14883, n14884,
    n14885, n14886_1, n14887, n14888, n14889, n14890, n14891_1, n14892,
    n14893, n14894, n14895, n14896_1, n14897, n14898, n14899, n14900,
    n14901_1, n14902, n14903, n14904, n14905, n14906_1, n14907, n14908,
    n14909, n14910, n14911_1, n14912, n14913, n14914, n14915, n14916_1,
    n14917, n14918, n14919, n14920, n14921_1, n14922, n14923, n14924,
    n14925, n14927, n14928, n14929, n14930, n14931_1, n14932, n14933,
    n14934, n14935, n14936_1, n14937, n14938, n14939, n14940, n14941_1,
    n14942, n14943, n14944, n14945, n14946_1, n14947, n14948, n14949,
    n14950, n14951_1, n14952, n14953, n14954, n14955, n14956_1, n14957,
    n14958, n14959, n14960, n14961_1, n14962, n14963, n14964, n14965,
    n14966_1, n14967, n14968, n14969, n14970, n14971_1, n14972, n14973,
    n14974, n14975, n14976_1, n14977, n14978, n14979, n14980, n14981_1,
    n14982, n14983, n14984, n14985, n14986_1, n14988, n14989, n14990,
    n14991_1, n14992, n14993, n14994, n14995, n14996_1, n14997, n14998,
    n14999, n15000, n15001_1, n15002, n15003, n15004, n15005, n15006_1,
    n15007, n15008, n15009, n15010, n15011_1, n15012, n15013, n15014,
    n15015, n15016_1, n15017, n15018, n15019, n15020, n15021_1, n15022,
    n15023, n15024, n15025, n15026_1, n15027, n15028, n15029, n15030,
    n15031_1, n15032, n15033, n15034, n15035, n15036_1, n15037, n15038,
    n15039, n15040, n15041_1, n15042, n15043, n15044, n15045, n15047,
    n15048, n15049, n15050, n15051_1, n15052, n15053, n15054, n15055,
    n15056_1, n15057, n15058, n15059, n15060, n15061_1, n15062, n15063,
    n15064, n15065, n15066_1, n15067, n15068, n15069, n15070, n15071_1,
    n15072, n15073, n15074, n15075, n15076_1, n15077, n15078, n15079,
    n15080, n15081_1, n15082, n15083, n15084, n15085, n15086_1, n15087,
    n15088, n15089, n15090, n15091_1, n15092, n15093, n15094, n15095,
    n15096_1, n15097, n15098, n15099, n15100, n15101_1, n15102, n15104,
    n15105, n15106_1, n15107, n15108, n15109, n15110, n15111_1, n15112,
    n15113, n15114, n15115, n15116_1, n15117, n15118, n15119, n15120,
    n15121_1, n15122, n15123, n15124, n15125, n15126_1, n15127, n15128,
    n15129, n15130, n15131_1, n15132, n15133, n15134, n15135, n15136_1,
    n15137, n15138, n15139, n15140, n15141_1, n15142, n15143, n15144,
    n15145, n15146_1, n15147, n15148, n15149, n15150, n15151_1, n15152,
    n15153, n15154, n15155, n15156_1, n15157, n15158, n15159, n15160,
    n15161_1, n15162, n15164, n15165, n15166_1, n15167, n15168, n15169,
    n15170, n15171_1, n15172, n15173, n15174, n15175, n15176_1, n15177,
    n15178, n15179, n15180, n15181_1, n15182, n15183, n15184, n15185,
    n15186_1, n15187, n15188, n15189, n15190, n15191_1, n15192, n15193,
    n15194, n15195, n15196_1, n15197, n15198, n15199, n15200, n15201_1,
    n15202, n15203, n15204, n15205, n15206_1, n15207, n15208, n15209,
    n15210, n15211_1, n15212, n15213, n15214, n15215, n15216_1, n15217,
    n15218, n15219, n15221_1, n15222, n15223, n15224, n15225, n15226_1,
    n15227, n15228, n15229, n15230, n15231_1, n15232, n15233, n15234,
    n15235, n15236_1, n15237, n15238, n15239, n15240, n15241_1, n15242,
    n15243, n15244, n15245, n15246_1, n15247, n15248, n15249, n15250,
    n15251_1, n15252, n15253, n15254, n15255, n15256_1, n15257, n15258,
    n15259, n15260, n15261_1, n15262, n15263, n15264, n15265, n15266_1,
    n15267, n15268, n15269, n15270, n15271_1, n15272, n15273, n15274,
    n15275, n15276_1, n15277, n15278, n15279, n15280, n15281_1, n15283,
    n15284, n15285, n15286_1, n15287, n15288, n15289, n15290, n15291_1,
    n15292, n15293, n15294, n15295, n15296_1, n15297, n15298, n15299,
    n15300, n15301_1, n15302, n15303, n15304, n15305, n15306_1, n15307,
    n15308, n15309, n15310, n15311_1, n15312, n15313, n15314, n15315,
    n15316_1, n15317, n15318, n15319, n15320, n15321_1, n15322, n15323,
    n15324, n15325, n15326_1, n15327, n15328, n15329, n15330, n15331_1,
    n15332, n15333, n15334, n15335, n15336_1, n15338, n15339, n15340,
    n15341_1, n15342, n15343, n15344, n15345, n15346_1, n15347, n15348,
    n15349, n15350, n15351_1, n15352, n15353, n15354, n15355, n15356_1,
    n15357, n15358, n15359, n15360, n15361_1, n15362, n15363, n15364,
    n15365, n15366_1, n15367, n15368, n15369, n15370, n15371_1, n15372,
    n15373, n15374, n15375, n15376_1, n15377, n15378, n15379, n15380,
    n15381_1, n15382, n15383, n15384, n15385, n15386_1, n15387, n15388,
    n15389, n15390, n15391_1, n15392, n15393, n15394, n15396_1, n15397,
    n15398, n15399, n15400, n15401_1, n15402, n15403, n15404, n15405,
    n15406_1, n15407, n15408, n15409, n15410, n15411_1, n15412, n15413,
    n15414, n15415, n15416_1, n15417, n15418, n15419, n15420, n15421_1,
    n15422, n15423, n15424, n15425, n15426_1, n15427, n15428, n15429,
    n15430, n15431_1, n15432, n15433, n15434, n15435, n15436_1, n15437,
    n15438, n15439, n15440, n15441_1, n15442, n15443, n15444, n15445,
    n15446_1, n15447, n15448, n15449, n15450, n15451_1, n15453, n15454,
    n15455, n15456_1, n15457, n15458, n15459, n15460, n15461_1, n15462,
    n15463, n15464, n15465, n15466_1, n15467, n15468, n15469, n15470,
    n15471_1, n15472, n15473, n15474, n15475, n15476_1, n15477, n15478,
    n15479, n15480, n15481_1, n15482, n15483, n15484, n15485, n15486_1,
    n15487, n15488, n15489, n15490, n15491_1, n15492, n15493, n15494,
    n15495, n15496_1, n15497, n15498, n15499, n15500, n15501_1, n15502,
    n15503, n15504, n15505, n15506_1, n15507, n15508, n15509, n15510,
    n15511_1, n15512, n15513, n15515, n15516_1, n15517, n15518, n15519,
    n15520, n15521_1, n15522, n15523, n15524, n15525, n15526_1, n15527,
    n15528, n15529, n15530, n15531_1, n15532, n15533, n15534, n15535,
    n15536_1, n15537, n15538, n15539, n15540, n15541_1, n15542, n15543,
    n15544, n15545, n15546_1, n15547, n15548, n15549, n15550, n15551_1,
    n15552, n15553, n15554, n15555, n15556_1, n15557, n15558, n15559,
    n15560, n15561_1, n15562, n15563, n15564, n15565, n15566_1, n15567,
    n15568, n15569, n15570, n15571_1, n15572, n15574, n15575, n15576_1,
    n15577, n15578, n15579, n15580, n15581_1, n15582, n15583, n15584,
    n15585, n15586_1, n15587, n15589, n15590, n15591_1, n15592, n15593,
    n15594, n15595, n15596_1, n15597, n15599, n15600, n15601_1, n15602,
    n15604, n15605, n15607, n15608, n15610, n15611_1, n15613, n15614,
    n15616_1, n15617, n15619, n15620, n15622, n15623, n15625, n15626_1,
    n15628, n15629, n15631_1, n15632, n15634, n15635, n15637, n15638,
    n15640, n15641_1, n15643, n15644, n15646_1, n15647, n15649, n15650,
    n15652, n15653, n15655, n15656_1, n15658, n15659, n15661_1, n15662,
    n15664, n15665, n15667, n15668, n15670, n15671_1, n15673, n15674,
    n15676_1, n15677, n15679, n15680, n15682, n15683, n15685, n15686_1,
    n15688, n15689, n15691_1, n15692, n15694, n15695, n15697, n15698,
    n15699, n15700, n15701_1, n15702, n15703, n15704, n15705, n15706_1,
    n15707, n15708, n15709, n15710, n15711_1, n15712, n15713, n15714,
    n15715, n15716_1, n15717, n15718, n15719, n15720, n15721_1, n15722,
    n15723, n15724, n15726_1, n15727, n15728, n15729, n15730, n15731_1,
    n15732, n15733, n15734, n15735, n15736_1, n15737, n15739, n15740,
    n15741_1, n15742, n15743, n15744, n15745, n15746_1, n15747, n15748,
    n15749, n15750, n15752, n15753, n15754, n15755, n15756_1, n15757,
    n15758, n15759, n15760, n15761_1, n15762, n15763, n15765, n15766_1,
    n15767, n15768, n15769, n15770, n15771_1, n15772, n15773, n15774,
    n15775, n15776_1, n15778, n15779, n15780, n15781_1, n15782, n15783,
    n15784, n15785, n15786_1, n15787, n15788, n15789, n15791_1, n15792,
    n15793, n15794, n15795, n15796_1, n15797, n15798, n15799, n15800,
    n15801_1, n15802, n15804, n15805, n15806_1, n15807, n15808, n15809,
    n15810, n15811_1, n15812, n15813, n15814, n15815, n15817, n15818,
    n15819, n15820, n15821_1, n15822, n15823, n15824, n15825, n15826_1,
    n15827, n15828, n15830, n15831_1, n15832, n15833, n15834, n15835,
    n15836_1, n15837, n15838, n15839, n15840, n15841_1, n15843, n15844,
    n15845, n15846_1, n15847, n15848, n15849, n15850, n15851_1, n15852,
    n15853, n15854, n15856_1, n15857, n15858, n15859, n15860, n15861_1,
    n15862, n15863, n15864, n15865, n15866_1, n15867, n15869, n15870,
    n15871_1, n15872, n15873, n15874, n15875, n15876_1, n15877, n15878,
    n15879, n15880, n15882, n15883, n15884, n15885, n15886_1, n15887,
    n15888, n15889, n15890, n15891_1, n15892, n15893, n15895, n15896_1,
    n15897, n15898, n15899, n15900, n15901_1, n15902, n15903, n15904,
    n15905, n15906_1, n15908, n15909, n15910, n15911_1, n15912, n15913,
    n15914, n15915, n15916_1, n15917, n15918, n15919, n15921_1, n15922,
    n15923, n15924, n15925, n15926_1, n15927, n15928, n15929, n15930,
    n15931_1, n15932, n15934, n15935, n15936_1, n15937, n15938, n15939,
    n15940, n15941_1, n15942, n15943, n15944, n15945, n15947, n15948,
    n15949, n15950, n15951_1, n15952, n15953, n15954, n15955, n15956_1,
    n15957, n15958, n15960, n15961_1, n15962, n15963, n15964, n15965,
    n15966_1, n15967, n15968, n15969, n15970, n15971_1, n15973, n15974,
    n15975, n15976_1, n15977, n15978, n15979, n15980, n15981_1, n15982,
    n15983, n15984, n15986_1, n15987, n15988, n15989, n15990, n15991_1,
    n15992, n15993, n15994, n15995, n15996_1, n15998, n15999, n16000,
    n16001_1, n16002, n16003, n16004, n16005, n16006_1, n16007, n16008,
    n16010, n16011_1, n16012, n16013, n16014, n16015, n16016_1, n16017,
    n16018, n16019, n16020, n16022, n16023, n16024, n16025, n16026_1,
    n16027, n16028, n16029, n16030, n16031_1, n16032, n16034, n16035,
    n16036_1, n16037, n16038, n16039, n16040, n16041_1, n16042, n16043,
    n16044, n16046_1, n16047, n16048, n16049, n16050, n16051_1, n16052,
    n16053, n16054, n16055, n16056_1, n16058, n16059, n16060, n16061_1,
    n16062, n16063, n16064, n16065, n16066_1, n16067, n16068, n16070,
    n16071_1, n16072, n16073, n16074, n16075, n16076_1, n16077, n16078,
    n16079, n16080, n16082, n16083, n16084, n16085, n16086_1, n16087,
    n16088, n16089, n16090, n16092, n16093, n16094, n16095, n16096_1,
    n16098, n16099, n16100, n16101_1, n16103, n16104, n16105, n16106_1,
    n16107, n16109, n16110, n16111_1, n16112, n16113, n16114, n16115,
    n16116_1, n16117, n16118, n16119, n16120, n16121_1, n16122, n16123,
    n16124, n16125, n16126_1, n16127, n16128, n16129, n16130, n16131_1,
    n16132, n16133, n16134, n16135, n16136_1, n16137, n16138, n16139,
    n16140, n16141_1, n16142, n16143, n16144, n16145, n16146_1, n16147,
    n16148, n16149, n16150, n16151_1, n16152, n16153, n16154, n16155,
    n16156_1, n16157, n16158, n16159, n16160, n16161_1, n16162, n16163,
    n16164, n16165, n16166_1, n16167, n16168, n16169, n16170, n16171_1,
    n16172, n16173, n16174, n16175, n16176_1, n16177, n16178, n16179,
    n16180, n16181_1, n16182, n16183, n16184, n16185, n16186_1, n16187,
    n16188, n16189, n16190, n16191_1, n16192, n16193, n16194, n16195,
    n16196_1, n16197, n16198, n16199, n16200, n16201_1, n16202, n16203,
    n16204, n16205, n16206_1, n16207, n16208, n16209, n16210, n16211_1,
    n16212, n16213, n16214, n16215, n16216_1, n16217, n16218, n16219,
    n16220, n16221_1, n16222, n16223, n16224, n16225, n16226_1, n16227,
    n16228, n16229, n16230, n16231_1, n16232, n16233, n16234, n16235,
    n16236_1, n16237, n16238, n16239, n16240, n16241_1, n16242, n16243,
    n16244, n16245, n16246_1, n16247, n16248, n16249, n16250, n16251_1,
    n16252, n16253, n16254, n16255, n16256_1, n16257, n16258, n16259,
    n16260, n16261_1, n16262, n16263, n16264, n16265, n16266_1, n16267,
    n16268, n16269, n16270, n16271_1, n16272, n16273, n16274, n16275,
    n16276_1, n16277, n16278, n16279, n16280, n16281_1, n16282, n16283,
    n16284, n16285, n16286_1, n16287, n16288, n16289, n16290, n16291_1,
    n16292, n16293, n16294, n16295, n16296_1, n16297, n16298, n16299,
    n16300, n16301_1, n16302, n16303, n16304, n16305, n16306_1, n16307,
    n16308, n16309, n16310, n16311_1, n16312, n16313, n16314, n16315,
    n16316_1, n16317, n16318, n16319, n16320, n16321_1, n16322, n16323,
    n16324, n16325, n16326_1, n16327, n16329, n16330, n16331_1, n16332,
    n16333, n16334, n16335, n16336_1, n16337, n16338, n16339, n16340,
    n16341_1, n16342, n16343, n16344, n16345, n16346_1, n16347, n16348,
    n16349, n16350, n16351_1, n16352, n16353, n16354, n16355, n16357,
    n16358, n16359, n16360, n16361_1, n16362, n16363, n16364, n16365,
    n16366_1, n16367, n16368, n16369, n16370, n16371_1, n16372, n16373,
    n16374, n16375, n16376_1, n16377, n16378, n16379, n16380, n16381_1,
    n16382, n16383, n16384, n16385, n16386_1, n16387, n16388, n16389,
    n16390, n16391_1, n16392, n16393, n16395, n16396_1, n16397, n16398,
    n16399, n16400, n16401_1, n16402, n16403, n16404, n16405, n16406_1,
    n16407, n16408, n16409, n16410, n16411_1, n16412, n16413, n16414,
    n16415, n16416_1, n16417, n16418, n16419, n16420, n16421_1, n16422,
    n16423, n16425, n16426_1, n16427, n16428, n16429, n16430, n16431_1,
    n16432, n16433, n16434, n16435, n16436_1, n16437, n16438, n16439,
    n16440, n16441_1, n16442, n16443, n16444, n16445, n16446_1, n16447,
    n16448, n16449, n16450, n16451_1, n16453, n16454, n16455, n16456_1,
    n16457, n16458, n16459, n16460, n16461_1, n16462, n16463, n16464,
    n16465, n16466_1, n16467, n16468, n16469, n16470, n16471_1, n16472,
    n16473, n16474, n16475, n16476_1, n16477, n16478, n16479, n16481_1,
    n16482, n16483, n16484, n16485, n16486_1, n16487, n16488, n16489,
    n16490, n16491_1, n16492, n16493, n16494, n16495, n16496_1, n16497,
    n16498, n16499, n16500, n16501_1, n16502, n16503, n16504, n16505,
    n16506_1, n16507, n16508, n16509, n16510, n16511_1, n16512, n16513,
    n16514, n16515, n16516_1, n16517, n16518, n16519, n16521_1, n16522,
    n16523, n16524, n16525, n16526_1, n16527, n16528, n16529, n16530,
    n16531_1, n16532, n16533, n16534, n16535, n16536_1, n16537, n16538,
    n16539, n16540, n16541_1, n16542, n16543, n16544, n16545, n16546_1,
    n16547, n16548, n16549, n16551_1, n16552, n16553, n16554, n16555,
    n16556_1, n16557, n16558, n16559, n16560, n16561_1, n16562, n16563,
    n16564, n16565, n16566_1, n16567, n16568, n16569, n16570, n16571_1,
    n16572, n16573, n16574, n16575, n16576_1, n16577, n16578, n16579,
    n16581_1, n16582, n16583, n16584, n16585, n16586_1, n16587, n16588,
    n16589, n16590, n16591_1, n16592, n16593, n16594, n16595, n16596_1,
    n16597, n16598, n16599, n16600, n16601_1, n16602, n16603, n16604,
    n16605, n16606_1, n16607, n16608, n16609, n16610, n16611_1, n16612,
    n16613, n16614, n16615, n16616_1, n16617, n16618, n16619, n16621_1,
    n16622, n16623, n16624, n16625, n16626_1, n16627, n16628, n16629,
    n16630, n16631_1, n16632, n16633, n16634, n16635, n16636_1, n16637,
    n16638, n16639, n16640, n16641_1, n16642, n16643, n16644, n16645,
    n16646_1, n16647, n16648, n16649, n16651_1, n16652, n16653, n16654,
    n16655, n16656_1, n16657, n16658, n16659, n16660, n16661_1, n16662,
    n16663, n16664, n16665, n16666_1, n16667, n16668, n16669, n16670,
    n16671_1, n16672, n16673, n16674, n16675, n16676_1, n16677, n16678,
    n16679, n16681_1, n16682, n16683, n16684, n16685, n16686_1, n16687,
    n16688, n16689, n16690, n16691_1, n16692, n16693, n16694, n16695,
    n16696_1, n16697, n16698, n16699, n16700, n16701_1, n16702, n16703,
    n16704, n16705, n16706_1, n16707, n16708, n16709, n16710, n16711_1,
    n16712, n16713, n16714, n16715, n16716_1, n16717, n16719, n16720,
    n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
    n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
    n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
    n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
    n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
    n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
    n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
    n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
    n16794, n16795, n16796, n16797, n16799, n16800, n16801, n16802, n16803,
    n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
    n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
    n16822, n16823, n16824, n16825, n16827, n16828, n16829, n16830, n16831,
    n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
    n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
    n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
    n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
    n16868, n16869, n16870, n16871, n16873, n16874, n16875, n16876, n16877,
    n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
    n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
    n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
    n16905, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
    n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
    n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
    n16933, n16934, n16935, n16936, n16937, n16939, n16940, n16941, n16942,
    n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
    n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
    n16961, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
    n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
    n16980, n16981, n16982, n16983, n16985, n16986, n16988, n16989, n16991,
    n16992, n16994, n16995, n16997, n16998, n17000, n17001, n17003, n17004,
    n17006, n17007, n17009, n17010, n17012, n17013, n17015, n17016, n17018,
    n17019, n17021, n17022, n17024, n17025, n17027, n17028, n17030, n17031,
    n17033, n17034, n17036, n17037, n17039, n17040, n17042, n17043, n17045,
    n17046, n17048, n17049, n17051, n17052, n17054, n17055, n17057, n17058,
    n17060, n17061, n17063, n17064, n17066, n17067, n17069, n17070, n17072,
    n17073, n17075, n17076, n17078, n17079, n17081, n17082, n17083, n17084,
    n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
    n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
    n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
    n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
    n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
    n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
    n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
    n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
    n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
    n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
    n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
    n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
    n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
    n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
    n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
    n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
    n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
    n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
    n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
    n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
    n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
    n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
    n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
    n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
    n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
    n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
    n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
    n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
    n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
    n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
    n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
    n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
    n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
    n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
    n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
    n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
    n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
    n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
    n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
    n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444,
    n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
    n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
    n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
    n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
    n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
    n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
    n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
    n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
    n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
    n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
    n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
    n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
    n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
    n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
    n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
    n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
    n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
    n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
    n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
    n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
    n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
    n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
    n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
    n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
    n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
    n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
    n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
    n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
    n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
    n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
    n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
    n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
    n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
    n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
    n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
    n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
    n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
    n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
    n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
    n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
    n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
    n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
    n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
    n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
    n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
    n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
    n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
    n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
    n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
    n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
    n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
    n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
    n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
    n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
    n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
    n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
    n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
    n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
    n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
    n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
    n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
    n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
    n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
    n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
    n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
    n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
    n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
    n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
    n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
    n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
    n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
    n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
    n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
    n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
    n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
    n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
    n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
    n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
    n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
    n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
    n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
    n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
    n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
    n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
    n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
    n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
    n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
    n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
    n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
    n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
    n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
    n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
    n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
    n18283, n18284, n18285, n18286, n18288, n18289, n18290, n18291, n18292,
    n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
    n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
    n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
    n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
    n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
    n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
    n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
    n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
    n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
    n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
    n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
    n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
    n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
    n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
    n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
    n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
    n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
    n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18455,
    n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
    n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
    n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
    n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
    n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
    n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
    n18512, n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
    n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
    n18531, n18532, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
    n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
    n18550, n18551, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
    n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
    n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18578,
    n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
    n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
    n18597, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
    n18607, n18608, n18609, n18611, n18612, n18613, n18614, n18615, n18616,
    n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
    n18626, n18627, n18628, n18630, n18631, n18632, n18633, n18634, n18635,
    n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
    n18645, n18646, n18647, n18649, n18650, n18651, n18652, n18653, n18654,
    n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
    n18664, n18665, n18666, n18667, n18669, n18670, n18671, n18672, n18673,
    n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
    n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
    n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
    n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
    n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
    n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
    n18730, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
    n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
    n18749, n18750, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
    n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
    n18768, n18769, n18770, n18772, n18773, n18774, n18775, n18776, n18777,
    n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
    n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18795, n18796,
    n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
    n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18814, n18815,
    n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
    n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18833, n18834,
    n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
    n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
    n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
    n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
    n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
    n18880, n18881, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
    n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
    n18899, n18900, n18901, n18903, n18904, n18905, n18906, n18907, n18908,
    n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
    n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18927,
    n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
    n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18946,
    n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
    n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18965,
    n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
    n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18984,
    n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
    n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
    n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
    n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
    n19022, n19023, n19024, n19025, n19026, n19028, n19029, n19030, n19031,
    n19032, n19033, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
    n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19052,
    n19053, n19054, n19055, n19056, n19057, n19058, n19060, n19061, n19062,
    n19063, n19064, n19065, n19066, n19067, n19069, n19070, n19071, n19072,
    n19073, n19074, n19075, n19077, n19078, n19079, n19080, n19081, n19082,
    n19083, n19084, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
    n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
    n19103, n19104, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
    n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19123,
    n19124, n19125, n19126, n19127, n19128, n19129, n19131, n19132, n19133,
    n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19142, n19143,
    n19144, n19145, n19146, n19147, n19148, n19150, n19151, n19152, n19153,
    n19154, n19155, n19156, n19157, n19159, n19160, n19161, n19162, n19163,
    n19164, n19165, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
    n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
    n19183, n19184, n19185, n19186, n19187, n19189, n19190, n19191, n19192,
    n19193, n19194, n19195, n19197, n19198, n19199, n19200, n19201, n19202,
    n19203, n19204, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
    n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
    n19222, n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
    n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
    n19241, n19242, n19243, n19244, n19246, n19247, n19248, n19249, n19250,
    n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
    n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
    n19269, n19270, n19271, n19272, n19273, n19275, n19276, n19277, n19278,
    n19279, n19280, n19281, n19283, n19284, n19285, n19286, n19287, n19288,
    n19289, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
    n19299, n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
    n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19317, n19318,
    n19319, n19320, n19321, n19322, n19323, n19325, n19326, n19327, n19328,
    n19329, n19330, n19331, n19332, n19333, n19335, n19336, n19337, n19338,
    n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
    n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
    n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
    n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
    n19376, n19377, n19378, n19379, n19381, n19382, n19383, n19384, n19385,
    n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19395,
    n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19405,
    n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
    n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
    n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19432, n19433,
    n19434, n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
    n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
    n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
    n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
    n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
    n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
    n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
    n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
    n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
    n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
    n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
    n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
    n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
    n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
    n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
    n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
    n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
    n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
    n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
    n19636, n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
    n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
    n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
    n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
    n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
    n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
    n19691, n19692, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
    n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
    n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
    n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
    n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
    n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
    n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19754, n19755,
    n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
    n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
    n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
    n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
    n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
    n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
    n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19819,
    n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
    n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
    n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
    n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
    n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
    n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
    n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
    n19883, n19884, n19885, n19886, n19887, n19888, n19890, n19891, n19892,
    n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
    n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
    n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
    n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
    n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
    n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
    n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19955, n19956,
    n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
    n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
    n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
    n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
    n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
    n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
    n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
    n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20029,
    n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
    n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
    n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
    n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
    n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
    n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
    n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
    n20093, n20094, n20095, n20096, n20097, n20099, n20100, n20101, n20102,
    n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
    n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
    n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
    n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
    n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
    n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
    n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
    n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
    n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
    n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
    n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
    n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
    n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
    n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
    n20230, n20231, n20232, n20233, n20234, n20235, n20237, n20238, n20239,
    n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
    n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
    n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
    n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
    n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
    n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
    n20294, n20295, n20296, n20297, n20298, n20299, n20301, n20302, n20303,
    n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
    n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
    n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
    n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
    n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
    n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
    n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
    n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
    n20376, n20377, n20378, n20380, n20381, n20382, n20383, n20384, n20385,
    n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
    n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
    n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
    n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
    n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
    n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
    n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
    n20449, n20450, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
    n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
    n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
    n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
    n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
    n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
    n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
    n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
    n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
    n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
    n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
    n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
    n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
    n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
    n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
    n20586, n20587, n20588, n20589, n20590, n20592, n20593, n20594, n20595,
    n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
    n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
    n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
    n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
    n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
    n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
    n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
    n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
    n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
    n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
    n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
    n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
    n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
    n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
    n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20732,
    n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
    n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
    n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
    n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
    n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
    n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
    n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
    n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
    n20805, n20806, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
    n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
    n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
    n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
    n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
    n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
    n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
    n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
    n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
    n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
    n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
    n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
    n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
    n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
    n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
    n20942, n20943, n20944, n20945, n20947, n20948, n20949, n20950, n20951,
    n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960,
    n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
    n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
    n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
    n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
    n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
    n21006, n21007, n21008, n21009, n21011, n21012, n21013, n21014, n21015,
    n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024,
    n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
    n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
    n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
    n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
    n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
    n21070, n21071, n21072, n21073, n21074, n21075, n21077, n21078, n21079,
    n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088,
    n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
    n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
    n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
    n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
    n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
    n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
    n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152,
    n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
    n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
    n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
    n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
    n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
    n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206,
    n21207, n21208, n21210, n21211, n21212, n21213, n21214, n21215, n21216,
    n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
    n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234,
    n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
    n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252,
    n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261,
    n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270,
    n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21279, n21280,
    n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
    n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
    n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
    n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
    n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
    n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334,
    n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21343, n21344,
    n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
    n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362,
    n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
    n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380,
    n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389,
    n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398,
    n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407,
    n21408, n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
    n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426,
    n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435,
    n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444,
    n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453,
    n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462,
    n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471,
    n21472, n21473, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
    n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490,
    n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
    n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508,
    n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517,
    n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526,
    n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535,
    n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544,
    n21545, n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554,
    n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
    n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572,
    n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581,
    n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590,
    n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599,
    n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608,
    n21609, n21610, n21611, n21612, n21614, n21615, n21616, n21617, n21618,
    n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627,
    n21628, n21629, n21630, n21632, n21633, n21634, n21635, n21636, n21637,
    n21638, n21639, n21640, n21641, n21643, n21644, n21645, n21646, n21648,
    n21649, n21651, n21652, n21654, n21655, n21657, n21658, n21660, n21661,
    n21663, n21664, n21666, n21667, n21669, n21670, n21672, n21673, n21675,
    n21676, n21678, n21679, n21681, n21682, n21684, n21685, n21687, n21688,
    n21690, n21691, n21693, n21694, n21696, n21697, n21699, n21700, n21702,
    n21703, n21705, n21706, n21708, n21709, n21711, n21712, n21714, n21715,
    n21717, n21718, n21720, n21721, n21723, n21724, n21726, n21727, n21729,
    n21730, n21732, n21733, n21735, n21736, n21738, n21739, n21741, n21742,
    n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751,
    n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760,
    n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21770,
    n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
    n21780, n21781, n21783, n21784, n21785, n21786, n21787, n21788, n21789,
    n21790, n21791, n21792, n21793, n21794, n21796, n21797, n21798, n21799,
    n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21809,
    n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818,
    n21819, n21820, n21822, n21823, n21824, n21825, n21826, n21827, n21828,
    n21829, n21830, n21831, n21832, n21833, n21835, n21836, n21837, n21838,
    n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21848,
    n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
    n21858, n21859, n21861, n21862, n21863, n21864, n21865, n21866, n21867,
    n21868, n21869, n21870, n21871, n21872, n21874, n21875, n21876, n21877,
    n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21887,
    n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896,
    n21897, n21898, n21900, n21901, n21902, n21903, n21904, n21905, n21906,
    n21907, n21908, n21909, n21910, n21911, n21913, n21914, n21915, n21916,
    n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21926,
    n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
    n21936, n21937, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
    n21946, n21947, n21948, n21949, n21950, n21952, n21953, n21954, n21955,
    n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21965,
    n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974,
    n21975, n21976, n21978, n21979, n21980, n21981, n21982, n21983, n21984,
    n21985, n21986, n21987, n21988, n21989, n21991, n21992, n21993, n21994,
    n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22004,
    n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013,
    n22014, n22015, n22017, n22018, n22019, n22020, n22021, n22022, n22023,
    n22024, n22025, n22026, n22027, n22028, n22030, n22031, n22032, n22033,
    n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22043,
    n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052,
    n22053, n22054, n22056, n22057, n22058, n22059, n22060, n22061, n22062,
    n22063, n22064, n22065, n22066, n22067, n22069, n22070, n22071, n22072,
    n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22082,
    n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091,
    n22092, n22093, n22095, n22096, n22097, n22098, n22099, n22100, n22101,
    n22102, n22103, n22104, n22105, n22106, n22108, n22109, n22110, n22111,
    n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22121,
    n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130,
    n22131, n22132, n22134, n22135, n22136, n22137, n22138, n22139, n22140,
    n22141, n22142, n22143, n22145, n22146, n22147, n22148, n22149, n22150,
    n22152, n22153, n22154, n22155, n22156, n22158, n22159, n22160, n22161,
    n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171,
    n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180,
    n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189,
    n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198,
    n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207,
    n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216,
    n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
    n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234,
    n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243,
    n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252,
    n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261,
    n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270,
    n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279,
    n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288,
    n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
    n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306,
    n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315,
    n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324,
    n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333,
    n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342,
    n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351,
    n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360,
    n22361, n22362, n22364, n22365, n22366, n22367, n22368, n22369, n22370,
    n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379,
    n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388,
    n22389, n22390, n22392, n22393, n22394, n22395, n22396, n22397, n22398,
    n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407,
    n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416,
    n22417, n22418, n22420, n22421, n22422, n22423, n22424, n22425, n22426,
    n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435,
    n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444,
    n22445, n22446, n22448, n22449, n22450, n22451, n22452, n22453, n22454,
    n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463,
    n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472,
    n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482,
    n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491,
    n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22500, n22501,
    n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510,
    n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519,
    n22520, n22521, n22522, n22523, n22524, n22526, n22527, n22528, n22529,
    n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538,
    n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547,
    n22548, n22549, n22550, n22551, n22552, n22554, n22555, n22556, n22557,
    n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566,
    n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575,
    n22576, n22577, n22578, n22579, n22580, n22582, n22583, n22584, n22585,
    n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594,
    n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603,
    n22604, n22605, n22606, n22608, n22609, n22610, n22611, n22612, n22613,
    n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622,
    n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631,
    n22632, n22633, n22634, n22636, n22637, n22638, n22639, n22640, n22641,
    n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650,
    n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659,
    n22660, n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669,
    n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678,
    n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687,
    n22688, n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
    n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706,
    n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715,
    n22716, n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725,
    n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734,
    n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22744,
    n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
    n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762,
    n22763, n22764, n22765, n22766, n22767, n22768, n22770, n22771, n22772,
    n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781,
    n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790,
    n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799,
    n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808,
    n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22817, n22818,
    n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827,
    n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836,
    n22837, n22838, n22839, n22840, n22841, n22842, n22844, n22845, n22846,
    n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855,
    n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864,
    n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22873, n22874,
    n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883,
    n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892,
    n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901,
    n22902, n22903, n22904, n22905, n22907, n22908, n22909, n22910, n22911,
    n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920,
    n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22929, n22930,
    n22932, n22933, n22935, n22936, n22938, n22939, n22941, n22942, n22944,
    n22945, n22947, n22948, n22950, n22951, n22953, n22954, n22956, n22957,
    n22959, n22960, n22962, n22963, n22965, n22966, n22968, n22969, n22971,
    n22972, n22974, n22975, n22977, n22978, n22980, n22981, n22983, n22984,
    n22986, n22987, n22989, n22990, n22992, n22993, n22995, n22996, n22998,
    n22999, n23001, n23002, n23004, n23005, n23007, n23008, n23010, n23011,
    n23013, n23014, n23016, n23017, n23019, n23020, n23022, n23023, n23025,
    n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034,
    n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043,
    n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052,
    n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061,
    n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070,
    n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079,
    n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088,
    n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
    n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106,
    n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115,
    n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124,
    n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133,
    n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142,
    n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151,
    n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160,
    n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
    n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178,
    n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187,
    n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196,
    n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205,
    n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214,
    n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223,
    n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232,
    n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
    n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250,
    n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259,
    n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268,
    n23269, n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277,
    n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286,
    n23287, n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295,
    n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304,
    n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
    n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322,
    n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331,
    n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340,
    n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349,
    n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358,
    n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367,
    n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376,
    n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
    n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394,
    n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403,
    n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412,
    n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421,
    n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430,
    n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439,
    n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448,
    n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
    n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466,
    n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475,
    n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484,
    n23485, n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493,
    n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502,
    n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511,
    n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520,
    n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
    n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538,
    n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547,
    n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556,
    n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565,
    n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574,
    n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583,
    n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592,
    n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
    n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610,
    n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619,
    n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628,
    n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637,
    n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646,
    n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655,
    n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664,
    n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
    n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682,
    n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691,
    n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700,
    n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709,
    n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718,
    n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727,
    n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736,
    n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
    n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754,
    n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763,
    n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772,
    n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781,
    n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790,
    n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799,
    n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808,
    n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
    n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826,
    n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835,
    n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844,
    n23845, n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853,
    n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862,
    n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871,
    n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880,
    n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
    n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898,
    n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907,
    n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916,
    n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925,
    n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934,
    n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943,
    n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952,
    n23953, n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
    n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970,
    n23971, n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979,
    n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988,
    n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997,
    n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006,
    n24007, n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015,
    n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024,
    n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
    n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042,
    n24043, n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051,
    n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24061,
    n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070,
    n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079,
    n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088,
    n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
    n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106,
    n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115,
    n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123, n24124,
    n24125, n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133,
    n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142,
    n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151,
    n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160,
    n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
    n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178,
    n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187,
    n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196,
    n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205,
    n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214,
    n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223,
    n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232,
    n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
    n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250,
    n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259,
    n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268,
    n24269, n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277,
    n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286,
    n24287, n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295,
    n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304,
    n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24313, n24314,
    n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323,
    n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331, n24332,
    n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341,
    n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349, n24350,
    n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359,
    n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368,
    n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
    n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386,
    n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395,
    n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403, n24404,
    n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412, n24413,
    n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421, n24422,
    n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24431,
    n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439, n24440,
    n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
    n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458,
    n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467,
    n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475, n24476,
    n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484, n24485,
    n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493, n24494,
    n24495, n24496, n24498, n24499, n24500, n24501, n24502, n24503, n24504,
    n24505, n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
    n24514, n24515, n24516, n24517, n24518, n24520, n24521, n24522, n24523,
    n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532,
    n24533, n24534, n24535, n24536, n24537, n24539, n24540, n24541, n24542,
    n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551,
    n24552, n24553, n24554, n24555, n24556, n24557, n24559, n24560, n24561,
    n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570,
    n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24579, n24580,
    n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589,
    n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597, n24599,
    n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608,
    n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
    n24618, n24619, n24620, n24621, n24622, n24624, n24625, n24626, n24627,
    n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636,
    n24637, n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645,
    n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655,
    n24656, n24657, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
    n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674,
    n24675, n24676, n24678, n24679, n24680, n24681, n24682, n24683, n24684,
    n24685, n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693,
    n24694, n24695, n24697, n24698, n24699, n24700, n24701, n24702, n24703,
    n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712,
    n24713, n24714, n24715, n24716, n24718, n24719, n24720, n24721, n24722,
    n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731,
    n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740,
    n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750,
    n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759,
    n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
    n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778,
    n24779, n24781, n24782, n24783, n24784, n24785, n24786, n24787, n24788,
    n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796, n24797,
    n24798, n24799, n24800, n24801, n24803, n24804, n24805, n24806, n24807,
    n24808, n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816,
    n24817, n24818, n24819, n24820, n24821, n24823, n24824, n24825, n24826,
    n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835,
    n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844,
    n24845, n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854,
    n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863,
    n24864, n24865, n24866, n24868, n24869, n24870, n24871, n24872, n24873,
    n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882,
    n24883, n24884, n24885, n24887, n24888, n24889, n24890, n24891, n24892,
    n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901,
    n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910,
    n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919,
    n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928,
    n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
    n24938, n24939, n24940, n24941, n24942, n24943, n24945, n24946, n24947,
    n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956,
    n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24965, n24966,
    n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975,
    n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984,
    n24985, n24986, n24987, n24989, n24990, n24991, n24992, n24993, n24994,
    n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003,
    n25004, n25005, n25006, n25008, n25009, n25010, n25011, n25012, n25013,
    n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022,
    n25023, n25024, n25025, n25026, n25028, n25029, n25030, n25031, n25032,
    n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
    n25042, n25043, n25044, n25045, n25047, n25048, n25049, n25050, n25051,
    n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060,
    n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25070,
    n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079,
    n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088,
    n25089, n25090, n25091, n25092, n25094, n25095, n25096, n25098, n25099,
    n25101, n25102, n25104, n25105, n25107, n25108, n25109, n25110, n25111,
    n25112, n25114, n25115, n25116, n25117, n25119, n25120, n25121, n25122,
    n25124, n25125, n25126, n25127, n25129, n25130, n25131, n25132, n25134,
    n25135, n25136, n25137, n25139, n25140, n25141, n25142, n25144, n25145,
    n25146, n25147, n25149, n25150, n25151, n25152, n25154, n25155, n25156,
    n25157, n25159, n25160, n25161, n25162, n25164, n25165, n25166, n25167,
    n25169, n25170, n25171, n25172, n25174, n25175, n25176, n25177, n25179,
    n25180, n25181, n25182, n25184, n25185, n25186, n25187, n25189, n25190,
    n25191, n25192, n25194, n25195, n25196, n25197, n25199, n25200, n25201,
    n25202, n25204, n25205, n25206, n25207, n25209, n25210, n25211, n25212,
    n25214, n25215, n25216, n25217, n25219, n25220, n25221, n25222, n25224,
    n25225, n25226, n25227, n25229, n25230, n25231, n25232, n25234, n25235,
    n25236, n25237, n25239, n25240, n25241, n25242, n25244, n25245, n25246,
    n25247, n25249, n25250, n25251, n25252, n25254, n25255, n25256, n25257,
    n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267,
    n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276,
    n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285,
    n25286, n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295,
    n25296, n25297, n25298, n25299, n25300, n25302, n25303, n25304, n25305,
    n25306, n25307, n25308, n25309, n25310, n25312, n25313, n25314, n25315,
    n25316, n25317, n25319, n25320, n25352, n25353, n25354, n25355, n25356,
    n25357, n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365,
    n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374,
    n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383,
    n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392,
    n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
    n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410,
    n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419,
    n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428,
    n25429, n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437,
    n25438, n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446,
    n25447, n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455,
    n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464,
    n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
    n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482,
    n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491,
    n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500,
    n25501, n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509,
    n25510, n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518,
    n25519, n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527,
    n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536,
    n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
    n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554,
    n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563,
    n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572,
    n25573, n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581,
    n25582, n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590,
    n25591, n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599,
    n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608,
    n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
    n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626,
    n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635,
    n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644,
    n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653,
    n25654, n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662,
    n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671,
    n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680,
    n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
    n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698,
    n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707,
    n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716,
    n25717, n25718, n25719, n25720, n25721, n25722, n25723, n25724, n25725,
    n25726, n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734,
    n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743,
    n25744, n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752,
    n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
    n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770,
    n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779,
    n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787, n25788,
    n25789, n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797,
    n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806,
    n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815,
    n25816, n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824,
    n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
    n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842,
    n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851,
    n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860,
    n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868, n25869,
    n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878,
    n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887,
    n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896,
    n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
    n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914,
    n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923,
    n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931, n25932,
    n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940, n25941,
    n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950,
    n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959,
    n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968,
    n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
    n25978, n25979, n25980, n25981, n25982, n25983, n25985, n25986, n25987,
    n25988, n25989, n25990, n25991, n25992, n25994, n25995, n25996, n25997,
    n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006,
    n26007, n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016,
    n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
    n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034,
    n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043,
    n26044, n26045, n26046, n26047, n26048, n26050, n26051, n26052, n26053,
    n26054, n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062,
    n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071,
    n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080,
    n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
    n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098,
    n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107,
    n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116,
    n26117, n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125,
    n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135,
    n26136, n26137, n26138, n26140, n26141, n26142, n26143, n26144, n26145,
    n26146, n26147, n26148, n26149, n26150, n26151, n26153, n26154, n26155,
    n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163, n26164,
    n26166, n26167, n26168, n26169, n26170, n26171, n26172, n26173, n26174,
    n26175, n26176, n26177, n26179, n26180, n26181, n26182, n26183, n26184,
    n26185, n26186, n26187, n26188, n26189, n26190, n26192, n26193, n26194,
    n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203,
    n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213,
    n26214, n26215, n26216, n26218, n26219, n26220, n26221, n26222, n26223,
    n26224, n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232,
    n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
    n26242, n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251,
    n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26262,
    n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26271, n26272,
    n26273, n26274, n26275, n26276, n26277, n26278, n26280, n26281, n26282,
    n26283, n26284, n26285, n26286, n26287, n26289, n26290, n26291, n26292,
    n26293, n26294, n26295, n26296, n26298, n26299, n26300, n26301, n26302,
    n26303, n26304, n26305, n26307, n26308, n26309, n26310, n26311, n26312,
    n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
    n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330,
    n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339, n26341,
    n26342, n26343, n26344, n26345, n26346, n26347, n26348, n26350, n26351,
    n26352, n26353, n26354, n26355, n26356, n26357, n26359, n26360, n26361,
    n26362, n26363, n26364, n26365, n26366, n26368, n26369, n26370, n26371,
    n26372, n26373, n26374, n26375, n26377, n26378, n26379, n26380, n26381,
    n26382, n26383, n26384, n26386, n26387, n26388, n26389, n26390, n26391,
    n26392, n26393, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
    n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410,
    n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26420,
    n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26429, n26430,
    n26431, n26432, n26433, n26434, n26435, n26436, n26438, n26439, n26440,
    n26441, n26442, n26443, n26444, n26445, n26447, n26448, n26449, n26450,
    n26451, n26452, n26453, n26454, n26456, n26457, n26458, n26459, n26460,
    n26461, n26462, n26463, n26465, n26466, n26467, n26468, n26469, n26470,
    n26471, n26472, n26474, n26475, n26476, n26477, n26478, n26479, n26480,
    n26481, n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490,
    n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499,
    n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26509,
    n26510, n26511, n26512, n26513, n26514, n26515, n26516, n26518, n26519,
    n26520, n26521, n26522, n26523, n26524, n26525, n26527, n26528, n26529,
    n26530, n26531, n26532, n26533, n26534, n26536, n26537, n26538, n26539,
    n26540, n26541, n26542, n26543, n26545, n26546, n26547, n26548, n26549,
    n26550, n26551, n26552, n26554, n26555, n26556, n26557, n26558, n26559,
    n26560, n26561, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
    n26570, n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579,
    n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588,
    n26589, n26590, n26591, n26592, n26593, n26594, n26596, n26597, n26598,
    n26599, n26600, n26601, n26602, n26603, n26605, n26606, n26607, n26608,
    n26609, n26610, n26611, n26612, n26614, n26615, n26616, n26617, n26618,
    n26619, n26620, n26621, n26623, n26624, n26625, n26626, n26627, n26628,
    n26629, n26630, n26632, n26633, n26634, n26635, n26636, n26637, n26638,
    n26639, n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648,
    n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26659,
    n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668,
    n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676, n26677,
    n26678, n26679, n26680, n26682, n26683, n26684, n26685, n26686, n26687,
    n26688, n26689, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
    n26698, n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707,
    n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716, n26718,
    n26719, n26720, n26721, n26722, n26723, n26724, n26725, n26727, n26728,
    n26729, n26730, n26731, n26732, n26733, n26734, n26736, n26737, n26738,
    n26739, n26740, n26741, n26742, n26743, n26745, n26746, n26747, n26748,
    n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756, n26757,
    n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765, n26767,
    n26768, n26769, n26770, n26771, n26772, n26773, n26774, n26776, n26777,
    n26778, n26779, n26780, n26781, n26782, n26783, n26785, n26786, n26787,
    n26788, n26789, n26790, n26791, n26792, n26794, n26795, n26796, n26797,
    n26798, n26799, n26800, n26801, n26803, n26804, n26805, n26806, n26807,
    n26808, n26809, n26810, n26812, n26813, n26814, n26815, n26816, n26817,
    n26818, n26819, n26821, n26822, n26823, n26824, n26825, n26826, n26827,
    n26828, n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837,
    n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845, n26846,
    n26847, n26848, n26849, n26851, n26852, n26853, n26854, n26855, n26856,
    n26857, n26858, n26860, n26861, n26862, n26863, n26864, n26865, n26866,
    n26867, n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876,
    n26878, n26879, n26880, n26881, n26882, n26883, n26884, n26885, n26887,
    n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26896, n26897,
    n26898, n26899, n26900, n26901, n26902, n26903, n26905, n26906, n26907,
    n26908, n26909, n26910, n26911, n26912, n26914, n26915, n26916, n26917,
    n26918, n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926,
    n26927, n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935,
    n26936, n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
    n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26956,
    n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26965, n26966,
    n26967, n26968, n26969, n26970, n26971, n26972, n26974, n26975, n26976,
    n26977, n26978, n26979, n26980, n26981, n26983, n26984, n26985, n26986,
    n26987, n26988, n26989, n26990, n26992, n26993, n26994, n26995, n26996,
    n26997, n26998, n26999, n27001, n27002, n27003, n27004, n27005, n27006,
    n27007, n27008, n27009, n27010, n27011, n27012, n27013, n27014, n27015,
    n27016, n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27025,
    n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27034, n27035,
    n27036, n27037, n27038, n27039, n27040, n27041, n27043, n27044, n27045,
    n27046, n27047, n27048, n27049, n27050, n27052, n27053, n27054, n27055,
    n27056, n27057, n27058, n27059, n27061, n27062, n27063, n27064, n27065,
    n27066, n27067, n27068, n27070, n27071, n27072, n27073, n27074, n27075,
    n27076, n27077, n27079, n27080, n27081, n27082, n27083, n27084, n27085,
    n27086, n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095,
    n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104,
    n27105, n27106, n27107, n27108, n27110, n27111, n27112, n27113, n27114,
    n27115, n27116, n27117, n27119, n27120, n27121, n27122, n27123, n27124,
    n27125, n27126, n27128, n27129, n27130, n27131, n27132, n27133, n27134,
    n27135, n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144,
    n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27155,
    n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27164, n27165,
    n27166, n27167, n27168, n27169, n27170, n27171, n27173, n27174, n27175,
    n27176, n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184,
    n27185, n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
    n27194, n27195, n27196, n27198, n27199, n27200, n27201, n27202, n27203,
    n27204, n27205, n27207, n27208, n27209, n27210, n27211, n27212, n27213,
    n27214, n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223,
    n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27234,
    n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27243, n27244,
    n27245, n27246, n27247, n27248, n27249, n27250, n27252, n27253, n27254,
    n27255, n27256, n27257, n27258, n27259, n27261, n27262, n27263, n27264,
    n27265, n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
    n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27282, n27283,
    n27284, n27285, n27286, n27287, n27288, n27289, n27291, n27292, n27293,
    n27294, n27295, n27296, n27297, n27298, n27300, n27301, n27302, n27303,
    n27304, n27305, n27306, n27307, n27309, n27310, n27311, n27312, n27313,
    n27314, n27315, n27316, n27318, n27319, n27320, n27321, n27322, n27323,
    n27324, n27325, n27327, n27328, n27329, n27330, n27331, n27332, n27333,
    n27334, n27336, n27337, n27338, n27339, n27340, n27341, n27342, n27343,
    n27345, n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
    n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361, n27362,
    n27363, n27364, n27366, n27367, n27368, n27369, n27370, n27371, n27372,
    n27373, n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382,
    n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27393,
    n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27402, n27403,
    n27404, n27405, n27406, n27407, n27408, n27409, n27411, n27412, n27413,
    n27414, n27415, n27416, n27417, n27418, n27420, n27421, n27422, n27423,
    n27424, n27425, n27426, n27427, n27429, n27430, n27431, n27432, n27433,
    n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441, n27442,
    n27443, n27444, n27445, n27446, n27447, n27449, n27450, n27451, n27452,
    n27453, n27454, n27455, n27456, n27458, n27459, n27460, n27461, n27462,
    n27463, n27464, n27465, n27467, n27468, n27469, n27470, n27471, n27472,
    n27473, n27474, n27476, n27477, n27478, n27479, n27480, n27481, n27482,
    n27483, n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492,
    n27494, n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27503,
    n27504, n27505, n27506, n27507, n27508, n27509, n27510, n27512, n27513,
    n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27523,
    n27524, n27525, n27526, n27527, n27528, n27530, n27531, n27532, n27533,
    n27534, n27535, n27536, n27537, n27539, n27540, n27541, n27542, n27543,
    n27544, n27545, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
    n27555, n27556, n27557, n27558, n27560, n27561, n27562, n27563, n27564,
    n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27574,
    n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583,
    n27584, n27585, n27586, n27588, n27589, n27590, n27591, n27592, n27593,
    n27594, n27595, n27596, n27597, n27598, n27599, n27601, n27602, n27603,
    n27604, n27605, n27607, n27608, n27609, n27610, n27611, n27612, n27613,
    n27614, n27615, n27616, n27617, n27618, n27619, n27620, n27621, n27622,
    n27623, n27624, n27625, n27626, n27627, n27628, n27629, n27630, n27631,
    n27632, n27633, n27634, n27635, n27636, n27637, n27638, n27639, n27640,
    n27641, n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
    n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657, n27658,
    n27659, n27660, n27661, n27662, n27663, n27664, n27665, n27666, n27667,
    n27668, n27669, n27670, n27671, n27672, n27673, n27674, n27675, n27676,
    n27677, n27678, n27679, n27680, n27681, n27682, n27683, n27684, n27685,
    n27686, n27687, n27688, n27689, n27690, n27691, n27692, n27693, n27694,
    n27695, n27696, n27697, n27698, n27699, n27700, n27701, n27702, n27703,
    n27704, n27705, n27706, n27707, n27708, n27709, n27710, n27711, n27712,
    n27713, n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
    n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729, n27730,
    n27731, n27732, n27733, n27734, n27735, n27736, n27737, n27738, n27739,
    n27740, n27741, n27742, n27743, n27744, n27745, n27746, n27747, n27748,
    n27749, n27750, n27751, n27752, n27753, n27754, n27755, n27756, n27757,
    n27758, n27759, n27760, n27761, n27762, n27763, n27764, n27765, n27766,
    n27767, n27768, n27769, n27770, n27771, n27772, n27773, n27774, n27775,
    n27776, n27777, n27778, n27779, n27780, n27781, n27783, n27784, n27785,
    n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794,
    n27795, n27796, n27797, n27798, n27799, n27800, n27801, n27802, n27803,
    n27804, n27805, n27806, n27807, n27808, n27809, n27810, n27811, n27812,
    n27813, n27814, n27815, n27816, n27817, n27818, n27819, n27820, n27821,
    n27822, n27823, n27824, n27825, n27826, n27827, n27828, n27829, n27830,
    n27831, n27832, n27833, n27834, n27835, n27836, n27837, n27838, n27839,
    n27840, n27841, n27842, n27843, n27844, n27845, n27846, n27847, n27848,
    n27849, n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
    n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865, n27866,
    n27867, n27868, n27869, n27870, n27871, n27872, n27873, n27874, n27875,
    n27876, n27877, n27878, n27879, n27881, n27882, n27883, n27884, n27885,
    n27886, n27887, n27888, n27889, n27890, n27891, n27892, n27893, n27894,
    n27895, n27896, n27897, n27898, n27899, n27900, n27901, n27902, n27903,
    n27904, n27905, n27906, n27907, n27908, n27909, n27910, n27911, n27912,
    n27913, n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
    n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929, n27930,
    n27931, n27932, n27933, n27934, n27935, n27936, n27937, n27938, n27939,
    n27940, n27941, n27942, n27943, n27944, n27945, n27946, n27947, n27948,
    n27949, n27950, n27951, n27952, n27953, n27954, n27955, n27956, n27957,
    n27958, n27959, n27960, n27961, n27962, n27963, n27964, n27965, n27966,
    n27967, n27968, n27969, n27970, n27971, n27972, n27973, n27974, n27975,
    n27976, n27977, n27978, n27979, n27980, n27981, n27982, n27983, n27984,
    n27985, n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
    n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001, n28002,
    n28004, n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012,
    n28013, n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28021,
    n28022, n28023, n28024, n28025, n28026, n28027, n28028, n28029, n28030,
    n28031, n28032, n28033, n28034, n28035, n28036, n28037, n28038, n28039,
    n28040, n28041, n28042, n28043, n28044, n28045, n28046, n28047, n28048,
    n28049, n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
    n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066,
    n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075,
    n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084,
    n28085, n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093,
    n28094, n28095, n28096, n28097, n28098, n28099, n28100, n28101, n28102,
    n28103, n28104, n28105, n28106, n28107, n28108, n28109, n28110, n28111,
    n28112, n28113, n28114, n28115, n28116, n28117, n28118, n28119, n28120,
    n28121, n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
    n28130, n28131, n28132, n28133, n28135, n28136, n28137, n28138, n28139,
    n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148,
    n28149, n28150, n28151, n28152, n28153, n28154, n28155, n28156, n28157,
    n28158, n28159, n28160, n28161, n28162, n28163, n28164, n28165, n28166,
    n28167, n28168, n28169, n28170, n28171, n28172, n28173, n28174, n28175,
    n28176, n28177, n28178, n28179, n28180, n28181, n28182, n28183, n28184,
    n28185, n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
    n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202,
    n28203, n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211,
    n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219, n28220,
    n28221, n28222, n28223, n28224, n28225, n28226, n28227, n28228, n28229,
    n28230, n28231, n28232, n28233, n28234, n28235, n28236, n28237, n28238,
    n28239, n28240, n28241, n28242, n28243, n28244, n28245, n28246, n28247,
    n28248, n28249, n28250, n28251, n28252, n28253, n28254, n28255, n28256,
    n28257, n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
    n28266, n28267, n28268, n28269, n28271, n28272, n28273, n28274, n28275,
    n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284,
    n28285, n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28293,
    n28294, n28295, n28296, n28297, n28298, n28299, n28300, n28301, n28302,
    n28303, n28304, n28305, n28306, n28307, n28308, n28309, n28310, n28311,
    n28312, n28313, n28314, n28315, n28316, n28317, n28318, n28319, n28320,
    n28321, n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
    n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338,
    n28339, n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347,
    n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355, n28356,
    n28357, n28358, n28359, n28360, n28361, n28362, n28363, n28364, n28365,
    n28366, n28367, n28368, n28369, n28370, n28371, n28372, n28373, n28374,
    n28375, n28376, n28377, n28378, n28379, n28380, n28381, n28382, n28383,
    n28384, n28385, n28386, n28387, n28388, n28389, n28390, n28391, n28392,
    n28393, n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
    n28402, n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411,
    n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420,
    n28421, n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429,
    n28430, n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438,
    n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446, n28447,
    n28448, n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456,
    n28457, n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
    n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474,
    n28475, n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483,
    n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492,
    n28493, n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501,
    n28502, n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510,
    n28511, n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519,
    n28520, n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528,
    n28529, n28530, n28531, n28532, n28533, n28535, n28536, n28537, n28538,
    n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547,
    n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555, n28556,
    n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564, n28565,
    n28566, n28567, n28568, n28569, n28570, n28571, n28572, n28573, n28574,
    n28575, n28576, n28577, n28578, n28579, n28580, n28581, n28582, n28583,
    n28584, n28585, n28586, n28587, n28588, n28589, n28590, n28591, n28592,
    n28593, n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
    n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610,
    n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619,
    n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627, n28628,
    n28629, n28630, n28631, n28633, n28634, n28635, n28636, n28637, n28638,
    n28639, n28640, n28641, n28642, n28643, n28644, n28645, n28646, n28647,
    n28648, n28649, n28650, n28651, n28652, n28653, n28654, n28655, n28656,
    n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
    n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673, n28674,
    n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683,
    n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691, n28692,
    n28693, n28694, n28695, n28696, n28697, n28698, n28699, n28700, n28701,
    n28702, n28703, n28704, n28705, n28706, n28707, n28708, n28709, n28710,
    n28711, n28712, n28713, n28714, n28715, n28716, n28717, n28718, n28719,
    n28720, n28721, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
    n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737, n28738,
    n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747,
    n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755, n28756,
    n28757, n28758, n28759, n28760, n28761, n28762, n28763, n28764, n28765,
    n28766, n28767, n28768, n28769, n28770, n28771, n28772, n28773, n28774,
    n28775, n28776, n28777, n28778, n28779, n28780, n28781, n28782, n28783,
    n28784, n28785, n28786, n28787, n28788, n28789, n28790, n28791, n28792,
    n28793, n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
    n28802, n28803, n28804, n28805, n28807, n28808, n28809, n28810, n28811,
    n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819, n28820,
    n28821, n28822, n28823, n28824, n28825, n28826, n28827, n28828, n28829,
    n28830, n28831, n28832, n28833, n28834, n28835, n28836, n28837, n28838,
    n28839, n28840, n28841, n28842, n28843, n28844, n28845, n28846, n28847,
    n28848, n28849, n28850, n28851, n28852, n28853, n28854, n28855, n28856,
    n28857, n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
    n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873, n28874,
    n28875, n28876, n28877, n28878, n28879, n28881, n28882, n28883, n28884,
    n28885, n28886, n28887, n28888, n28889, n28890, n28891, n28892, n28893,
    n28894, n28895, n28896, n28897, n28898, n28899, n28900, n28901, n28902,
    n28903, n28904, n28905, n28906, n28907, n28908, n28909, n28910, n28911,
    n28912, n28913, n28914, n28915, n28916, n28917, n28918, n28919, n28920,
    n28921, n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
    n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937, n28938,
    n28939, n28940, n28941, n28942, n28943, n28944, n28945, n28946, n28947,
    n28948, n28949, n28950, n28951, n28953, n28954, n28955, n28956, n28957,
    n28958, n28959, n28960, n28961, n28962, n28963, n28964, n28965, n28966,
    n28967, n28968, n28969, n28970, n28971, n28972, n28973, n28974, n28975,
    n28976, n28977, n28978, n28979, n28980, n28981, n28982, n28983, n28984,
    n28985, n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
    n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001, n29002,
    n29003, n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011,
    n29012, n29013, n29014, n29015, n29016, n29017, n29018, n29019, n29020,
    n29021, n29022, n29023, n29024, n29025, n29026, n29027, n29028, n29029,
    n29030, n29031, n29033, n29034, n29035, n29036, n29037, n29038, n29039,
    n29040, n29041, n29042, n29043, n29044, n29045, n29046, n29047, n29048,
    n29049, n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
    n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065, n29066,
    n29067, n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075,
    n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083, n29084,
    n29085, n29086, n29087, n29088, n29089, n29090, n29091, n29092, n29093,
    n29094, n29095, n29096, n29097, n29098, n29099, n29100, n29101, n29102,
    n29103, n29104, n29105, n29106, n29108, n29109, n29110, n29111, n29112,
    n29113, n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
    n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129, n29130,
    n29131, n29132, n29133, n29134, n29135, n29136, n29137, n29138, n29139,
    n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147, n29148,
    n29149, n29150, n29151, n29152, n29153, n29154, n29155, n29156, n29157,
    n29158, n29159, n29160, n29161, n29162, n29163, n29164, n29165, n29166,
    n29167, n29168, n29169, n29170, n29171, n29172, n29173, n29174, n29175,
    n29176, n29177, n29178, n29179, n29181, n29182, n29183, n29184, n29185,
    n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193, n29194,
    n29195, n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203,
    n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211, n29212,
    n29213, n29214, n29215, n29216, n29217, n29218, n29219, n29220, n29221,
    n29222, n29223, n29224, n29225, n29226, n29227, n29228, n29229, n29230,
    n29231, n29232, n29233, n29234, n29235, n29236, n29237, n29238, n29239,
    n29240, n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248,
    n29249, n29250, n29251, n29252, n29253, n29254, n29255, n29257, n29258,
    n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267,
    n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275, n29276,
    n29277, n29278, n29279, n29280, n29281, n29282, n29283, n29284, n29285,
    n29286, n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29294,
    n29295, n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303,
    n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311, n29312,
    n29313, n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
    n29322, n29323, n29324, n29325, n29326, n29327, n29329, n29330, n29331,
    n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339, n29340,
    n29341, n29342, n29343, n29344, n29345, n29346, n29347, n29348, n29349,
    n29350, n29351, n29352, n29353, n29354, n29355, n29356, n29357, n29358,
    n29359, n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367,
    n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375, n29376,
    n29377, n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
    n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394,
    n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403,
    n29404, n29405, n29406, n29408, n29409, n29410, n29411, n29412, n29413,
    n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422,
    n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431,
    n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440,
    n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
    n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458,
    n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467,
    n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476,
    n29477, n29479, n29480, n29481, n29482, n29483, n29484, n29485, n29486,
    n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494, n29495,
    n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29504,
    n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
    n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521, n29522,
    n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531,
    n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539, n29540,
    n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548, n29549,
    n29550, n29551, n29552, n29553, n29554, n29555, n29557, n29558, n29559,
    n29560, n29561, n29562, n29563, n29564, n29565, n29566, n29567, n29568,
    n29569, n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
    n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585, n29586,
    n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595,
    n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603, n29604,
    n29605, n29606, n29607, n29608, n29609, n29610, n29611, n29612, n29613,
    n29614, n29615, n29616, n29617, n29618, n29619, n29620, n29621, n29622,
    n29623, n29624, n29625, n29626, n29627, n29628, n29629, n29630, n29631,
    n29633, n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
    n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649, n29650,
    n29651, n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659,
    n29660, n29661, n29662, n29663, n29664, n29665, n29666, n29667, n29668,
    n29669, n29670, n29671, n29672, n29673, n29674, n29675, n29676, n29677,
    n29678, n29679, n29680, n29681, n29682, n29683, n29684, n29685, n29686,
    n29687, n29688, n29689, n29690, n29691, n29692, n29693, n29694, n29695,
    n29696, n29697, n29698, n29699, n29700, n29701, n29702, n29703, n29704,
    n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713, n29714,
    n29715, n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723,
    n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731, n29732,
    n29733, n29734, n29735, n29736, n29737, n29738, n29739, n29740, n29741,
    n29742, n29743, n29744, n29745, n29746, n29747, n29748, n29749, n29750,
    n29751, n29752, n29753, n29754, n29755, n29756, n29757, n29758, n29759,
    n29760, n29761, n29762, n29763, n29764, n29765, n29766, n29767, n29768,
    n29769, n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777,
    n29778, n29779, n29780, n29781, n29783, n29784, n29785, n29786, n29787,
    n29788, n29789, n29790, n29791, n29792, n29793, n29794, n29795, n29796,
    n29797, n29798, n29799, n29800, n29801, n29802, n29803, n29804, n29805,
    n29806, n29807, n29808, n29809, n29810, n29811, n29812, n29813, n29814,
    n29815, n29816, n29817, n29818, n29819, n29820, n29821, n29822, n29823,
    n29824, n29825, n29826, n29827, n29828, n29829, n29830, n29831, n29832,
    n29833, n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
    n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849, n29850,
    n29851, n29852, n29853, n29854, n29855, n29856, n29857, n29858, n29860,
    n29861, n29862, n29863, n29864, n29865, n29866, n29867, n29868, n29869,
    n29870, n29871, n29872, n29873, n29874, n29875, n29876, n29877, n29878,
    n29879, n29880, n29881, n29882, n29883, n29884, n29885, n29886, n29887,
    n29888, n29889, n29890, n29891, n29892, n29893, n29894, n29895, n29896,
    n29897, n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
    n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913, n29914,
    n29915, n29916, n29917, n29918, n29919, n29920, n29921, n29922, n29923,
    n29924, n29925, n29926, n29927, n29928, n29929, n29930, n29931, n29932,
    n29934, n29935, n29936, n29937, n29938, n29939, n29940, n29941, n29942,
    n29943, n29944, n29945, n29946, n29947, n29948, n29949, n29950, n29951,
    n29952, n29953, n29954, n29955, n29956, n29957, n29958, n29959, n29960,
    n29961, n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
    n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977, n29978,
    n29979, n29980, n29981, n29982, n29983, n29984, n29985, n29986, n29987,
    n29988, n29989, n29990, n29991, n29992, n29993, n29994, n29995, n29996,
    n29997, n29998, n29999, n30000, n30001, n30002, n30003, n30004, n30005,
    n30006, n30007, n30008, n30009, n30010, n30011, n30012, n30014, n30015,
    n30016, n30017, n30018, n30019, n30020, n30021, n30022, n30023, n30024,
    n30025, n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
    n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041, n30042,
    n30043, n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051,
    n30052, n30053, n30054, n30055, n30056, n30057, n30058, n30059, n30060,
    n30061, n30062, n30063, n30064, n30065, n30066, n30067, n30068, n30069,
    n30070, n30071, n30072, n30073, n30074, n30075, n30076, n30077, n30078,
    n30079, n30080, n30081, n30082, n30083, n30084, n30085, n30086, n30087,
    n30089, n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
    n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106,
    n30107, n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115,
    n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123, n30124,
    n30125, n30126, n30127, n30128, n30129, n30130, n30131, n30132, n30133,
    n30134, n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142,
    n30143, n30144, n30145, n30146, n30147, n30148, n30149, n30150, n30151,
    n30152, n30153, n30154, n30155, n30156, n30157, n30158, n30160, n30161,
    n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169, n30170,
    n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178, n30179,
    n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187, n30188,
    n30189, n30190, n30191, n30192, n30193, n30194, n30195, n30196, n30197,
    n30198, n30199, n30200, n30201, n30202, n30203, n30204, n30205, n30206,
    n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214, n30215,
    n30216, n30217, n30218, n30219, n30220, n30221, n30222, n30223, n30224,
    n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233,
    n30234, n30235, n30236, n30237, n30238, n30240, n30241, n30242, n30243,
    n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251, n30252,
    n30253, n30254, n30255, n30256, n30257, n30258, n30259, n30260, n30261,
    n30262, n30263, n30264, n30265, n30266, n30267, n30268, n30269, n30270,
    n30271, n30272, n30273, n30274, n30275, n30276, n30277, n30278, n30279,
    n30280, n30281, n30282, n30283, n30284, n30285, n30286, n30287, n30288,
    n30289, n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297,
    n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305, n30306,
    n30307, n30308, n30309, n30311, n30312, n30313, n30314, n30315, n30316,
    n30317, n30318, n30319, n30320, n30321, n30322, n30323, n30324, n30325,
    n30326, n30327, n30328, n30329, n30330, n30331, n30332, n30333, n30334,
    n30335, n30336, n30337, n30338, n30339, n30340, n30341, n30342, n30343,
    n30344, n30345, n30346, n30347, n30348, n30349, n30350, n30351, n30352,
    n30353, n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
    n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369, n30370,
    n30371, n30372, n30373, n30374, n30375, n30376, n30377, n30378, n30379,
    n30380, n30381, n30382, n30384, n30385, n30386, n30387, n30388, n30389,
    n30390, n30391, n30392, n30393, n30394, n30395, n30396, n30397, n30398,
    n30399, n30400, n30401, n30402, n30403, n30404, n30405, n30406, n30407,
    n30408, n30409, n30410, n30411, n30412, n30413, n30414, n30415, n30416,
    n30417, n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425,
    n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433, n30434,
    n30435, n30436, n30437, n30438, n30439, n30440, n30441, n30442, n30443,
    n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451, n30452,
    n30453, n30454, n30455, n30456, n30457, n30458, n30459, n30460, n30461,
    n30462, n30463, n30464, n30466, n30467, n30468, n30469, n30470, n30471,
    n30472, n30473, n30474, n30475, n30476, n30477, n30478, n30479, n30480,
    n30481, n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489,
    n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497, n30499,
    n30500, n30501, n30502, n30503, n30504, n30505, n30506, n30507, n30508,
    n30509, n30510, n30511, n30512, n30514, n30515, n30516, n30517, n30518,
    n30519, n30520, n30521, n30522, n30523, n30524, n30525, n30526, n30527,
    n30528, n30529, n30530, n30532, n30533, n30534, n30535, n30536, n30537,
    n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545, n30546,
    n30547, n30548, n30549, n30550, n30551, n30552, n30554, n30555, n30556,
    n30557, n30558, n30559, n30560, n30561, n30562, n30563, n30564, n30565,
    n30566, n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574,
    n30575, n30577, n30578, n30579, n30580, n30581, n30582, n30583, n30584,
    n30585, n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593,
    n30594, n30595, n30596, n30597, n30598, n30600, n30601, n30602, n30603,
    n30604, n30605, n30606, n30607, n30608, n30609, n30610, n30611, n30612,
    n30613, n30614, n30615, n30616, n30617, n30618, n30619, n30620, n30621,
    n30623, n30624, n30625, n30626, n30627, n30628, n30629, n30630, n30631,
    n30632, n30633, n30634, n30635, n30636, n30637, n30638, n30639, n30640,
    n30641, n30642, n30643, n30644, n30646, n30647, n30648, n30649, n30650,
    n30651, n30652, n30653, n30654, n30655, n30656, n30657, n30658, n30659,
    n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667, n30669,
    n30670, n30671, n30672, n30673, n30674, n30675, n30676, n30677, n30678,
    n30679, n30680, n30681, n30682, n30683, n30684, n30685, n30686, n30687,
    n30688, n30689, n30690, n30692, n30693, n30694, n30695, n30696, n30697,
    n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705, n30706,
    n30707, n30708, n30709, n30710, n30711, n30712, n30713, n30715, n30716,
    n30717, n30718, n30719, n30720, n30721, n30722, n30723, n30724, n30725,
    n30726, n30727, n30728, n30729, n30730, n30731, n30732, n30733, n30734,
    n30735, n30736, n30738, n30739, n30740, n30741, n30742, n30743, n30744,
    n30745, n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753,
    n30754, n30755, n30756, n30757, n30758, n30759, n30761, n30762, n30763,
    n30764, n30765, n30766, n30767, n30768, n30769, n30770, n30771, n30772,
    n30773, n30774, n30775, n30776, n30777, n30778, n30779, n30780, n30781,
    n30782, n30784, n30785, n30786, n30787, n30788, n30789, n30790, n30791,
    n30792, n30793, n30794, n30795, n30796, n30797, n30798, n30799, n30800,
    n30801, n30802, n30803, n30804, n30805, n30807, n30808, n30809, n30810,
    n30811, n30812, n30813, n30814, n30815, n30816, n30817, n30818, n30819,
    n30820, n30821, n30822, n30823, n30824, n30825, n30826, n30827, n30828,
    n30830, n30831, n30832, n30833, n30834, n30835, n30836, n30837, n30838,
    n30839, n30840, n30841, n30842, n30843, n30844, n30845, n30846, n30847,
    n30848, n30849, n30850, n30851, n30853, n30854, n30855, n30856, n30857,
    n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865, n30866,
    n30867, n30868, n30869, n30870, n30871, n30872, n30873, n30874, n30876,
    n30877, n30878, n30879, n30880, n30881, n30882, n30883, n30884, n30885,
    n30886, n30887, n30888, n30889, n30890, n30891, n30892, n30893, n30894,
    n30895, n30896, n30897, n30899, n30900, n30901, n30902, n30903, n30904,
    n30905, n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913,
    n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30922, n30923,
    n30924, n30925, n30926, n30927, n30928, n30929, n30930, n30931, n30932,
    n30933, n30934, n30935, n30936, n30937, n30938, n30939, n30940, n30941,
    n30942, n30943, n30945, n30946, n30947, n30948, n30949, n30950, n30951,
    n30952, n30953, n30954, n30955, n30956, n30957, n30958, n30959, n30960,
    n30961, n30962, n30963, n30964, n30965, n30966, n30968, n30969, n30970,
    n30971, n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979,
    n30980, n30981, n30982, n30983, n30984, n30985, n30986, n30987, n30988,
    n30989, n30991, n30992, n30993, n30994, n30995, n30996, n30997, n30998,
    n30999, n31000, n31001, n31002, n31003, n31004, n31005, n31006, n31007,
    n31008, n31009, n31010, n31011, n31012, n31014, n31015, n31016, n31017,
    n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025, n31026,
    n31027, n31028, n31029, n31030, n31031, n31032, n31033, n31034, n31035,
    n31037, n31038, n31039, n31040, n31041, n31042, n31043, n31044, n31045,
    n31046, n31047, n31048, n31049, n31050, n31051, n31052, n31053, n31054,
    n31055, n31056, n31057, n31058, n31060, n31061, n31062, n31063, n31064,
    n31065, n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073,
    n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081, n31083,
    n31084, n31085, n31086, n31087, n31088, n31089, n31090, n31091, n31092,
    n31093, n31094, n31095, n31096, n31097, n31098, n31099, n31100, n31101,
    n31102, n31103, n31104, n31106, n31107, n31108, n31109, n31110, n31111,
    n31112, n31113, n31114, n31115, n31116, n31117, n31118, n31119, n31120,
    n31121, n31122, n31123, n31124, n31125, n31126, n31127, n31129, n31130,
    n31131, n31132, n31133, n31134, n31135, n31136, n31137, n31138, n31139,
    n31140, n31141, n31142, n31143, n31144, n31145, n31146, n31147, n31148,
    n31149, n31150, n31152, n31153, n31154, n31155, n31156, n31157, n31158,
    n31159, n31160, n31161, n31162, n31163, n31164, n31165, n31166, n31167,
    n31168, n31169, n31170, n31171, n31172, n31173, n31175, n31176, n31177,
    n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185, n31186,
    n31187, n31188, n31189, n31190, n31191, n31192, n31193, n31194, n31195,
    n31196, n31198, n31199, n31200, n31201, n31202, n31203, n31204, n31205,
    n31206, n31207, n31209, n31210, n31211, n31212, n31214, n31215, n31216,
    n31217, n31219, n31220, n31221, n31222, n31224, n31225, n31226, n31227,
    n31229, n31230, n31231, n31232, n31234, n31235, n31236, n31237, n31239,
    n31240, n31241, n31242, n31244, n31245, n31246, n31247, n31249, n31250,
    n31251, n31252, n31254, n31255, n31256, n31257, n31259, n31260, n31261,
    n31262, n31264, n31265, n31266, n31267, n31269, n31270, n31271, n31272,
    n31274, n31275, n31276, n31277, n31279, n31280, n31281, n31282, n31284,
    n31285, n31286, n31288, n31289, n31290, n31292, n31293, n31294, n31296,
    n31297, n31298, n31300, n31301, n31302, n31304, n31305, n31306, n31308,
    n31309, n31310, n31312, n31313, n31314, n31316, n31317, n31318, n31320,
    n31321, n31322, n31324, n31325, n31326, n31328, n31329, n31330, n31332,
    n31333, n31334, n31336, n31337, n31338, n31340, n31341, n31342, n31344,
    n31345, n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353,
    n31355, n31356, n31357, n31358, n31360, n31361, n31362, n31363, n31365,
    n31366, n31367, n31368, n31370, n31371, n31372, n31373, n31375, n31376,
    n31377, n31378, n31380, n31381, n31382, n31383, n31385, n31386, n31387,
    n31388, n31390, n31391, n31392, n31393, n31395, n31396, n31397, n31398,
    n31400, n31401, n31402, n31403, n31405, n31406, n31407, n31408, n31410,
    n31411, n31412, n31413, n31415, n31416, n31417, n31418, n31420, n31421,
    n31422, n31423, n31425, n31426, n31427, n31428, n31430, n31431, n31432,
    n31433, n31434, n31436, n31437, n31438, n31439, n31441, n31442, n31443,
    n31444, n31446, n31447, n31448, n31449, n31451, n31452, n31453, n31454,
    n31456, n31457, n31458, n31459, n31461, n31462, n31463, n31464, n31466,
    n31467, n31468, n31469, n31471, n31472, n31473, n31474, n31476, n31477,
    n31478, n31479, n31481, n31482, n31483, n31484, n31486, n31487, n31488,
    n31489, n31491, n31492, n31493, n31494, n31496, n31497, n31498, n31499,
    n31501, n31502, n31503, n31504, n31507, n31508, n31509, n31510, n31511,
    n31512, n31513, n31514, n31515, n31516, n31517, n31518, n31520, n31521,
    n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31530, n31531,
    n31532, n31533, n31534, n31535, n31536, n31537, n31538, n31539, n31541,
    n31542, n31543, n31544, n31545, n31546, n31547, n31548, n31549, n31550,
    n31551, n31553, n31554, n31555, n31556, n31557, n31558, n31559, n31560,
    n31561, n31562, n31564, n31565, n31566, n31567, n31568, n31569, n31570,
    n31571, n31572, n31573, n31574, n31576, n31577, n31578, n31579, n31580,
    n31581, n31582, n31583, n31584, n31585, n31587, n31588, n31589, n31590,
    n31591, n31592, n31593, n31594, n31595, n31596, n31597, n31599, n31600,
    n31601, n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
    n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617, n31618,
    n31619, n31620, n31621, n31622, n31623, n31624, n31625, n31626, n31627,
    n31628, n31629, n31630, n31631, n31632, n31633, n31634, n31635, n31636,
    n31637, n31638, n31639, n31640, n31641, n31642, n31643, n31644, n31645,
    n31646, n31647, n31648, n31649, n31650, n31651, n31652, n31653, n31654,
    n31655, n31656, n31657, n31658, n31659, n31660, n31662, n31663, n31664,
    n31665, n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673,
    n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681, n31682,
    n31683, n31684, n31685, n31686, n31687, n31688, n31689, n31690, n31691,
    n31692, n31693, n31694, n31695, n31696, n31697, n31698, n31699, n31700,
    n31701, n31702, n31703, n31705, n31706, n31707, n31708, n31709, n31710,
    n31711, n31712, n31713, n31714, n31715, n31716, n31717, n31718, n31719,
    n31720, n31721, n31722, n31723, n31724, n31725, n31726, n31727, n31728,
    n31729, n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737,
    n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745, n31747,
    n31748, n31749, n31750, n31751, n31752, n31753, n31754, n31755, n31756,
    n31757, n31758, n31759, n31760, n31761, n31762, n31763, n31764, n31765,
    n31766, n31767, n31768, n31769, n31770, n31771, n31772, n31773, n31774,
    n31775, n31776, n31777, n31778, n31779, n31780, n31781, n31782, n31783,
    n31784, n31785, n31786, n31787, n31788, n31790, n31791, n31792, n31793,
    n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801, n31802,
    n31803, n31804, n31805, n31806, n31807, n31808, n31809, n31810, n31811,
    n31812, n31813, n31814, n31815, n31816, n31817, n31818, n31819, n31820,
    n31821, n31822, n31823, n31824, n31825, n31826, n31827, n31828, n31829,
    n31830, n31832, n31833, n31834, n31835, n31836, n31837, n31838, n31839,
    n31840, n31841, n31842, n31843, n31844, n31845, n31846, n31847, n31848,
    n31849, n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857,
    n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865, n31866,
    n31867, n31868, n31869, n31870, n31871, n31872, n31873, n31875, n31876,
    n31877, n31878, n31879, n31880, n31881, n31882, n31883, n31884, n31885,
    n31886, n31887, n31888, n31889, n31890, n31891, n31892, n31893, n31894,
    n31895, n31896, n31897, n31898, n31899, n31900, n31901, n31902, n31903,
    n31904, n31905, n31906, n31907, n31908, n31909, n31910, n31911, n31912,
    n31913, n31914, n31915, n31917, n31918, n31919, n31920, n31921, n31922,
    n31923, n31924, n31925, n31926, n31927, n31928, n31929, n31930, n31931,
    n31932, n31933, n31934, n31935, n31936, n31937, n31938, n31939, n31940,
    n31941, n31942, n31943, n31944, n31945, n31946, n31947, n31948, n31949,
    n31950, n31951, n31952, n31953, n31954, n31955, n31956, n31957, n31958,
    n31960, n31961, n31962, n31963, n31964, n31965, n31966, n31967, n31968,
    n31969, n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977,
    n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985, n31986,
    n31987, n31988, n31989, n31990, n31991, n31992, n31993, n31994, n31995,
    n31996, n31997, n31998, n31999, n32000, n32001, n32002, n32003, n32004,
    n32005, n32006, n32007, n32008, n32009, n32010, n32011, n32012, n32013,
    n32014, n32015, n32016, n32017, n32018, n32019, n32020, n32021, n32022,
    n32023, n32024, n32025, n32026, n32027, n32028, n32029, n32031, n32032,
    n32033, n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
    n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049, n32050,
    n32051, n32052, n32053, n32054, n32055, n32056, n32057, n32058, n32059,
    n32060, n32061, n32062, n32063, n32064, n32065, n32066, n32067, n32068,
    n32069, n32070, n32071, n32072, n32073, n32074, n32076, n32077, n32078,
    n32079, n32080, n32081, n32082, n32083, n32084, n32085, n32086, n32087,
    n32088, n32089, n32090, n32091, n32092, n32093, n32094, n32095, n32096,
    n32097, n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105,
    n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113, n32114,
    n32115, n32116, n32117, n32118, n32120, n32121, n32122, n32123, n32124,
    n32125, n32126, n32127, n32128, n32129, n32130, n32131, n32132, n32133,
    n32134, n32135, n32136, n32137, n32138, n32139, n32140, n32141, n32142,
    n32143, n32144, n32145, n32146, n32147, n32148, n32149, n32150, n32151,
    n32152, n32153, n32154, n32155, n32156, n32157, n32158, n32159, n32160,
    n32161, n32162, n32163, n32165, n32166, n32167, n32168, n32169, n32170,
    n32171, n32172, n32173, n32174, n32175, n32176, n32177, n32178, n32179,
    n32180, n32181, n32182, n32183, n32184, n32185, n32186, n32187, n32188,
    n32189, n32190, n32191, n32192, n32193, n32194, n32195, n32196, n32197,
    n32198, n32199, n32200, n32201, n32202, n32203, n32204, n32205, n32206,
    n32207, n32209, n32210, n32211, n32212, n32213, n32214, n32215, n32216,
    n32217, n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225,
    n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233, n32234,
    n32235, n32236, n32237, n32238, n32239, n32240, n32241, n32242, n32243,
    n32244, n32245, n32246, n32247, n32248, n32249, n32250, n32251, n32252,
    n32254, n32255, n32256, n32257, n32258, n32259, n32260, n32261, n32262,
    n32263, n32264, n32265, n32266, n32267, n32268, n32269, n32270, n32271,
    n32272, n32273, n32274, n32275, n32276, n32277, n32278, n32279, n32280,
    n32281, n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289,
    n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32298, n32299,
    n32300, n32301, n32302, n32303, n32304, n32305, n32306, n32307, n32308,
    n32309, n32310, n32311, n32312, n32313, n32314, n32315, n32316, n32317,
    n32318, n32319, n32320, n32321, n32322, n32323, n32324, n32325, n32326,
    n32327, n32328, n32329, n32330, n32331, n32332, n32333, n32334, n32335,
    n32336, n32337, n32338, n32339, n32340, n32341, n32342, n32343, n32344,
    n32345, n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
    n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361, n32362,
    n32363, n32364, n32365, n32366, n32367, n32368, n32369, n32370, n32371,
    n32372, n32373, n32374, n32375, n32376, n32377, n32378, n32379, n32380,
    n32381, n32382, n32383, n32384, n32385, n32386, n32387, n32388, n32389,
    n32390, n32391, n32392, n32393, n32394, n32395, n32397, n32398, n32399,
    n32400, n32401, n32402, n32403, n32404, n32405, n32406, n32407, n32408,
    n32409, n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
    n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425, n32426,
    n32427, n32428, n32429, n32430, n32431, n32432, n32433, n32434, n32435,
    n32436, n32437, n32438, n32439, n32440, n32441, n32442, n32443, n32445,
    n32446, n32447, n32448, n32449, n32450, n32451, n32452, n32453, n32454,
    n32455, n32456, n32457, n32458, n32459, n32460, n32461, n32462, n32463,
    n32464, n32465, n32466, n32467, n32468, n32469, n32470, n32471, n32472,
    n32473, n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481,
    n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489, n32490,
    n32491, n32492, n32494, n32495, n32496, n32497, n32498, n32499, n32500,
    n32501, n32502, n32503, n32504, n32505, n32506, n32507, n32508, n32509,
    n32510, n32511, n32512, n32513, n32514, n32515, n32516, n32517, n32518,
    n32519, n32520, n32521, n32522, n32523, n32524, n32525, n32526, n32527,
    n32528, n32529, n32530, n32531, n32532, n32533, n32534, n32535, n32536,
    n32537, n32538, n32539, n32540, n32542, n32543, n32544, n32545, n32546,
    n32547, n32548, n32549, n32550, n32551, n32552, n32553, n32554, n32555,
    n32556, n32557, n32558, n32559, n32560, n32561, n32562, n32563, n32564,
    n32565, n32566, n32567, n32568, n32569, n32570, n32571, n32572, n32573,
    n32574, n32575, n32576, n32577, n32578, n32579, n32580, n32581, n32582,
    n32583, n32584, n32585, n32586, n32587, n32588, n32589, n32591, n32592,
    n32593, n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601,
    n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609, n32610,
    n32611, n32612, n32613, n32614, n32615, n32616, n32617, n32618, n32619,
    n32620, n32621, n32622, n32623, n32624, n32625, n32626, n32627, n32628,
    n32629, n32630, n32631, n32632, n32633, n32634, n32635, n32636, n32637,
    n32639, n32640, n32641, n32642, n32643, n32644, n32645, n32646, n32647,
    n32648, n32649, n32650, n32651, n32652, n32653, n32654, n32655, n32656,
    n32657, n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665,
    n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673, n32674,
    n32675, n32676, n32677, n32678, n32679, n32680, n32681, n32682, n32683,
    n32684, n32685, n32686, n32688, n32689, n32690, n32691, n32692, n32693,
    n32694, n32695, n32696, n32697, n32698, n32699, n32700, n32701, n32702,
    n32703, n32704, n32705, n32706, n32707, n32708, n32709, n32710, n32711,
    n32712, n32713, n32714, n32715, n32716, n32717, n32718, n32719, n32720,
    n32721, n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729,
    n32730, n32731, n32732, n32733, n32734, n32736, n32737, n32738, n32739,
    n32740, n32741, n32742, n32743, n32745, n32746, n32747, n32748, n32749,
    n32750, n32751, n32752, n32754, n32755, n32756, n32757, n32758, n32759,
    n32760, n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769,
    n32771, n32772, n32773, n32774, n32775, n32776, n32777, n32778, n32779,
    n32781, n32782, n32783, n32784, n32785, n32786, n32787, n32788, n32790,
    n32791, n32792, n32793, n32794, n32795, n32796, n32797, n32798, n32800,
    n32801, n32802, n32803, n32804, n32805, n32806, n32807, n32809, n32810,
    n32811, n32812, n32813, n32814, n32815, n32816, n32817, n32819, n32820,
    n32821, n32822, n32823, n32824, n32825, n32826, n32828, n32829, n32830,
    n32831, n32832, n32833, n32834, n32835, n32836, n32838, n32839, n32840,
    n32841, n32842, n32843, n32844, n32845, n32847, n32848, n32849, n32850,
    n32851, n32852, n32853, n32854, n32855, n32857, n32858, n32859, n32860,
    n32861, n32862, n32863, n32864, n32866, n32867, n32868, n32869, n32870,
    n32871, n32872, n32873, n32874, n32876, n32877, n32878, n32879, n32880,
    n32881, n32882, n32883, n32885, n32886, n32887, n32888, n32889, n32890,
    n32891, n32892, n32893, n32895, n32896, n32897, n32898, n32899, n32900,
    n32901, n32902, n32904, n32905, n32906, n32907, n32908, n32909, n32910,
    n32911, n32912, n32914, n32915, n32916, n32917, n32918, n32919, n32920,
    n32921, n32923, n32924, n32925, n32926, n32927, n32928, n32929, n32930,
    n32931, n32933, n32934, n32935, n32936, n32937, n32938, n32939, n32940,
    n32942, n32943, n32944, n32945, n32946, n32947, n32948, n32949, n32950,
    n32952, n32953, n32954, n32955, n32956, n32957, n32958, n32959, n32961,
    n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969, n32971,
    n32972, n32973, n32974, n32975, n32976, n32977, n32978, n32980, n32981,
    n32982, n32983, n32984, n32985, n32986, n32987, n32988, n32990, n32991,
    n32992, n32993, n32994, n32995, n32996, n32997, n32999, n33000, n33001,
    n33002, n33003, n33004, n33005, n33006, n33007, n33009, n33010, n33011,
    n33012, n33013, n33014, n33015, n33016, n33018, n33019, n33020, n33021,
    n33022, n33023, n33024, n33025, n33026, n33028, n33029, n33030, n33031,
    n33032, n33033, n33034, n33035, n33037, n33038, n33039, n33040, n33041,
    n33042, n33044, n33045, n33046, n33047, n33048, n33049, n33050, n33051,
    n33052, n33053, n33054, n33055, n33056, n33057, n33058, n33059, n33060,
    n33061, n33062, n33063, n33064, n33065, n33066, n33067, n33068, n33069,
    n33070, n33071, n33072, n33073, n33074, n33075, n33076, n33077, n33078,
    n33079, n33080, n33081, n33082, n33083, n33084, n33085, n33087, n33088,
    n33089, n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097,
    n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105, n33106,
    n33107, n33108, n33110, n33111, n33112, n33113, n33114, n33115, n33116,
    n33117, n33118, n33119, n33120, n33121, n33122, n33123, n33124, n33125,
    n33126, n33127, n33128, n33129, n33130, n33131, n33132, n33133, n33134,
    n33135, n33136, n33137, n33138, n33140, n33141, n33142, n33143, n33144,
    n33145, n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153,
    n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161, n33162,
    n33163, n33164, n33165, n33166, n33167, n33168, n33169, n33171, n33172,
    n33173, n33174, n33175, n33176, n33177, n33178, n33179, n33180, n33181,
    n33182, n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190,
    n33191, n33192, n33193, n33194, n33195, n33196, n33197, n33198, n33199,
    n33200, n33201, n33202, n33203, n33204, n33205, n33206, n33208, n33209,
    n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217, n33218,
    n33219, n33220, n33221, n33222, n33223, n33224, n33225, n33226, n33227,
    n33228, n33229, n33230, n33231, n33232, n33233, n33234, n33235, n33236,
    n33237, n33239, n33240, n33241, n33242, n33243, n33244, n33245, n33246,
    n33247, n33248, n33249, n33250, n33251, n33252, n33253, n33254, n33255,
    n33256, n33257, n33258, n33259, n33260, n33261, n33262, n33263, n33264,
    n33265, n33267, n33268, n33269, n33270, n33271, n33272, n33273, n33274,
    n33275, n33276, n33277, n33278, n33279, n33280, n33281, n33282, n33283,
    n33284, n33285, n33286, n33287, n33288, n33289, n33290, n33291, n33293,
    n33294, n33295, n33296, n33297, n33298, n33299, n33300, n33301, n33302,
    n33303, n33304, n33305, n33306, n33307, n33308, n33309, n33310, n33311,
    n33312, n33313, n33314, n33315, n33316, n33317, n33318, n33319, n33321,
    n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329, n33330,
    n33331, n33332, n33333, n33334, n33335, n33336, n33337, n33338, n33339,
    n33340, n33341, n33342, n33343, n33344, n33345, n33347, n33348, n33349,
    n33350, n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358,
    n33359, n33360, n33361, n33362, n33363, n33364, n33365, n33366, n33367,
    n33368, n33369, n33370, n33371, n33372, n33373, n33375, n33376, n33377,
    n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385, n33386,
    n33387, n33388, n33389, n33390, n33391, n33392, n33393, n33394, n33395,
    n33396, n33397, n33398, n33399, n33401, n33402, n33403, n33404, n33405,
    n33406, n33407, n33408, n33409, n33410, n33411, n33412, n33413, n33414,
    n33415, n33416, n33417, n33418, n33419, n33420, n33421, n33422, n33423,
    n33424, n33425, n33426, n33427, n33429, n33430, n33431, n33432, n33433,
    n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441, n33442,
    n33443, n33444, n33445, n33446, n33447, n33448, n33449, n33450, n33451,
    n33452, n33453, n33455, n33456, n33457, n33458, n33459, n33460, n33461,
    n33462, n33463, n33464, n33465, n33466, n33467, n33468, n33469, n33470,
    n33471, n33472, n33473, n33474, n33475, n33476, n33477, n33478, n33479,
    n33480, n33481, n33483, n33484, n33485, n33486, n33487, n33488, n33489,
    n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497, n33498,
    n33499, n33500, n33501, n33502, n33503, n33504, n33505, n33506, n33507,
    n33509, n33510, n33511, n33512, n33513, n33514, n33515, n33516, n33517,
    n33518, n33519, n33520, n33521, n33522, n33523, n33524, n33525, n33526,
    n33527, n33528, n33529, n33530, n33531, n33532, n33533, n33534, n33535,
    n33537, n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545,
    n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553, n33554,
    n33555, n33556, n33557, n33558, n33559, n33560, n33561, n33563, n33564,
    n33565, n33566, n33567, n33568, n33569, n33570, n33571, n33572, n33573,
    n33574, n33575, n33576, n33577, n33578, n33579, n33580, n33581, n33582,
    n33583, n33584, n33585, n33586, n33587, n33588, n33589, n33591, n33592,
    n33593, n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601,
    n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609, n33610,
    n33611, n33612, n33613, n33614, n33615, n33617, n33618, n33619, n33620,
    n33621, n33622, n33623, n33624, n33625, n33626, n33627, n33628, n33629,
    n33630, n33631, n33632, n33633, n33634, n33635, n33636, n33637, n33638,
    n33639, n33640, n33641, n33642, n33644, n33645, n33646, n33647, n33648,
    n33649, n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657,
    n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665, n33666,
    n33667, n33669, n33670, n33671, n33672, n33673, n33674, n33675, n33676,
    n33677, n33678, n33679, n33680, n33681, n33682, n33683, n33684, n33685,
    n33686, n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694,
    n33696, n33697, n33698, n33699, n33700, n33701, n33702, n33703, n33704,
    n33705, n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713,
    n33714, n33715, n33716, n33717, n33718, n33719, n33721, n33722, n33723,
    n33724, n33725, n33726, n33727, n33728, n33729, n33730, n33731, n33732,
    n33733, n33734, n33735, n33736, n33737, n33738, n33739, n33740, n33741,
    n33742, n33743, n33744, n33745, n33746, n33748, n33749, n33750, n33751,
    n33752, n33753, n33754, n33755, n33756, n33757, n33758, n33759, n33760,
    n33761, n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
    n33770, n33771, n33773, n33774, n33775, n33776, n33777, n33778, n33779,
    n33780, n33781, n33782, n33783, n33784, n33785, n33786, n33787, n33788,
    n33789, n33790, n33791, n33792, n33793, n33794, n33795, n33796, n33797,
    n33798, n33800, n33801, n33802, n33803, n33804, n33805, n33806, n33807,
    n33808, n33809, n33810, n33811, n33812, n33813, n33814, n33815, n33816,
    n33817, n33818, n33819, n33820, n33821, n33822, n33823, n33825, n33826,
    n33827, n33828, n33829, n33830, n33831, n33832, n33833, n33834, n33835,
    n33836, n33837, n33838, n33839, n33840, n33841, n33842, n33843, n33844,
    n33845, n33846, n33847, n33848, n33849, n33850, n33852, n33853, n33854,
    n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862, n33863,
    n33864, n33865, n33866, n33867, n33868, n33869, n33870, n33871, n33872,
    n33873, n33874, n33875, n33877, n33878, n33879, n33880, n33881, n33882,
    n33883, n33884, n33885, n33886, n33887, n33888, n33889, n33890, n33891,
    n33892, n33893, n33894, n33895, n33896, n33897, n33898, n33899, n33900,
    n33902, n33903, n33904, n33905, n33906, n33907, n33908, n33909, n33910,
    n33911, n33912, n33913, n33914, n33915, n33916, n33917, n33918, n33919,
    n33920, n33921, n33922, n33923, n33924, n33925, n33926, n33927, n33929,
    n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937, n33938,
    n33939, n33940, n33941, n33942, n33943, n33944, n33945, n33946, n33947,
    n33948, n33949, n33950, n33951, n33952, n33953, n33954, n33955, n33956,
    n33957, n33958, n33959, n33960, n33961, n33962, n33963, n33964, n33965,
    n33966, n33968, n33969, n33970, n33971, n33972, n33973, n33974, n33975,
    n33977, n33978, n33979, n33981, n33982, n33983, n33985, n33986, n33988,
    n33989, n33990, n33992, n33993, n33995, n33996, n33997, n33998, n34000,
    n34001, n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
    n34010, n34011, n34012, n34013, n34014, n34016, n34017, n34018, n34020,
    n34021, n34023, n34024, n34025, n34027, n34029, n34030, n34031, n34032,
    n34033, n34035, n34036, n34037, n34039, n34040, n34041, n34043, n34044,
    n34046, n34047, n34049, n34050, n34052, n34053, n34054, n34055, n34056,
    n34057, n34059, n34060, n34061, n34062, n34064, n34065, n34066, n34067,
    n34069, n34070, n34071, n34072, n34074, n34075, n34076, n34077, n34079,
    n34080, n34081, n34082, n34084, n34085, n34086, n34087, n34089, n34090,
    n34091, n34092, n34094, n34095, n34096, n34097, n34099, n34100, n34101,
    n34102, n34104, n34105, n34106, n34107, n34109, n34110, n34111, n34112,
    n34114, n34115, n34116, n34117, n34119, n34120, n34121, n34122, n34124,
    n34125, n34126, n34127, n34129, n34130, n34131, n34132, n34134, n34135,
    n34136, n34137, n34139, n34140, n34141, n34142, n34144, n34145, n34146,
    n34147, n34149, n34150, n34151, n34152, n34154, n34155, n34156, n34157,
    n34159, n34160, n34161, n34162, n34164, n34165, n34166, n34167, n34169,
    n34170, n34171, n34172, n34174, n34175, n34176, n34177, n34179, n34180,
    n34181, n34182, n34184, n34185, n34186, n34187, n34189, n34190, n34191,
    n34192, n34194, n34195, n34196, n34197, n34199, n34200, n34201, n34202,
    n34204, n34205, n34206, n34207, n34208, n34209, n34210, n34211, n34212,
    n34213, n34214, n34215, n34216, n34217, n34218, n34219, n34220, n34221,
    n34222, n34223, n34224, n34225, n34226, n34227, n34229, n34230, n34231,
    n34232, n34233, n34234, n34235, n34236, n34237, n34238, n34239, n34240,
    n34241, n34243, n34244, n34245, n34246, n34247, n34248, n34249, n34250,
    n34251, n34253, n34254, n34255, n34256, n34257, n34258, n34260, n34261,
    n34293, n34294, n34295, n34296, n34297, n34298, n34299, n34300, n34301,
    n34302, n34303, n34304, n34305, n34306, n34307, n34308, n34309, n34310,
    n34311, n34312, n34313, n34314, n34315, n34316, n34317, n34318, n34319,
    n34320, n34321, n34322, n34323, n34324, n34325, n34326, n34327, n34328,
    n34329, n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337,
    n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345, n34346,
    n34347, n34348, n34349, n34350, n34351, n34352, n34353, n34354, n34355,
    n34356, n34357, n34358, n34359, n34360, n34361, n34362, n34363, n34364,
    n34365, n34366, n34367, n34368, n34369, n34370, n34371, n34372, n34373,
    n34374, n34375, n34376, n34377, n34378, n34379, n34380, n34381, n34382,
    n34383, n34384, n34385, n34386, n34387, n34388, n34389, n34390, n34391,
    n34392, n34393, n34394, n34395, n34396, n34397, n34398, n34399, n34400,
    n34401, n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409,
    n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417, n34418,
    n34419, n34420, n34421, n34422, n34423, n34424, n34425, n34426, n34427,
    n34428, n34429, n34430, n34431, n34432, n34433, n34434, n34435, n34436,
    n34437, n34438, n34439, n34440, n34441, n34442, n34443, n34444, n34445,
    n34446, n34447, n34448, n34449, n34450, n34451, n34452, n34453, n34454,
    n34455, n34456, n34457, n34458, n34459, n34460, n34461, n34462, n34463,
    n34464, n34465, n34466, n34467, n34468, n34469, n34470, n34471, n34472,
    n34473, n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481,
    n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489, n34490,
    n34491, n34492, n34493, n34494, n34495, n34496, n34497, n34498, n34499,
    n34500, n34501, n34502, n34503, n34504, n34505, n34506, n34507, n34508,
    n34509, n34510, n34511, n34512, n34513, n34514, n34515, n34516, n34517,
    n34518, n34519, n34520, n34521, n34522, n34523, n34524, n34525, n34526,
    n34527, n34528, n34529, n34530, n34531, n34532, n34533, n34534, n34535,
    n34536, n34537, n34538, n34539, n34540, n34541, n34542, n34543, n34544,
    n34545, n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553,
    n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561, n34562,
    n34563, n34564, n34565, n34566, n34567, n34568, n34569, n34570, n34571,
    n34572, n34573, n34574, n34575, n34576, n34577, n34578, n34579, n34580,
    n34581, n34582, n34583, n34584, n34585, n34586, n34587, n34588, n34589,
    n34590, n34591, n34592, n34593, n34594, n34595, n34596, n34597, n34598,
    n34599, n34600, n34601, n34602, n34603, n34604, n34605, n34606, n34607,
    n34608, n34609, n34610, n34611, n34612, n34613, n34614, n34615, n34616,
    n34617, n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625,
    n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633, n34634,
    n34635, n34636, n34637, n34638, n34639, n34640, n34641, n34642, n34643,
    n34644, n34645, n34646, n34647, n34648, n34649, n34650, n34651, n34652,
    n34653, n34654, n34655, n34656, n34657, n34658, n34659, n34660, n34661,
    n34662, n34663, n34664, n34665, n34666, n34667, n34668, n34669, n34670,
    n34671, n34672, n34673, n34674, n34675, n34676, n34677, n34678, n34679,
    n34680, n34681, n34682, n34683, n34684, n34685, n34686, n34687, n34688,
    n34689, n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697,
    n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705, n34706,
    n34707, n34708, n34709, n34710, n34711, n34712, n34713, n34714, n34715,
    n34716, n34717, n34718, n34719, n34720, n34721, n34722, n34723, n34724,
    n34725, n34726, n34727, n34728, n34729, n34730, n34731, n34732, n34733,
    n34734, n34735, n34736, n34737, n34738, n34739, n34740, n34741, n34742,
    n34743, n34744, n34745, n34746, n34747, n34748, n34749, n34750, n34751,
    n34752, n34753, n34754, n34755, n34756, n34757, n34758, n34759, n34760,
    n34761, n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769,
    n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777, n34778,
    n34779, n34780, n34781, n34782, n34783, n34784, n34785, n34786, n34787,
    n34788, n34789, n34790, n34791, n34792, n34793, n34794, n34795, n34796,
    n34797, n34798, n34799, n34800, n34801, n34802, n34803, n34804, n34805,
    n34806, n34807, n34808, n34809, n34810, n34811, n34812, n34813, n34814,
    n34815, n34816, n34817, n34818, n34819, n34820, n34821, n34822, n34823,
    n34824, n34825, n34826, n34827, n34828, n34829, n34830, n34831, n34832,
    n34833, n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841,
    n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849, n34850,
    n34851, n34852, n34853, n34854, n34855, n34856, n34857, n34858, n34859,
    n34860, n34861, n34862, n34863, n34864, n34865, n34866, n34867, n34868,
    n34869, n34870, n34871, n34872, n34873, n34874, n34875, n34876, n34877,
    n34878, n34879, n34880, n34881, n34882, n34883, n34884, n34885, n34886,
    n34887, n34888, n34889, n34890, n34891, n34892, n34893, n34894, n34895,
    n34896, n34897, n34898, n34899, n34900, n34901, n34902, n34903, n34904,
    n34905, n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913,
    n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921, n34922,
    n34923, n34924, n34926, n34927, n34928, n34929, n34930, n34931, n34932,
    n34933, n34935, n34936, n34937, n34938, n34939, n34940, n34941, n34942,
    n34943, n34944, n34945, n34946, n34947, n34948, n34950, n34951, n34952,
    n34953, n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
    n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969, n34970,
    n34971, n34972, n34973, n34974, n34975, n34976, n34977, n34978, n34979,
    n34980, n34981, n34982, n34983, n34984, n34985, n34986, n34987, n34988,
    n34989, n34991, n34992, n34993, n34994, n34995, n34996, n34997, n34998,
    n34999, n35000, n35001, n35002, n35003, n35004, n35005, n35006, n35007,
    n35008, n35009, n35010, n35011, n35012, n35013, n35014, n35015, n35016,
    n35017, n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025,
    n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033, n35034,
    n35035, n35036, n35037, n35038, n35039, n35040, n35041, n35042, n35043,
    n35044, n35045, n35046, n35047, n35048, n35049, n35050, n35051, n35052,
    n35053, n35054, n35055, n35056, n35057, n35058, n35059, n35060, n35061,
    n35062, n35063, n35064, n35065, n35066, n35067, n35068, n35069, n35070,
    n35071, n35072, n35073, n35074, n35075, n35077, n35078, n35079, n35080,
    n35081, n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089,
    n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097, n35099,
    n35100, n35101, n35102, n35103, n35104, n35105, n35106, n35107, n35108,
    n35109, n35110, n35111, n35112, n35113, n35114, n35115, n35116, n35117,
    n35118, n35119, n35121, n35122, n35123, n35124, n35125, n35126, n35127,
    n35128, n35129, n35130, n35131, n35132, n35133, n35134, n35135, n35136,
    n35137, n35138, n35139, n35140, n35141, n35143, n35144, n35145, n35146,
    n35147, n35148, n35149, n35150, n35151, n35152, n35153, n35154, n35155,
    n35156, n35157, n35158, n35159, n35160, n35161, n35162, n35163, n35165,
    n35166, n35167, n35168, n35169, n35170, n35171, n35172, n35173, n35174,
    n35175, n35176, n35177, n35178, n35179, n35180, n35181, n35182, n35183,
    n35184, n35185, n35187, n35188, n35189, n35190, n35191, n35192, n35193,
    n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201, n35202,
    n35203, n35204, n35205, n35206, n35207, n35209, n35210, n35211, n35212,
    n35213, n35214, n35215, n35216, n35217, n35218, n35219, n35220, n35221,
    n35222, n35223, n35224, n35225, n35226, n35227, n35228, n35229, n35231,
    n35232, n35233, n35234, n35235, n35236, n35237, n35238, n35239, n35240,
    n35241, n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249,
    n35250, n35251, n35252, n35253, n35254, n35255, n35257, n35258, n35259,
    n35260, n35261, n35262, n35263, n35264, n35266, n35267, n35268, n35269,
    n35270, n35271, n35272, n35273, n35275, n35276, n35277, n35278, n35279,
    n35280, n35281, n35282, n35284, n35285, n35286, n35287, n35288, n35289,
    n35290, n35291, n35293, n35294, n35295, n35296, n35297, n35298, n35299,
    n35300, n35302, n35303, n35304, n35305, n35306, n35307, n35308, n35309,
    n35311, n35312, n35313, n35314, n35315, n35316, n35317, n35318, n35320,
    n35321, n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
    n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337, n35338,
    n35339, n35340, n35341, n35342, n35343, n35345, n35346, n35347, n35348,
    n35349, n35350, n35351, n35352, n35354, n35355, n35356, n35357, n35358,
    n35359, n35360, n35361, n35363, n35364, n35365, n35366, n35367, n35368,
    n35369, n35370, n35372, n35373, n35374, n35375, n35376, n35377, n35378,
    n35379, n35381, n35382, n35383, n35384, n35385, n35386, n35387, n35388,
    n35390, n35391, n35392, n35393, n35394, n35395, n35396, n35397, n35399,
    n35400, n35401, n35402, n35403, n35404, n35405, n35406, n35408, n35409,
    n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417, n35418,
    n35419, n35420, n35421, n35422, n35423, n35424, n35425, n35426, n35427,
    n35428, n35429, n35430, n35431, n35433, n35434, n35435, n35436, n35437,
    n35438, n35439, n35440, n35442, n35443, n35444, n35445, n35446, n35447,
    n35448, n35449, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
    n35458, n35460, n35461, n35462, n35463, n35464, n35465, n35466, n35467,
    n35469, n35470, n35471, n35472, n35473, n35474, n35475, n35476, n35478,
    n35479, n35480, n35481, n35482, n35483, n35484, n35485, n35487, n35488,
    n35489, n35490, n35491, n35492, n35493, n35494, n35496, n35497, n35498,
    n35499, n35500, n35501, n35502, n35503, n35504, n35505, n35506, n35507,
    n35508, n35509, n35510, n35511, n35512, n35513, n35514, n35515, n35516,
    n35517, n35518, n35519, n35520, n35522, n35523, n35524, n35525, n35526,
    n35527, n35528, n35529, n35531, n35532, n35533, n35534, n35535, n35536,
    n35537, n35538, n35540, n35541, n35542, n35543, n35544, n35545, n35546,
    n35547, n35549, n35550, n35551, n35552, n35553, n35554, n35555, n35556,
    n35558, n35559, n35560, n35561, n35562, n35563, n35564, n35565, n35567,
    n35568, n35569, n35570, n35571, n35572, n35573, n35574, n35576, n35577,
    n35578, n35579, n35580, n35581, n35582, n35583, n35585, n35586, n35587,
    n35588, n35589, n35590, n35591, n35592, n35593, n35594, n35595, n35596,
    n35597, n35598, n35599, n35600, n35601, n35602, n35603, n35604, n35605,
    n35606, n35607, n35609, n35610, n35611, n35612, n35613, n35614, n35615,
    n35616, n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625,
    n35627, n35628, n35629, n35630, n35631, n35632, n35633, n35634, n35636,
    n35637, n35638, n35639, n35640, n35641, n35642, n35643, n35645, n35646,
    n35647, n35648, n35649, n35650, n35651, n35652, n35654, n35655, n35656,
    n35657, n35658, n35659, n35660, n35661, n35663, n35664, n35665, n35666,
    n35667, n35668, n35669, n35670, n35672, n35673, n35674, n35675, n35676,
    n35677, n35678, n35679, n35680, n35681, n35682, n35683, n35684, n35685,
    n35686, n35687, n35688, n35689, n35690, n35691, n35692, n35693, n35695,
    n35696, n35697, n35698, n35699, n35700, n35701, n35702, n35704, n35705,
    n35706, n35707, n35708, n35709, n35710, n35711, n35713, n35714, n35715,
    n35716, n35717, n35718, n35719, n35720, n35722, n35723, n35724, n35725,
    n35726, n35727, n35728, n35729, n35731, n35732, n35733, n35734, n35735,
    n35736, n35737, n35738, n35740, n35741, n35742, n35743, n35744, n35745,
    n35746, n35747, n35749, n35750, n35751, n35752, n35753, n35754, n35755,
    n35756, n35758, n35759, n35760, n35761, n35762, n35763, n35764, n35765,
    n35766, n35767, n35768, n35769, n35770, n35771, n35772, n35773, n35774,
    n35775, n35776, n35777, n35778, n35780, n35781, n35782, n35783, n35784,
    n35785, n35786, n35787, n35789, n35790, n35791, n35792, n35793, n35794,
    n35795, n35796, n35798, n35799, n35800, n35801, n35802, n35803, n35804,
    n35805, n35807, n35808, n35809, n35810, n35811, n35812, n35813, n35814,
    n35816, n35817, n35818, n35819, n35820, n35821, n35822, n35823, n35825,
    n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35834, n35835,
    n35836, n35837, n35838, n35839, n35840, n35841, n35843, n35844, n35845,
    n35846, n35847, n35848, n35849, n35850, n35851, n35852, n35853, n35854,
    n35855, n35856, n35857, n35858, n35859, n35860, n35861, n35862, n35864,
    n35865, n35866, n35867, n35868, n35869, n35870, n35871, n35873, n35874,
    n35875, n35876, n35877, n35878, n35879, n35880, n35882, n35883, n35884,
    n35885, n35886, n35887, n35888, n35889, n35891, n35892, n35893, n35894,
    n35895, n35896, n35897, n35898, n35900, n35901, n35902, n35903, n35904,
    n35905, n35906, n35907, n35909, n35910, n35911, n35912, n35913, n35914,
    n35915, n35916, n35918, n35919, n35920, n35921, n35922, n35923, n35924,
    n35925, n35927, n35928, n35929, n35930, n35931, n35932, n35933, n35934,
    n35935, n35936, n35937, n35938, n35939, n35940, n35941, n35942, n35943,
    n35944, n35945, n35946, n35947, n35948, n35949, n35951, n35952, n35953,
    n35954, n35955, n35956, n35957, n35958, n35960, n35961, n35962, n35963,
    n35964, n35965, n35966, n35967, n35969, n35970, n35971, n35972, n35973,
    n35974, n35975, n35976, n35978, n35979, n35980, n35981, n35982, n35983,
    n35984, n35985, n35987, n35988, n35989, n35990, n35991, n35992, n35993,
    n35994, n35996, n35997, n35998, n35999, n36000, n36001, n36002, n36003,
    n36005, n36006, n36007, n36008, n36009, n36010, n36011, n36012, n36014,
    n36015, n36016, n36017, n36018, n36019, n36020, n36021, n36022, n36023,
    n36024, n36025, n36026, n36027, n36028, n36029, n36030, n36031, n36032,
    n36033, n36034, n36035, n36036, n36038, n36039, n36040, n36041, n36042,
    n36043, n36044, n36045, n36047, n36048, n36049, n36050, n36051, n36052,
    n36053, n36054, n36056, n36057, n36058, n36059, n36060, n36061, n36062,
    n36063, n36065, n36066, n36067, n36068, n36069, n36070, n36071, n36072,
    n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081, n36083,
    n36084, n36085, n36086, n36087, n36088, n36089, n36090, n36092, n36093,
    n36094, n36095, n36096, n36097, n36098, n36099, n36101, n36102, n36103,
    n36104, n36105, n36106, n36107, n36108, n36109, n36110, n36111, n36112,
    n36113, n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121,
    n36123, n36124, n36125, n36126, n36127, n36128, n36129, n36130, n36132,
    n36133, n36134, n36135, n36136, n36137, n36138, n36139, n36141, n36142,
    n36143, n36144, n36145, n36146, n36147, n36148, n36150, n36151, n36152,
    n36153, n36154, n36155, n36156, n36157, n36159, n36160, n36161, n36162,
    n36163, n36164, n36165, n36166, n36168, n36169, n36170, n36171, n36172,
    n36173, n36174, n36175, n36177, n36178, n36179, n36180, n36181, n36182,
    n36183, n36184, n36186, n36187, n36188, n36189, n36190, n36191, n36192,
    n36193, n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201,
    n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209, n36211,
    n36212, n36213, n36214, n36215, n36216, n36217, n36218, n36220, n36221,
    n36222, n36223, n36224, n36225, n36226, n36227, n36229, n36230, n36231,
    n36232, n36233, n36234, n36235, n36236, n36238, n36239, n36240, n36241,
    n36242, n36243, n36244, n36245, n36247, n36248, n36249, n36250, n36251,
    n36252, n36253, n36254, n36256, n36257, n36258, n36259, n36260, n36261,
    n36262, n36263, n36265, n36266, n36267, n36268, n36269, n36270, n36271,
    n36272, n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281,
    n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289, n36290,
    n36291, n36292, n36293, n36295, n36296, n36297, n36298, n36299, n36300,
    n36301, n36302, n36304, n36305, n36306, n36307, n36308, n36309, n36310,
    n36311, n36313, n36314, n36315, n36316, n36317, n36318, n36319, n36320,
    n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329, n36331,
    n36332, n36333, n36334, n36335, n36336, n36337, n36338, n36340, n36341,
    n36342, n36343, n36344, n36345, n36346, n36347, n36349, n36350, n36351,
    n36352, n36353, n36354, n36355, n36356, n36358, n36359, n36360, n36361,
    n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369, n36370,
    n36371, n36372, n36373, n36374, n36375, n36376, n36377, n36379, n36380,
    n36381, n36382, n36383, n36384, n36385, n36386, n36388, n36389, n36390,
    n36391, n36392, n36393, n36394, n36395, n36397, n36398, n36399, n36400,
    n36401, n36402, n36403, n36404, n36406, n36407, n36408, n36409, n36410,
    n36411, n36412, n36413, n36415, n36416, n36417, n36418, n36419, n36420,
    n36421, n36422, n36424, n36425, n36426, n36427, n36428, n36429, n36430,
    n36431, n36433, n36434, n36435, n36436, n36437, n36438, n36439, n36440,
    n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449, n36450,
    n36451, n36452, n36453, n36454, n36455, n36456, n36457, n36458, n36459,
    n36460, n36462, n36463, n36464, n36465, n36466, n36467, n36468, n36469,
    n36471, n36472, n36473, n36474, n36475, n36476, n36477, n36478, n36480,
    n36481, n36482, n36483, n36484, n36485, n36486, n36487, n36489, n36490,
    n36491, n36492, n36493, n36494, n36495, n36496, n36498, n36499, n36500,
    n36501, n36502, n36503, n36504, n36505, n36507, n36508, n36509, n36510,
    n36511, n36512, n36513, n36514, n36516, n36517, n36518, n36519, n36520,
    n36521, n36522, n36523, n36525, n36526, n36527, n36528, n36529, n36530,
    n36531, n36532, n36533, n36534, n36536, n36537, n36538, n36539, n36540,
    n36541, n36543, n36544, n36545, n36546, n36547, n36548, n36549, n36550,
    n36552, n36553, n36554, n36555, n36556, n36557, n36558, n36560, n36561,
    n36562, n36563, n36564, n36565, n36566, n36568, n36569, n36570, n36571,
    n36573, n36574, n36575, n36576, n36577, n36578, n36579, n36580, n36581,
    n36582, n36583, n36584, n36585, n36587, n36588, n36589, n36590, n36591,
    n36592, n36593, n36594, n36595, n36596, n36597, n36598, n36599, n36601,
    n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609, n36610,
    n36611, n36612, n36614, n36615, n36616, n36617, n36618, n36620, n36621,
    n36622, n36623, n36624, n36625, n36626, n36627, n36628, n36629, n36630,
    n36631, n36632, n36633, n36634, n36635, n36636, n36637, n36638, n36639,
    n36640, n36641, n36642, n36643, n36644, n36645, n36646, n36647, n36648,
    n36649, n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657,
    n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665, n36666,
    n36667, n36668, n36669, n36670, n36671, n36672, n36673, n36674, n36675,
    n36676, n36677, n36678, n36679, n36680, n36681, n36682, n36683, n36684,
    n36685, n36686, n36687, n36688, n36689, n36690, n36691, n36692, n36693,
    n36694, n36695, n36696, n36697, n36698, n36699, n36700, n36701, n36702,
    n36703, n36704, n36705, n36706, n36707, n36708, n36709, n36710, n36711,
    n36712, n36713, n36714, n36715, n36716, n36717, n36718, n36719, n36720,
    n36721, n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729,
    n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737, n36738,
    n36739, n36740, n36741, n36742, n36743, n36744, n36745, n36746, n36747,
    n36748, n36749, n36750, n36751, n36752, n36753, n36754, n36755, n36756,
    n36757, n36758, n36759, n36760, n36761, n36762, n36763, n36764, n36765,
    n36766, n36767, n36768, n36769, n36770, n36771, n36772, n36773, n36774,
    n36775, n36776, n36777, n36778, n36779, n36780, n36781, n36782, n36783,
    n36784, n36785, n36786, n36787, n36788, n36789, n36790, n36791, n36792,
    n36793, n36794, n36796, n36797, n36798, n36799, n36800, n36801, n36802,
    n36803, n36804, n36805, n36806, n36807, n36808, n36809, n36810, n36811,
    n36812, n36813, n36814, n36815, n36816, n36817, n36818, n36819, n36820,
    n36821, n36822, n36823, n36824, n36825, n36826, n36827, n36828, n36829,
    n36830, n36831, n36832, n36833, n36834, n36835, n36836, n36837, n36838,
    n36839, n36840, n36841, n36842, n36843, n36844, n36845, n36846, n36847,
    n36848, n36849, n36850, n36851, n36852, n36853, n36854, n36855, n36856,
    n36857, n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865,
    n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873, n36874,
    n36875, n36876, n36877, n36878, n36879, n36880, n36881, n36882, n36883,
    n36884, n36885, n36886, n36887, n36888, n36889, n36890, n36891, n36892,
    n36893, n36894, n36895, n36896, n36897, n36898, n36899, n36900, n36901,
    n36902, n36904, n36905, n36906, n36907, n36908, n36909, n36910, n36911,
    n36912, n36913, n36914, n36915, n36916, n36917, n36918, n36919, n36920,
    n36921, n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929,
    n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937, n36938,
    n36939, n36940, n36941, n36942, n36943, n36944, n36945, n36946, n36947,
    n36948, n36949, n36950, n36951, n36952, n36953, n36954, n36955, n36956,
    n36957, n36958, n36959, n36960, n36961, n36962, n36963, n36964, n36965,
    n36966, n36967, n36968, n36969, n36970, n36971, n36972, n36973, n36974,
    n36975, n36976, n36977, n36978, n36979, n36980, n36981, n36982, n36983,
    n36984, n36985, n36986, n36987, n36988, n36989, n36990, n36991, n36992,
    n36993, n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001,
    n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009, n37010,
    n37011, n37012, n37013, n37014, n37015, n37016, n37017, n37018, n37019,
    n37020, n37021, n37022, n37023, n37025, n37026, n37027, n37028, n37029,
    n37030, n37031, n37032, n37033, n37034, n37035, n37036, n37037, n37038,
    n37039, n37040, n37041, n37042, n37043, n37044, n37045, n37046, n37047,
    n37048, n37049, n37050, n37051, n37052, n37053, n37054, n37055, n37056,
    n37057, n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065,
    n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073, n37074,
    n37075, n37076, n37077, n37078, n37079, n37080, n37081, n37082, n37083,
    n37084, n37085, n37086, n37087, n37088, n37089, n37090, n37091, n37092,
    n37093, n37094, n37095, n37096, n37097, n37098, n37099, n37100, n37101,
    n37102, n37103, n37104, n37105, n37106, n37107, n37108, n37109, n37110,
    n37111, n37112, n37113, n37114, n37115, n37116, n37117, n37118, n37119,
    n37120, n37121, n37122, n37123, n37124, n37125, n37126, n37127, n37128,
    n37129, n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137,
    n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145, n37146,
    n37147, n37148, n37149, n37150, n37151, n37152, n37153, n37154, n37156,
    n37157, n37158, n37159, n37160, n37161, n37162, n37163, n37164, n37165,
    n37166, n37167, n37168, n37169, n37170, n37171, n37172, n37173, n37174,
    n37175, n37176, n37177, n37178, n37179, n37180, n37181, n37182, n37183,
    n37184, n37185, n37186, n37187, n37188, n37189, n37190, n37191, n37192,
    n37193, n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201,
    n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209, n37210,
    n37211, n37212, n37213, n37214, n37215, n37216, n37217, n37218, n37219,
    n37220, n37221, n37222, n37223, n37224, n37225, n37226, n37227, n37228,
    n37229, n37230, n37231, n37232, n37233, n37234, n37235, n37236, n37237,
    n37238, n37239, n37240, n37241, n37242, n37243, n37244, n37245, n37246,
    n37247, n37248, n37249, n37250, n37251, n37252, n37253, n37254, n37255,
    n37256, n37257, n37258, n37259, n37260, n37261, n37262, n37263, n37264,
    n37265, n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273,
    n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281, n37282,
    n37283, n37284, n37285, n37286, n37287, n37288, n37289, n37290, n37292,
    n37293, n37294, n37295, n37296, n37297, n37298, n37299, n37300, n37301,
    n37302, n37303, n37304, n37305, n37306, n37307, n37308, n37309, n37310,
    n37311, n37312, n37313, n37314, n37315, n37316, n37317, n37318, n37319,
    n37320, n37321, n37322, n37323, n37324, n37325, n37326, n37327, n37328,
    n37329, n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337,
    n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345, n37346,
    n37347, n37348, n37349, n37350, n37351, n37352, n37353, n37354, n37355,
    n37356, n37357, n37358, n37359, n37360, n37361, n37362, n37363, n37364,
    n37365, n37366, n37367, n37368, n37369, n37370, n37371, n37372, n37373,
    n37374, n37375, n37376, n37377, n37378, n37379, n37380, n37381, n37382,
    n37383, n37384, n37385, n37386, n37387, n37388, n37389, n37390, n37391,
    n37392, n37393, n37394, n37395, n37396, n37397, n37398, n37399, n37400,
    n37401, n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409,
    n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417, n37418,
    n37419, n37420, n37421, n37422, n37423, n37425, n37426, n37427, n37428,
    n37429, n37430, n37431, n37432, n37433, n37434, n37435, n37436, n37437,
    n37438, n37439, n37440, n37441, n37442, n37443, n37444, n37445, n37446,
    n37447, n37448, n37449, n37450, n37451, n37452, n37453, n37454, n37455,
    n37456, n37457, n37458, n37459, n37460, n37461, n37462, n37463, n37464,
    n37465, n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473,
    n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481, n37482,
    n37483, n37484, n37485, n37486, n37487, n37488, n37489, n37490, n37491,
    n37492, n37493, n37494, n37495, n37496, n37497, n37498, n37499, n37500,
    n37501, n37502, n37503, n37504, n37505, n37506, n37507, n37508, n37509,
    n37510, n37511, n37512, n37513, n37514, n37515, n37516, n37517, n37518,
    n37519, n37520, n37521, n37522, n37523, n37524, n37525, n37526, n37527,
    n37528, n37529, n37530, n37531, n37532, n37533, n37534, n37535, n37536,
    n37537, n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545,
    n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553, n37554,
    n37556, n37557, n37558, n37559, n37560, n37561, n37562, n37563, n37564,
    n37565, n37566, n37567, n37568, n37569, n37570, n37571, n37572, n37573,
    n37574, n37575, n37576, n37577, n37578, n37579, n37580, n37581, n37582,
    n37583, n37584, n37585, n37586, n37587, n37588, n37589, n37590, n37591,
    n37592, n37593, n37594, n37595, n37596, n37597, n37598, n37599, n37600,
    n37601, n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609,
    n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617, n37618,
    n37619, n37620, n37621, n37622, n37623, n37624, n37625, n37626, n37627,
    n37628, n37629, n37630, n37631, n37632, n37633, n37634, n37635, n37636,
    n37637, n37638, n37639, n37640, n37641, n37642, n37643, n37644, n37645,
    n37646, n37647, n37648, n37649, n37650, n37651, n37652, n37654, n37655,
    n37656, n37657, n37658, n37659, n37660, n37661, n37662, n37663, n37664,
    n37665, n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673,
    n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681, n37682,
    n37683, n37684, n37685, n37686, n37687, n37688, n37689, n37690, n37691,
    n37692, n37693, n37694, n37695, n37696, n37697, n37698, n37699, n37700,
    n37701, n37702, n37703, n37704, n37705, n37706, n37707, n37708, n37709,
    n37710, n37711, n37712, n37713, n37714, n37715, n37716, n37717, n37718,
    n37719, n37720, n37721, n37722, n37723, n37724, n37725, n37726, n37727,
    n37728, n37729, n37730, n37731, n37732, n37733, n37734, n37735, n37736,
    n37737, n37738, n37739, n37740, n37741, n37742, n37744, n37745, n37746,
    n37747, n37748, n37749, n37750, n37751, n37752, n37753, n37754, n37755,
    n37756, n37757, n37758, n37759, n37760, n37761, n37762, n37763, n37764,
    n37765, n37766, n37767, n37768, n37769, n37770, n37771, n37772, n37773,
    n37774, n37775, n37776, n37777, n37778, n37779, n37780, n37781, n37782,
    n37783, n37784, n37785, n37786, n37787, n37788, n37789, n37790, n37791,
    n37792, n37793, n37794, n37795, n37796, n37797, n37798, n37799, n37800,
    n37801, n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809,
    n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817, n37818,
    n37819, n37820, n37821, n37822, n37823, n37824, n37825, n37827, n37828,
    n37829, n37830, n37831, n37832, n37833, n37834, n37835, n37836, n37837,
    n37838, n37839, n37840, n37841, n37842, n37843, n37844, n37845, n37846,
    n37847, n37848, n37849, n37850, n37851, n37852, n37853, n37854, n37855,
    n37856, n37857, n37858, n37859, n37860, n37861, n37862, n37863, n37864,
    n37865, n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873,
    n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881, n37882,
    n37883, n37884, n37885, n37886, n37887, n37888, n37889, n37890, n37891,
    n37892, n37893, n37894, n37895, n37896, n37897, n37898, n37899, n37900,
    n37901, n37903, n37904, n37905, n37906, n37907, n37908, n37909, n37910,
    n37911, n37912, n37913, n37914, n37915, n37916, n37917, n37918, n37919,
    n37920, n37921, n37922, n37923, n37924, n37925, n37926, n37927, n37928,
    n37929, n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937,
    n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945, n37946,
    n37947, n37948, n37949, n37950, n37951, n37952, n37953, n37954, n37955,
    n37956, n37957, n37958, n37959, n37960, n37961, n37962, n37963, n37964,
    n37965, n37966, n37967, n37968, n37969, n37970, n37971, n37972, n37973,
    n37975, n37976, n37977, n37978, n37979, n37980, n37981, n37982, n37983,
    n37984, n37985, n37986, n37987, n37988, n37989, n37990, n37991, n37992,
    n37993, n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001,
    n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009, n38010,
    n38011, n38012, n38013, n38014, n38015, n38016, n38017, n38018, n38019,
    n38020, n38021, n38022, n38023, n38024, n38025, n38026, n38027, n38028,
    n38029, n38030, n38031, n38032, n38033, n38034, n38035, n38036, n38037,
    n38038, n38039, n38040, n38041, n38042, n38043, n38044, n38045, n38046,
    n38047, n38048, n38049, n38050, n38051, n38053, n38054, n38055, n38056,
    n38057, n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065,
    n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073, n38074,
    n38075, n38076, n38077, n38078, n38079, n38080, n38081, n38082, n38083,
    n38084, n38085, n38086, n38087, n38088, n38089, n38090, n38091, n38092,
    n38093, n38094, n38095, n38096, n38097, n38098, n38099, n38100, n38101,
    n38102, n38103, n38104, n38105, n38106, n38107, n38108, n38109, n38110,
    n38111, n38112, n38113, n38114, n38115, n38116, n38117, n38118, n38119,
    n38120, n38121, n38122, n38123, n38124, n38125, n38126, n38128, n38129,
    n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137, n38138,
    n38139, n38140, n38141, n38142, n38143, n38144, n38145, n38146, n38147,
    n38148, n38149, n38150, n38151, n38152, n38153, n38154, n38155, n38156,
    n38157, n38158, n38159, n38160, n38161, n38162, n38163, n38164, n38165,
    n38166, n38167, n38168, n38169, n38170, n38171, n38172, n38173, n38174,
    n38175, n38176, n38177, n38178, n38179, n38180, n38181, n38182, n38183,
    n38184, n38185, n38186, n38187, n38188, n38189, n38190, n38191, n38192,
    n38193, n38194, n38195, n38196, n38197, n38198, n38199, n38201, n38202,
    n38203, n38204, n38205, n38206, n38207, n38208, n38209, n38210, n38211,
    n38212, n38213, n38214, n38215, n38216, n38217, n38218, n38219, n38220,
    n38221, n38222, n38223, n38224, n38225, n38226, n38227, n38228, n38229,
    n38230, n38231, n38232, n38233, n38234, n38235, n38236, n38237, n38238,
    n38239, n38240, n38241, n38242, n38243, n38244, n38245, n38246, n38247,
    n38248, n38249, n38250, n38251, n38252, n38253, n38254, n38255, n38256,
    n38257, n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265,
    n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273, n38274,
    n38275, n38276, n38277, n38279, n38280, n38281, n38282, n38283, n38284,
    n38285, n38286, n38287, n38288, n38289, n38290, n38291, n38292, n38293,
    n38294, n38295, n38296, n38297, n38298, n38299, n38300, n38301, n38302,
    n38303, n38304, n38305, n38306, n38307, n38308, n38309, n38310, n38311,
    n38312, n38313, n38314, n38315, n38316, n38317, n38318, n38319, n38320,
    n38321, n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329,
    n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337, n38338,
    n38339, n38340, n38341, n38342, n38343, n38344, n38345, n38346, n38347,
    n38348, n38349, n38351, n38352, n38353, n38354, n38355, n38356, n38357,
    n38358, n38359, n38360, n38361, n38362, n38363, n38364, n38365, n38366,
    n38367, n38368, n38369, n38370, n38371, n38372, n38373, n38374, n38375,
    n38376, n38377, n38378, n38379, n38380, n38381, n38382, n38383, n38384,
    n38385, n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393,
    n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401, n38402,
    n38403, n38404, n38405, n38406, n38407, n38408, n38409, n38410, n38411,
    n38412, n38413, n38414, n38415, n38416, n38417, n38418, n38419, n38420,
    n38421, n38422, n38423, n38424, n38425, n38426, n38427, n38428, n38430,
    n38431, n38432, n38433, n38434, n38435, n38436, n38437, n38438, n38439,
    n38440, n38441, n38442, n38443, n38444, n38445, n38446, n38447, n38448,
    n38449, n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457,
    n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465, n38466,
    n38467, n38468, n38469, n38470, n38471, n38472, n38473, n38474, n38475,
    n38476, n38477, n38478, n38479, n38480, n38481, n38482, n38483, n38484,
    n38485, n38486, n38487, n38488, n38489, n38490, n38491, n38492, n38493,
    n38494, n38495, n38496, n38497, n38498, n38499, n38501, n38502, n38503,
    n38504, n38505, n38506, n38507, n38508, n38509, n38510, n38511, n38512,
    n38513, n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521,
    n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529, n38530,
    n38531, n38532, n38533, n38534, n38535, n38536, n38537, n38538, n38539,
    n38540, n38541, n38542, n38543, n38544, n38545, n38546, n38547, n38548,
    n38549, n38550, n38551, n38552, n38553, n38554, n38555, n38556, n38557,
    n38558, n38559, n38560, n38561, n38562, n38563, n38564, n38565, n38566,
    n38567, n38568, n38569, n38570, n38571, n38572, n38573, n38574, n38575,
    n38576, n38577, n38579, n38580, n38581, n38582, n38583, n38584, n38585,
    n38586, n38587, n38588, n38589, n38590, n38591, n38592, n38593, n38594,
    n38595, n38596, n38597, n38598, n38599, n38600, n38601, n38602, n38603,
    n38604, n38605, n38606, n38607, n38608, n38609, n38610, n38611, n38612,
    n38613, n38614, n38615, n38616, n38617, n38618, n38619, n38620, n38621,
    n38622, n38623, n38624, n38625, n38626, n38627, n38628, n38629, n38630,
    n38631, n38632, n38633, n38634, n38635, n38636, n38637, n38638, n38639,
    n38640, n38641, n38642, n38643, n38644, n38645, n38646, n38647, n38648,
    n38649, n38650, n38651, n38652, n38653, n38655, n38656, n38657, n38658,
    n38659, n38660, n38661, n38662, n38663, n38664, n38665, n38666, n38667,
    n38668, n38669, n38670, n38671, n38672, n38673, n38674, n38675, n38676,
    n38677, n38678, n38679, n38680, n38681, n38682, n38683, n38684, n38685,
    n38686, n38687, n38688, n38689, n38690, n38691, n38692, n38693, n38694,
    n38695, n38696, n38697, n38698, n38699, n38700, n38701, n38702, n38703,
    n38704, n38705, n38706, n38707, n38708, n38709, n38710, n38711, n38712,
    n38713, n38714, n38715, n38716, n38717, n38718, n38719, n38720, n38721,
    n38722, n38723, n38724, n38725, n38726, n38728, n38729, n38730, n38731,
    n38732, n38733, n38734, n38735, n38736, n38737, n38738, n38739, n38740,
    n38741, n38742, n38743, n38744, n38745, n38746, n38747, n38748, n38749,
    n38750, n38751, n38752, n38753, n38754, n38755, n38756, n38757, n38758,
    n38759, n38760, n38761, n38762, n38763, n38764, n38765, n38766, n38767,
    n38768, n38769, n38770, n38771, n38772, n38773, n38774, n38775, n38776,
    n38777, n38778, n38779, n38780, n38781, n38782, n38783, n38784, n38785,
    n38786, n38787, n38788, n38789, n38790, n38791, n38792, n38793, n38794,
    n38795, n38796, n38797, n38798, n38799, n38800, n38801, n38802, n38803,
    n38805, n38806, n38807, n38808, n38809, n38810, n38811, n38812, n38813,
    n38814, n38815, n38816, n38817, n38818, n38819, n38820, n38821, n38822,
    n38823, n38824, n38825, n38826, n38827, n38828, n38829, n38830, n38831,
    n38832, n38833, n38834, n38835, n38836, n38837, n38838, n38839, n38840,
    n38841, n38842, n38843, n38844, n38845, n38846, n38847, n38848, n38849,
    n38850, n38851, n38852, n38853, n38854, n38855, n38856, n38857, n38858,
    n38859, n38860, n38861, n38862, n38863, n38864, n38865, n38866, n38867,
    n38868, n38869, n38870, n38871, n38872, n38873, n38874, n38875, n38876,
    n38877, n38878, n38879, n38880, n38882, n38883, n38884, n38885, n38886,
    n38887, n38888, n38889, n38890, n38891, n38892, n38893, n38894, n38895,
    n38896, n38897, n38898, n38899, n38900, n38901, n38902, n38903, n38904,
    n38905, n38906, n38907, n38908, n38909, n38910, n38911, n38912, n38913,
    n38914, n38915, n38916, n38917, n38918, n38919, n38920, n38921, n38922,
    n38923, n38924, n38925, n38926, n38927, n38928, n38929, n38930, n38931,
    n38932, n38933, n38934, n38935, n38936, n38937, n38938, n38939, n38940,
    n38941, n38942, n38943, n38944, n38945, n38946, n38947, n38948, n38949,
    n38950, n38951, n38952, n38953, n38954, n38956, n38957, n38958, n38959,
    n38960, n38961, n38962, n38963, n38964, n38965, n38966, n38967, n38968,
    n38969, n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977,
    n38978, n38979, n38980, n38981, n38982, n38983, n38984, n38985, n38986,
    n38987, n38988, n38989, n38990, n38991, n38992, n38993, n38994, n38995,
    n38996, n38997, n38998, n38999, n39000, n39001, n39002, n39003, n39004,
    n39005, n39006, n39007, n39008, n39009, n39010, n39011, n39012, n39013,
    n39014, n39015, n39016, n39017, n39018, n39019, n39020, n39021, n39022,
    n39023, n39024, n39025, n39026, n39027, n39028, n39029, n39030, n39031,
    n39032, n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041,
    n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049, n39050,
    n39051, n39052, n39053, n39054, n39055, n39056, n39057, n39058, n39059,
    n39060, n39061, n39062, n39063, n39064, n39065, n39066, n39067, n39068,
    n39069, n39070, n39071, n39072, n39073, n39074, n39075, n39076, n39077,
    n39078, n39079, n39080, n39081, n39082, n39083, n39084, n39085, n39086,
    n39087, n39088, n39089, n39090, n39091, n39092, n39093, n39094, n39095,
    n39096, n39097, n39098, n39099, n39100, n39101, n39102, n39103, n39104,
    n39105, n39106, n39107, n39109, n39110, n39111, n39112, n39113, n39114,
    n39115, n39116, n39117, n39118, n39119, n39120, n39121, n39122, n39123,
    n39124, n39125, n39126, n39127, n39128, n39129, n39130, n39131, n39132,
    n39133, n39134, n39135, n39136, n39137, n39138, n39139, n39140, n39141,
    n39142, n39143, n39144, n39145, n39146, n39147, n39148, n39149, n39150,
    n39151, n39152, n39153, n39154, n39155, n39156, n39157, n39158, n39159,
    n39160, n39161, n39162, n39163, n39164, n39165, n39166, n39167, n39168,
    n39169, n39170, n39171, n39172, n39173, n39174, n39175, n39176, n39177,
    n39178, n39180, n39181, n39182, n39183, n39184, n39185, n39186, n39187,
    n39188, n39189, n39190, n39191, n39192, n39193, n39194, n39195, n39196,
    n39197, n39198, n39199, n39200, n39201, n39202, n39203, n39204, n39205,
    n39206, n39207, n39208, n39209, n39210, n39211, n39212, n39213, n39214,
    n39215, n39216, n39217, n39218, n39219, n39220, n39221, n39222, n39223,
    n39224, n39225, n39226, n39227, n39228, n39229, n39230, n39231, n39232,
    n39233, n39234, n39235, n39236, n39237, n39238, n39239, n39240, n39241,
    n39242, n39243, n39244, n39245, n39246, n39247, n39248, n39249, n39250,
    n39251, n39252, n39253, n39254, n39255, n39256, n39257, n39258, n39260,
    n39261, n39262, n39263, n39264, n39265, n39266, n39267, n39268, n39269,
    n39270, n39271, n39272, n39273, n39274, n39275, n39276, n39277, n39278,
    n39279, n39280, n39281, n39282, n39283, n39284, n39285, n39286, n39287,
    n39288, n39289, n39290, n39291, n39292, n39293, n39294, n39295, n39296,
    n39297, n39298, n39299, n39300, n39301, n39302, n39303, n39304, n39305,
    n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313, n39314,
    n39315, n39316, n39317, n39318, n39319, n39320, n39321, n39322, n39323,
    n39324, n39325, n39326, n39327, n39328, n39329, n39331, n39332, n39333,
    n39334, n39335, n39336, n39337, n39338, n39339, n39340, n39341, n39342,
    n39343, n39344, n39345, n39346, n39347, n39348, n39349, n39350, n39351,
    n39352, n39353, n39354, n39355, n39356, n39357, n39358, n39359, n39360,
    n39361, n39362, n39363, n39364, n39365, n39366, n39367, n39368, n39369,
    n39370, n39371, n39372, n39373, n39374, n39375, n39376, n39377, n39378,
    n39379, n39380, n39381, n39382, n39383, n39384, n39385, n39386, n39387,
    n39388, n39389, n39390, n39391, n39392, n39393, n39394, n39395, n39396,
    n39397, n39398, n39399, n39400, n39401, n39403, n39404, n39405, n39406,
    n39407, n39408, n39409, n39410, n39411, n39412, n39413, n39414, n39415,
    n39416, n39417, n39418, n39419, n39420, n39421, n39422, n39423, n39424,
    n39425, n39426, n39427, n39428, n39429, n39430, n39431, n39432, n39433,
    n39434, n39435, n39436, n39437, n39438, n39439, n39440, n39441, n39442,
    n39443, n39444, n39445, n39446, n39447, n39448, n39449, n39450, n39451,
    n39452, n39453, n39454, n39455, n39456, n39457, n39458, n39459, n39460,
    n39461, n39462, n39463, n39464, n39465, n39466, n39467, n39468, n39469,
    n39470, n39471, n39472, n39473, n39474, n39475, n39476, n39477, n39478,
    n39479, n39480, n39481, n39482, n39483, n39485, n39486, n39487, n39488,
    n39489, n39490, n39491, n39492, n39493, n39494, n39495, n39496, n39497,
    n39498, n39499, n39500, n39501, n39502, n39503, n39504, n39505, n39506,
    n39507, n39508, n39509, n39510, n39511, n39512, n39513, n39514, n39515,
    n39516, n39518, n39519, n39520, n39521, n39522, n39523, n39524, n39525,
    n39526, n39527, n39528, n39529, n39530, n39531, n39533, n39534, n39535,
    n39536, n39537, n39538, n39539, n39540, n39541, n39542, n39543, n39544,
    n39545, n39546, n39547, n39548, n39549, n39551, n39552, n39553, n39554,
    n39555, n39556, n39557, n39558, n39559, n39560, n39561, n39562, n39563,
    n39564, n39565, n39566, n39567, n39568, n39569, n39570, n39571, n39573,
    n39574, n39575, n39576, n39577, n39578, n39579, n39580, n39581, n39582,
    n39583, n39584, n39585, n39586, n39587, n39588, n39589, n39590, n39591,
    n39592, n39593, n39594, n39596, n39597, n39598, n39599, n39600, n39601,
    n39602, n39603, n39604, n39605, n39606, n39607, n39608, n39609, n39610,
    n39611, n39612, n39613, n39614, n39615, n39616, n39617, n39619, n39620,
    n39621, n39622, n39623, n39624, n39625, n39626, n39627, n39628, n39629,
    n39630, n39631, n39632, n39633, n39634, n39635, n39636, n39637, n39638,
    n39639, n39640, n39642, n39643, n39644, n39645, n39646, n39647, n39648,
    n39649, n39650, n39651, n39652, n39653, n39654, n39655, n39656, n39657,
    n39658, n39659, n39660, n39661, n39662, n39663, n39665, n39666, n39667,
    n39668, n39669, n39670, n39671, n39672, n39673, n39674, n39675, n39676,
    n39677, n39678, n39679, n39680, n39681, n39682, n39683, n39684, n39685,
    n39686, n39688, n39689, n39690, n39691, n39692, n39693, n39694, n39695,
    n39696, n39697, n39698, n39699, n39700, n39701, n39702, n39703, n39704,
    n39705, n39706, n39707, n39708, n39709, n39711, n39712, n39713, n39714,
    n39715, n39716, n39717, n39718, n39719, n39720, n39721, n39722, n39723,
    n39724, n39725, n39726, n39727, n39728, n39729, n39730, n39731, n39732,
    n39734, n39735, n39736, n39737, n39738, n39739, n39740, n39741, n39742,
    n39743, n39744, n39745, n39746, n39747, n39748, n39749, n39750, n39751,
    n39752, n39753, n39754, n39755, n39757, n39758, n39759, n39760, n39761,
    n39762, n39763, n39764, n39765, n39766, n39767, n39768, n39769, n39770,
    n39771, n39772, n39773, n39774, n39775, n39776, n39777, n39778, n39780,
    n39781, n39782, n39783, n39784, n39785, n39786, n39787, n39788, n39789,
    n39790, n39791, n39792, n39793, n39794, n39795, n39796, n39797, n39798,
    n39799, n39800, n39801, n39803, n39804, n39805, n39806, n39807, n39808,
    n39809, n39810, n39811, n39812, n39813, n39814, n39815, n39816, n39817,
    n39818, n39819, n39820, n39821, n39822, n39823, n39824, n39826, n39827,
    n39828, n39829, n39830, n39831, n39832, n39833, n39834, n39835, n39836,
    n39837, n39838, n39839, n39840, n39841, n39842, n39843, n39844, n39845,
    n39846, n39847, n39849, n39850, n39851, n39852, n39853, n39854, n39855,
    n39856, n39857, n39858, n39859, n39860, n39861, n39862, n39863, n39864,
    n39865, n39866, n39867, n39868, n39869, n39870, n39872, n39873, n39874,
    n39875, n39876, n39877, n39878, n39879, n39880, n39881, n39882, n39883,
    n39884, n39885, n39886, n39887, n39888, n39889, n39890, n39891, n39892,
    n39893, n39895, n39896, n39897, n39898, n39899, n39900, n39901, n39902,
    n39903, n39904, n39905, n39906, n39907, n39908, n39909, n39910, n39911,
    n39912, n39913, n39914, n39915, n39916, n39918, n39919, n39920, n39921,
    n39922, n39923, n39924, n39925, n39926, n39927, n39928, n39929, n39930,
    n39931, n39932, n39933, n39934, n39935, n39936, n39937, n39938, n39939,
    n39941, n39942, n39943, n39944, n39945, n39946, n39947, n39948, n39949,
    n39950, n39951, n39952, n39953, n39954, n39955, n39956, n39957, n39958,
    n39959, n39960, n39961, n39962, n39964, n39965, n39966, n39967, n39968,
    n39969, n39970, n39971, n39972, n39973, n39974, n39975, n39976, n39977,
    n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985, n39987,
    n39988, n39989, n39990, n39991, n39992, n39993, n39994, n39995, n39996,
    n39997, n39998, n39999, n40000, n40001, n40002, n40003, n40004, n40005,
    n40006, n40007, n40008, n40010, n40011, n40012, n40013, n40014, n40015,
    n40016, n40017, n40018, n40019, n40020, n40021, n40022, n40023, n40024,
    n40025, n40026, n40027, n40028, n40029, n40030, n40031, n40033, n40034,
    n40035, n40036, n40037, n40038, n40039, n40040, n40041, n40042, n40043,
    n40044, n40045, n40046, n40047, n40048, n40049, n40050, n40051, n40052,
    n40053, n40054, n40056, n40057, n40058, n40059, n40060, n40061, n40062,
    n40063, n40064, n40065, n40066, n40067, n40068, n40069, n40070, n40071,
    n40072, n40073, n40074, n40075, n40076, n40077, n40079, n40080, n40081,
    n40082, n40083, n40084, n40085, n40086, n40087, n40088, n40089, n40090,
    n40091, n40092, n40093, n40094, n40095, n40096, n40097, n40098, n40099,
    n40100, n40102, n40103, n40104, n40105, n40106, n40107, n40108, n40109,
    n40110, n40111, n40112, n40113, n40114, n40115, n40116, n40117, n40118,
    n40119, n40120, n40121, n40122, n40123, n40125, n40126, n40127, n40128,
    n40129, n40130, n40131, n40132, n40133, n40134, n40135, n40136, n40137,
    n40138, n40139, n40140, n40141, n40142, n40143, n40144, n40145, n40146,
    n40148, n40149, n40150, n40151, n40152, n40153, n40154, n40155, n40156,
    n40157, n40158, n40159, n40160, n40161, n40162, n40163, n40164, n40165,
    n40166, n40167, n40168, n40169, n40171, n40172, n40173, n40174, n40175,
    n40176, n40177, n40178, n40179, n40180, n40181, n40182, n40183, n40184,
    n40185, n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40194,
    n40195, n40196, n40197, n40198, n40199, n40200, n40201, n40202, n40203,
    n40204, n40205, n40206, n40207, n40208, n40209, n40210, n40211, n40212,
    n40213, n40214, n40215, n40217, n40218, n40219, n40220, n40221, n40222,
    n40223, n40224, n40225, n40226, n40227, n40228, n40229, n40231, n40232,
    n40233, n40234, n40235, n40236, n40237, n40239, n40240, n40241, n40242,
    n40243, n40244, n40245, n40247, n40248, n40249, n40250, n40251, n40252,
    n40253, n40255, n40256, n40257, n40258, n40259, n40260, n40261, n40263,
    n40264, n40265, n40266, n40267, n40268, n40269, n40271, n40272, n40273,
    n40274, n40275, n40276, n40277, n40279, n40280, n40281, n40282, n40283,
    n40284, n40285, n40287, n40288, n40289, n40290, n40292, n40293, n40294,
    n40295, n40297, n40298, n40299, n40300, n40302, n40303, n40304, n40305,
    n40307, n40308, n40309, n40310, n40312, n40313, n40314, n40315, n40317,
    n40318, n40319, n40320, n40322, n40323, n40324, n40325, n40327, n40328,
    n40329, n40331, n40332, n40333, n40335, n40336, n40337, n40339, n40340,
    n40341, n40343, n40344, n40345, n40347, n40348, n40349, n40351, n40352,
    n40353, n40355, n40356, n40357, n40359, n40360, n40361, n40363, n40364,
    n40365, n40367, n40368, n40369, n40371, n40372, n40373, n40375, n40376,
    n40377, n40379, n40380, n40381, n40383, n40384, n40385, n40387, n40388,
    n40389, n40390, n40391, n40392, n40393, n40394, n40395, n40396, n40398,
    n40399, n40400, n40401, n40403, n40404, n40405, n40406, n40408, n40409,
    n40410, n40411, n40413, n40414, n40415, n40416, n40418, n40419, n40420,
    n40421, n40423, n40424, n40425, n40426, n40428, n40429, n40430, n40431,
    n40433, n40434, n40435, n40436, n40438, n40439, n40440, n40441, n40443,
    n40444, n40445, n40446, n40448, n40449, n40450, n40451, n40453, n40454,
    n40455, n40456, n40458, n40459, n40460, n40461, n40463, n40464, n40465,
    n40466, n40468, n40469, n40470, n40471, n40473, n40474, n40475, n40476,
    n40477, n40479, n40480, n40481, n40482, n40484, n40485, n40486, n40487,
    n40489, n40490, n40491, n40492, n40494, n40495, n40496, n40497, n40499,
    n40500, n40501, n40502, n40504, n40505, n40506, n40507, n40509, n40510,
    n40511, n40512, n40514, n40515, n40516, n40517, n40519, n40520, n40521,
    n40522, n40524, n40525, n40526, n40527, n40529, n40530, n40531, n40532,
    n40534, n40535, n40536, n40537, n40539, n40540, n40541, n40542, n40544,
    n40545, n40546, n40547, n40550, n40551, n40552, n40553, n40554, n40555,
    n40556, n40557, n40558, n40559, n40560, n40561, n40563, n40564, n40565,
    n40566, n40567, n40568, n40569, n40570, n40571, n40573, n40574, n40575,
    n40576, n40577, n40578, n40579, n40580, n40581, n40582, n40584, n40585,
    n40586, n40587, n40588, n40589, n40590, n40591, n40592, n40593, n40594,
    n40596, n40597, n40598, n40599, n40600, n40601, n40602, n40603, n40604,
    n40605, n40607, n40608, n40609, n40610, n40611, n40612, n40613, n40614,
    n40615, n40616, n40617, n40619, n40620, n40621, n40622, n40623, n40624,
    n40625, n40626, n40627, n40628, n40630, n40631, n40632, n40633, n40634,
    n40635, n40636, n40637, n40638, n40639, n40640, n40642, n40643, n40644,
    n40645, n40646, n40647, n40648, n40649, n40650, n40651, n40652, n40653,
    n40654, n40655, n40656, n40657, n40658, n40659, n40660, n40661, n40662,
    n40663, n40664, n40665, n40666, n40667, n40668, n40669, n40670, n40671,
    n40672, n40673, n40674, n40675, n40676, n40677, n40678, n40679, n40680,
    n40681, n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689,
    n40690, n40691, n40692, n40693, n40694, n40695, n40696, n40697, n40698,
    n40699, n40700, n40701, n40702, n40703, n40705, n40706, n40707, n40708,
    n40709, n40710, n40711, n40712, n40713, n40714, n40715, n40716, n40717,
    n40718, n40719, n40720, n40721, n40722, n40723, n40724, n40725, n40726,
    n40727, n40728, n40729, n40730, n40731, n40732, n40733, n40734, n40735,
    n40736, n40737, n40738, n40739, n40740, n40741, n40742, n40743, n40744,
    n40745, n40746, n40748, n40749, n40750, n40751, n40752, n40753, n40754,
    n40755, n40756, n40757, n40758, n40759, n40760, n40761, n40762, n40763,
    n40764, n40765, n40766, n40767, n40768, n40769, n40770, n40771, n40772,
    n40773, n40774, n40775, n40776, n40777, n40778, n40779, n40780, n40781,
    n40782, n40783, n40784, n40785, n40786, n40787, n40788, n40790, n40791,
    n40792, n40793, n40794, n40795, n40796, n40797, n40798, n40799, n40800,
    n40801, n40802, n40803, n40804, n40805, n40806, n40807, n40808, n40809,
    n40810, n40811, n40812, n40813, n40814, n40815, n40816, n40817, n40818,
    n40819, n40820, n40821, n40822, n40823, n40824, n40825, n40826, n40827,
    n40828, n40829, n40830, n40831, n40833, n40834, n40835, n40836, n40837,
    n40838, n40839, n40840, n40841, n40842, n40843, n40844, n40845, n40846,
    n40847, n40848, n40849, n40850, n40851, n40852, n40853, n40854, n40855,
    n40856, n40857, n40858, n40859, n40860, n40861, n40862, n40863, n40864,
    n40865, n40866, n40867, n40868, n40869, n40870, n40871, n40872, n40873,
    n40875, n40876, n40877, n40878, n40879, n40880, n40881, n40882, n40883,
    n40884, n40885, n40886, n40887, n40888, n40889, n40890, n40891, n40892,
    n40893, n40894, n40895, n40896, n40897, n40898, n40899, n40900, n40901,
    n40902, n40903, n40904, n40905, n40906, n40907, n40908, n40909, n40910,
    n40911, n40912, n40913, n40914, n40915, n40916, n40918, n40919, n40920,
    n40921, n40922, n40923, n40924, n40925, n40926, n40927, n40928, n40929,
    n40930, n40931, n40932, n40933, n40934, n40935, n40936, n40937, n40938,
    n40939, n40940, n40941, n40942, n40943, n40944, n40945, n40946, n40947,
    n40948, n40949, n40950, n40951, n40952, n40953, n40954, n40955, n40956,
    n40957, n40958, n40960, n40961, n40962, n40963, n40964, n40965, n40966,
    n40967, n40968, n40969, n40970, n40971, n40972, n40973, n40974, n40975,
    n40976, n40977, n40978, n40979, n40980, n40981, n40982, n40983, n40984,
    n40985, n40986, n40987, n40988, n40989, n40990, n40991, n40992, n40993,
    n40994, n40995, n40996, n40997, n40998, n40999, n41000, n41001, n41003,
    n41004, n41005, n41006, n41007, n41008, n41009, n41010, n41011, n41012,
    n41013, n41014, n41015, n41016, n41017, n41018, n41019, n41020, n41021,
    n41022, n41023, n41024, n41025, n41026, n41027, n41028, n41029, n41030,
    n41031, n41032, n41033, n41034, n41035, n41036, n41037, n41038, n41039,
    n41040, n41041, n41042, n41043, n41044, n41045, n41046, n41047, n41048,
    n41049, n41050, n41051, n41052, n41053, n41054, n41055, n41056, n41057,
    n41058, n41059, n41060, n41061, n41062, n41063, n41064, n41065, n41066,
    n41067, n41068, n41069, n41070, n41071, n41072, n41074, n41075, n41076,
    n41077, n41078, n41079, n41080, n41081, n41082, n41083, n41084, n41085,
    n41086, n41087, n41088, n41089, n41090, n41091, n41092, n41093, n41094,
    n41095, n41096, n41097, n41098, n41099, n41100, n41101, n41102, n41103,
    n41104, n41105, n41106, n41107, n41108, n41109, n41110, n41111, n41112,
    n41113, n41114, n41115, n41116, n41117, n41119, n41120, n41121, n41122,
    n41123, n41124, n41125, n41126, n41127, n41128, n41129, n41130, n41131,
    n41132, n41133, n41134, n41135, n41136, n41137, n41138, n41139, n41140,
    n41141, n41142, n41143, n41144, n41145, n41146, n41147, n41148, n41149,
    n41150, n41151, n41152, n41153, n41154, n41155, n41156, n41157, n41158,
    n41159, n41160, n41161, n41163, n41164, n41165, n41166, n41167, n41168,
    n41169, n41170, n41171, n41172, n41173, n41174, n41175, n41176, n41177,
    n41178, n41179, n41180, n41181, n41182, n41183, n41184, n41185, n41186,
    n41187, n41188, n41189, n41190, n41191, n41192, n41193, n41194, n41195,
    n41196, n41197, n41198, n41199, n41200, n41201, n41202, n41203, n41204,
    n41205, n41206, n41208, n41209, n41210, n41211, n41212, n41213, n41214,
    n41215, n41216, n41217, n41218, n41219, n41220, n41221, n41222, n41223,
    n41224, n41225, n41226, n41227, n41228, n41229, n41230, n41231, n41232,
    n41233, n41234, n41235, n41236, n41237, n41238, n41239, n41240, n41241,
    n41242, n41243, n41244, n41245, n41246, n41247, n41248, n41249, n41250,
    n41252, n41253, n41254, n41255, n41256, n41257, n41258, n41259, n41260,
    n41261, n41262, n41263, n41264, n41265, n41266, n41267, n41268, n41269,
    n41270, n41271, n41272, n41273, n41274, n41275, n41276, n41277, n41278,
    n41279, n41280, n41281, n41282, n41283, n41284, n41285, n41286, n41287,
    n41288, n41289, n41290, n41291, n41292, n41293, n41294, n41295, n41297,
    n41298, n41299, n41300, n41301, n41302, n41303, n41304, n41305, n41306,
    n41307, n41308, n41309, n41310, n41311, n41312, n41313, n41314, n41315,
    n41316, n41317, n41318, n41319, n41320, n41321, n41322, n41323, n41324,
    n41325, n41326, n41327, n41328, n41329, n41330, n41331, n41332, n41333,
    n41334, n41335, n41336, n41337, n41338, n41339, n41341, n41342, n41343,
    n41344, n41345, n41346, n41347, n41348, n41349, n41350, n41351, n41352,
    n41353, n41354, n41355, n41356, n41357, n41358, n41359, n41360, n41361,
    n41362, n41363, n41364, n41365, n41366, n41367, n41368, n41369, n41370,
    n41371, n41372, n41373, n41374, n41375, n41376, n41377, n41378, n41379,
    n41380, n41381, n41382, n41383, n41384, n41385, n41386, n41387, n41388,
    n41389, n41390, n41391, n41392, n41393, n41394, n41395, n41396, n41397,
    n41398, n41399, n41400, n41401, n41402, n41403, n41404, n41405, n41406,
    n41407, n41408, n41409, n41410, n41411, n41412, n41413, n41414, n41415,
    n41416, n41417, n41418, n41419, n41420, n41421, n41422, n41423, n41424,
    n41425, n41426, n41427, n41428, n41429, n41430, n41431, n41432, n41433,
    n41434, n41435, n41436, n41437, n41438, n41440, n41441, n41442, n41443,
    n41444, n41445, n41446, n41447, n41448, n41449, n41450, n41451, n41452,
    n41453, n41454, n41455, n41456, n41457, n41458, n41459, n41460, n41461,
    n41462, n41463, n41464, n41465, n41466, n41467, n41468, n41469, n41470,
    n41471, n41472, n41473, n41474, n41475, n41476, n41477, n41478, n41479,
    n41480, n41481, n41482, n41483, n41484, n41485, n41486, n41488, n41489,
    n41490, n41491, n41492, n41493, n41494, n41495, n41496, n41497, n41498,
    n41499, n41500, n41501, n41502, n41503, n41504, n41505, n41506, n41507,
    n41508, n41509, n41510, n41511, n41512, n41513, n41514, n41515, n41516,
    n41517, n41518, n41519, n41520, n41521, n41522, n41523, n41524, n41525,
    n41526, n41527, n41528, n41529, n41530, n41531, n41532, n41533, n41534,
    n41535, n41537, n41538, n41539, n41540, n41541, n41542, n41543, n41544,
    n41545, n41546, n41547, n41548, n41549, n41550, n41551, n41552, n41553,
    n41554, n41555, n41556, n41557, n41558, n41559, n41560, n41561, n41562,
    n41563, n41564, n41565, n41566, n41567, n41568, n41569, n41570, n41571,
    n41572, n41573, n41574, n41575, n41576, n41577, n41578, n41579, n41580,
    n41581, n41582, n41583, n41585, n41586, n41587, n41588, n41589, n41590,
    n41591, n41592, n41593, n41594, n41595, n41596, n41597, n41598, n41599,
    n41600, n41601, n41602, n41603, n41604, n41605, n41606, n41607, n41608,
    n41609, n41610, n41611, n41612, n41613, n41614, n41615, n41616, n41617,
    n41618, n41619, n41620, n41621, n41622, n41623, n41624, n41625, n41626,
    n41627, n41628, n41629, n41630, n41631, n41632, n41634, n41635, n41636,
    n41637, n41638, n41639, n41640, n41641, n41642, n41643, n41644, n41645,
    n41646, n41647, n41648, n41649, n41650, n41651, n41652, n41653, n41654,
    n41655, n41656, n41657, n41658, n41659, n41660, n41661, n41662, n41663,
    n41664, n41665, n41666, n41667, n41668, n41669, n41670, n41671, n41672,
    n41673, n41674, n41675, n41676, n41677, n41678, n41679, n41680, n41682,
    n41683, n41684, n41685, n41686, n41687, n41688, n41689, n41690, n41691,
    n41692, n41693, n41694, n41695, n41696, n41697, n41698, n41699, n41700,
    n41701, n41702, n41703, n41704, n41705, n41706, n41707, n41708, n41709,
    n41710, n41711, n41712, n41713, n41714, n41715, n41716, n41717, n41718,
    n41719, n41720, n41721, n41722, n41723, n41724, n41725, n41726, n41727,
    n41728, n41729, n41731, n41732, n41733, n41734, n41735, n41736, n41737,
    n41738, n41739, n41740, n41741, n41742, n41743, n41744, n41745, n41746,
    n41747, n41748, n41749, n41750, n41751, n41752, n41753, n41754, n41755,
    n41756, n41757, n41758, n41759, n41760, n41761, n41762, n41763, n41764,
    n41765, n41766, n41767, n41768, n41769, n41770, n41771, n41772, n41773,
    n41774, n41775, n41776, n41777, n41779, n41780, n41781, n41782, n41783,
    n41784, n41785, n41786, n41788, n41789, n41790, n41791, n41792, n41793,
    n41794, n41795, n41797, n41798, n41799, n41800, n41801, n41802, n41803,
    n41805, n41806, n41807, n41808, n41809, n41810, n41811, n41812, n41814,
    n41815, n41816, n41817, n41818, n41819, n41820, n41821, n41822, n41824,
    n41825, n41826, n41827, n41828, n41829, n41830, n41831, n41833, n41834,
    n41835, n41836, n41837, n41838, n41839, n41840, n41841, n41843, n41844,
    n41845, n41846, n41847, n41848, n41849, n41850, n41852, n41853, n41854,
    n41855, n41856, n41857, n41858, n41859, n41860, n41862, n41863, n41864,
    n41865, n41866, n41867, n41868, n41869, n41871, n41872, n41873, n41874,
    n41875, n41876, n41877, n41878, n41879, n41881, n41882, n41883, n41884,
    n41885, n41886, n41887, n41888, n41890, n41891, n41892, n41893, n41894,
    n41895, n41896, n41897, n41898, n41900, n41901, n41902, n41903, n41904,
    n41905, n41906, n41907, n41909, n41910, n41911, n41912, n41913, n41914,
    n41915, n41916, n41917, n41919, n41920, n41921, n41922, n41923, n41924,
    n41925, n41926, n41928, n41929, n41930, n41931, n41932, n41933, n41934,
    n41935, n41936, n41938, n41939, n41940, n41941, n41942, n41943, n41944,
    n41945, n41947, n41948, n41949, n41950, n41951, n41952, n41953, n41954,
    n41955, n41957, n41958, n41959, n41960, n41961, n41962, n41963, n41964,
    n41966, n41967, n41968, n41969, n41970, n41971, n41972, n41973, n41974,
    n41976, n41977, n41978, n41979, n41980, n41981, n41982, n41983, n41985,
    n41986, n41987, n41988, n41989, n41990, n41991, n41992, n41993, n41995,
    n41996, n41997, n41998, n41999, n42000, n42001, n42002, n42004, n42005,
    n42006, n42007, n42008, n42009, n42010, n42011, n42012, n42014, n42015,
    n42016, n42017, n42018, n42019, n42020, n42021, n42023, n42024, n42025,
    n42026, n42027, n42028, n42029, n42030, n42031, n42033, n42034, n42035,
    n42036, n42037, n42038, n42039, n42040, n42042, n42043, n42044, n42045,
    n42046, n42047, n42048, n42049, n42050, n42052, n42053, n42054, n42055,
    n42056, n42057, n42058, n42059, n42061, n42062, n42063, n42064, n42065,
    n42066, n42067, n42068, n42069, n42071, n42072, n42073, n42074, n42075,
    n42076, n42077, n42078, n42080, n42081, n42082, n42083, n42084, n42085,
    n42087, n42088, n42089, n42090, n42091, n42092, n42093, n42094, n42095,
    n42096, n42097, n42098, n42099, n42100, n42101, n42102, n42103, n42104,
    n42105, n42106, n42107, n42108, n42109, n42110, n42111, n42112, n42113,
    n42114, n42115, n42116, n42117, n42118, n42119, n42120, n42121, n42122,
    n42123, n42124, n42125, n42126, n42127, n42128, n42130, n42131, n42132,
    n42133, n42134, n42135, n42136, n42137, n42138, n42139, n42140, n42141,
    n42142, n42143, n42144, n42145, n42146, n42147, n42148, n42149, n42150,
    n42151, n42153, n42154, n42155, n42156, n42157, n42158, n42159, n42160,
    n42161, n42162, n42163, n42164, n42165, n42166, n42167, n42168, n42169,
    n42170, n42171, n42172, n42173, n42174, n42175, n42176, n42177, n42178,
    n42179, n42180, n42181, n42183, n42184, n42185, n42186, n42187, n42188,
    n42189, n42190, n42191, n42192, n42193, n42194, n42195, n42196, n42197,
    n42198, n42199, n42200, n42201, n42202, n42203, n42204, n42205, n42206,
    n42207, n42208, n42209, n42210, n42211, n42212, n42214, n42215, n42216,
    n42217, n42218, n42219, n42220, n42221, n42222, n42223, n42224, n42225,
    n42226, n42227, n42228, n42229, n42230, n42231, n42232, n42233, n42234,
    n42235, n42236, n42237, n42238, n42239, n42240, n42241, n42242, n42243,
    n42244, n42245, n42246, n42247, n42248, n42249, n42251, n42252, n42253,
    n42254, n42255, n42256, n42257, n42258, n42259, n42260, n42261, n42262,
    n42263, n42264, n42265, n42266, n42267, n42268, n42269, n42270, n42271,
    n42272, n42273, n42274, n42275, n42276, n42277, n42278, n42279, n42280,
    n42282, n42283, n42284, n42285, n42286, n42287, n42288, n42289, n42290,
    n42291, n42292, n42293, n42294, n42295, n42296, n42297, n42298, n42299,
    n42300, n42301, n42302, n42303, n42304, n42305, n42306, n42307, n42308,
    n42310, n42311, n42312, n42313, n42314, n42315, n42316, n42317, n42318,
    n42319, n42320, n42321, n42322, n42323, n42324, n42325, n42326, n42327,
    n42328, n42329, n42330, n42331, n42332, n42333, n42334, n42336, n42337,
    n42338, n42339, n42340, n42341, n42342, n42343, n42344, n42345, n42346,
    n42347, n42348, n42349, n42350, n42351, n42352, n42353, n42354, n42355,
    n42356, n42357, n42358, n42359, n42360, n42361, n42362, n42364, n42365,
    n42366, n42367, n42368, n42369, n42370, n42371, n42372, n42373, n42374,
    n42375, n42376, n42377, n42378, n42379, n42380, n42381, n42382, n42383,
    n42384, n42385, n42386, n42387, n42388, n42390, n42391, n42392, n42393,
    n42394, n42395, n42396, n42397, n42398, n42399, n42400, n42401, n42402,
    n42403, n42404, n42405, n42406, n42407, n42408, n42409, n42410, n42411,
    n42412, n42413, n42414, n42415, n42416, n42418, n42419, n42420, n42421,
    n42422, n42423, n42424, n42425, n42426, n42427, n42428, n42429, n42430,
    n42431, n42432, n42433, n42434, n42435, n42436, n42437, n42438, n42439,
    n42440, n42441, n42442, n42444, n42445, n42446, n42447, n42448, n42449,
    n42450, n42451, n42452, n42453, n42454, n42455, n42456, n42457, n42458,
    n42459, n42460, n42461, n42462, n42463, n42464, n42465, n42466, n42467,
    n42468, n42469, n42470, n42472, n42473, n42474, n42475, n42476, n42477,
    n42478, n42479, n42480, n42481, n42482, n42483, n42484, n42485, n42486,
    n42487, n42488, n42489, n42490, n42491, n42492, n42493, n42494, n42495,
    n42496, n42498, n42499, n42500, n42501, n42502, n42503, n42504, n42505,
    n42506, n42507, n42508, n42509, n42510, n42511, n42512, n42513, n42514,
    n42515, n42516, n42517, n42518, n42519, n42520, n42521, n42522, n42523,
    n42524, n42526, n42527, n42528, n42529, n42530, n42531, n42532, n42533,
    n42534, n42535, n42536, n42537, n42538, n42539, n42540, n42541, n42542,
    n42543, n42544, n42545, n42546, n42547, n42548, n42549, n42550, n42552,
    n42553, n42554, n42555, n42556, n42557, n42558, n42559, n42560, n42561,
    n42562, n42563, n42564, n42565, n42566, n42567, n42568, n42569, n42570,
    n42571, n42572, n42573, n42574, n42575, n42576, n42577, n42578, n42580,
    n42581, n42582, n42583, n42584, n42585, n42586, n42587, n42588, n42589,
    n42590, n42591, n42592, n42593, n42594, n42595, n42596, n42597, n42598,
    n42599, n42600, n42601, n42602, n42603, n42604, n42606, n42607, n42608,
    n42609, n42610, n42611, n42612, n42613, n42614, n42615, n42616, n42617,
    n42618, n42619, n42620, n42621, n42622, n42623, n42624, n42625, n42626,
    n42627, n42628, n42629, n42630, n42631, n42632, n42634, n42635, n42636,
    n42637, n42638, n42639, n42640, n42641, n42642, n42643, n42644, n42645,
    n42646, n42647, n42648, n42649, n42650, n42651, n42652, n42653, n42654,
    n42655, n42656, n42657, n42658, n42660, n42661, n42662, n42663, n42664,
    n42665, n42666, n42667, n42668, n42669, n42670, n42671, n42672, n42673,
    n42674, n42675, n42676, n42677, n42678, n42679, n42680, n42681, n42682,
    n42683, n42684, n42685, n42687, n42688, n42689, n42690, n42691, n42692,
    n42693, n42694, n42695, n42696, n42697, n42698, n42699, n42700, n42701,
    n42702, n42703, n42704, n42705, n42706, n42707, n42708, n42709, n42710,
    n42712, n42713, n42714, n42715, n42716, n42717, n42718, n42719, n42720,
    n42721, n42722, n42723, n42724, n42725, n42726, n42727, n42728, n42729,
    n42730, n42731, n42732, n42733, n42734, n42735, n42736, n42737, n42739,
    n42740, n42741, n42742, n42743, n42744, n42745, n42746, n42747, n42748,
    n42749, n42750, n42751, n42752, n42753, n42754, n42755, n42756, n42757,
    n42758, n42759, n42760, n42761, n42762, n42764, n42765, n42766, n42767,
    n42768, n42769, n42770, n42771, n42772, n42773, n42774, n42775, n42776,
    n42777, n42778, n42779, n42780, n42781, n42782, n42783, n42784, n42785,
    n42786, n42787, n42788, n42789, n42791, n42792, n42793, n42794, n42795,
    n42796, n42797, n42798, n42799, n42800, n42801, n42802, n42803, n42804,
    n42805, n42806, n42807, n42808, n42809, n42810, n42811, n42812, n42813,
    n42814, n42816, n42817, n42818, n42819, n42820, n42821, n42822, n42823,
    n42824, n42825, n42826, n42827, n42828, n42829, n42830, n42831, n42832,
    n42833, n42834, n42835, n42836, n42837, n42838, n42839, n42840, n42841,
    n42843, n42844, n42845, n42846, n42847, n42848, n42849, n42850, n42851,
    n42852, n42853, n42854, n42855, n42856, n42857, n42858, n42859, n42860,
    n42861, n42862, n42863, n42864, n42865, n42866, n42868, n42869, n42870,
    n42871, n42872, n42873, n42874, n42875, n42876, n42877, n42878, n42879,
    n42880, n42881, n42882, n42883, n42884, n42885, n42886, n42887, n42888,
    n42889, n42890, n42891, n42892, n42893, n42895, n42896, n42897, n42898,
    n42899, n42900, n42901, n42902, n42903, n42904, n42905, n42906, n42907,
    n42908, n42909, n42910, n42911, n42912, n42913, n42914, n42915, n42916,
    n42917, n42918, n42920, n42921, n42922, n42923, n42924, n42925, n42926,
    n42927, n42928, n42929, n42930, n42931, n42932, n42933, n42934, n42935,
    n42936, n42937, n42938, n42939, n42940, n42941, n42942, n42943, n42945,
    n42946, n42947, n42948, n42949, n42950, n42951, n42952, n42953, n42954,
    n42955, n42956, n42957, n42958, n42959, n42960, n42961, n42962, n42963,
    n42964, n42965, n42966, n42967, n42968, n42969, n42970, n42972, n42973,
    n42974, n42975, n42976, n42977, n42978, n42979, n42980, n42981, n42982,
    n42983, n42984, n42985, n42986, n42987, n42988, n42989, n42990, n42991,
    n42992, n42993, n42994, n42995, n42996, n42997, n42998, n42999, n43000,
    n43001, n43002, n43003, n43004, n43005, n43006, n43007, n43008, n43009,
    n43011, n43012, n43013, n43014, n43015, n43016, n43017, n43018, n43020,
    n43021, n43022, n43024, n43025, n43026, n43028, n43029, n43031, n43032,
    n43033, n43035, n43036, n43038, n43039, n43040, n43041, n43043, n43044,
    n43045, n43046, n43047, n43048, n43049, n43050, n43051, n43052, n43053,
    n43054, n43055, n43056, n43057, n43059, n43060, n43061, n43063, n43064,
    n43066, n43067, n43068, n43070, n43072, n43073, n43074, n43075, n43076,
    n43078, n43079, n43080, n43082, n43083, n43084, n43086, n43087, n43089,
    n43090, n43092, n43093, n43095, n43096, n43097, n43098, n43099, n43100,
    n43102, n43103, n43104, n43105, n43107, n43108, n43109, n43110, n43112,
    n43113, n43114, n43115, n43117, n43118, n43119, n43120, n43122, n43123,
    n43124, n43125, n43127, n43128, n43129, n43130, n43132, n43133, n43134,
    n43135, n43137, n43138, n43139, n43140, n43142, n43143, n43144, n43145,
    n43147, n43148, n43149, n43150, n43152, n43153, n43154, n43155, n43157,
    n43158, n43159, n43160, n43162, n43163, n43164, n43165, n43167, n43168,
    n43169, n43170, n43172, n43173, n43174, n43175, n43177, n43178, n43179,
    n43180, n43182, n43183, n43184, n43185, n43187, n43188, n43189, n43190,
    n43192, n43193, n43194, n43195, n43197, n43198, n43199, n43200, n43202,
    n43203, n43204, n43205, n43207, n43208, n43209, n43210, n43212, n43213,
    n43214, n43215, n43217, n43218, n43219, n43220, n43222, n43223, n43224,
    n43225, n43227, n43228, n43229, n43230, n43232, n43233, n43234, n43235,
    n43237, n43238, n43239, n43240, n43242, n43243, n43244, n43245, n43247,
    n43248, n43249, n43250, n43251, n43252, n43253, n43254, n43255, n43256,
    n43257, n43258, n43259, n43260, n43261, n43262, n43263, n43264, n43265,
    n43266, n43267, n43268, n43269, n43270, n43272, n43273, n43274, n43275,
    n43276, n43277, n43278, n43279, n43280, n43281, n43282, n43283, n43284,
    n43286, n43287, n43288, n43289, n43290, n43291, n43292, n43293, n43294,
    n43296, n43297, n43298, n43299, n43300, n43301, n43303, n43304, n43336,
    n43337, n43338, n43339, n43340, n43341, n43342, n43343, n43344, n43345,
    n43346, n43347, n43348, n43349, n43350, n43351, n43352, n43353, n43354,
    n43355, n43356, n43357, n43358, n43359, n43360, n43361, n43362, n43363,
    n43364, n43365, n43366, n43367, n43368, n43369, n43370, n43371, n43372,
    n43373, n43374, n43375, n43376, n43377, n43378, n43379, n43380, n43381,
    n43382, n43383, n43384, n43385, n43386, n43387, n43388, n43389, n43390,
    n43391, n43392, n43393, n43394, n43395, n43396, n43397, n43398, n43399,
    n43400, n43401, n43402, n43403, n43404, n43405, n43406, n43407, n43408,
    n43409, n43410, n43411, n43412, n43413, n43414, n43415, n43416, n43417,
    n43418, n43419, n43420, n43421, n43422, n43423, n43424, n43425, n43426,
    n43427, n43428, n43429, n43430, n43431, n43432, n43433, n43434, n43435,
    n43436, n43437, n43438, n43439, n43440, n43441, n43442, n43443, n43444,
    n43445, n43446, n43447, n43448, n43449, n43450, n43451, n43452, n43453,
    n43454, n43455, n43456, n43457, n43458, n43459, n43460, n43461, n43462,
    n43463, n43464, n43465, n43466, n43467, n43468, n43469, n43470, n43471,
    n43472, n43473, n43474, n43475, n43476, n43477, n43478, n43479, n43480,
    n43481, n43482, n43483, n43484, n43485, n43486, n43487, n43488, n43489,
    n43490, n43491, n43492, n43493, n43494, n43495, n43496, n43497, n43498,
    n43499, n43500, n43501, n43502, n43503, n43504, n43505, n43506, n43507,
    n43508, n43509, n43510, n43511, n43512, n43513, n43514, n43515, n43516,
    n43517, n43518, n43519, n43520, n43521, n43522, n43523, n43524, n43525,
    n43526, n43527, n43528, n43529, n43530, n43531, n43532, n43533, n43534,
    n43535, n43536, n43537, n43538, n43539, n43540, n43541, n43542, n43543,
    n43544, n43545, n43546, n43547, n43548, n43549, n43550, n43551, n43552,
    n43553, n43554, n43555, n43556, n43557, n43558, n43559, n43560, n43561,
    n43562, n43563, n43564, n43565, n43566, n43567, n43568, n43569, n43570,
    n43571, n43572, n43573, n43574, n43575, n43576, n43577, n43578, n43579,
    n43580, n43581, n43582, n43583, n43584, n43585, n43586, n43587, n43588,
    n43589, n43590, n43591, n43592, n43593, n43594, n43595, n43596, n43597,
    n43598, n43599, n43600, n43601, n43602, n43603, n43604, n43605, n43606,
    n43607, n43608, n43609, n43610, n43611, n43612, n43613, n43614, n43615,
    n43616, n43617, n43618, n43619, n43620, n43621, n43622, n43623, n43624,
    n43625, n43626, n43627, n43628, n43629, n43630, n43631, n43632, n43633,
    n43634, n43635, n43636, n43637, n43638, n43639, n43640, n43641, n43642,
    n43643, n43644, n43645, n43646, n43647, n43648, n43649, n43650, n43651,
    n43652, n43653, n43654, n43655, n43656, n43657, n43658, n43659, n43660,
    n43661, n43662, n43663, n43664, n43665, n43666, n43667, n43668, n43669,
    n43670, n43671, n43672, n43673, n43674, n43675, n43676, n43677, n43678,
    n43679, n43680, n43681, n43682, n43683, n43684, n43685, n43686, n43687,
    n43688, n43689, n43690, n43691, n43692, n43693, n43694, n43695, n43696,
    n43697, n43698, n43699, n43700, n43701, n43702, n43703, n43704, n43705,
    n43706, n43707, n43708, n43709, n43710, n43711, n43712, n43713, n43714,
    n43715, n43716, n43717, n43718, n43719, n43720, n43721, n43722, n43723,
    n43724, n43725, n43726, n43727, n43728, n43729, n43730, n43731, n43732,
    n43733, n43734, n43735, n43736, n43737, n43738, n43739, n43740, n43741,
    n43742, n43743, n43744, n43745, n43746, n43747, n43748, n43749, n43750,
    n43751, n43752, n43753, n43754, n43755, n43756, n43757, n43758, n43759,
    n43760, n43761, n43762, n43763, n43764, n43765, n43766, n43767, n43768,
    n43769, n43770, n43771, n43772, n43773, n43774, n43775, n43776, n43777,
    n43778, n43779, n43780, n43781, n43782, n43783, n43784, n43785, n43786,
    n43787, n43788, n43789, n43790, n43791, n43792, n43793, n43794, n43795,
    n43796, n43797, n43798, n43799, n43800, n43801, n43802, n43803, n43804,
    n43805, n43806, n43807, n43808, n43809, n43810, n43811, n43812, n43813,
    n43814, n43815, n43816, n43817, n43818, n43819, n43820, n43821, n43822,
    n43823, n43824, n43825, n43826, n43827, n43828, n43829, n43830, n43831,
    n43832, n43833, n43834, n43835, n43836, n43837, n43838, n43839, n43840,
    n43841, n43842, n43843, n43844, n43845, n43846, n43847, n43848, n43849,
    n43850, n43851, n43852, n43853, n43854, n43855, n43856, n43857, n43858,
    n43859, n43860, n43861, n43862, n43863, n43864, n43865, n43866, n43867,
    n43868, n43869, n43870, n43871, n43872, n43873, n43874, n43875, n43876,
    n43877, n43878, n43879, n43880, n43881, n43882, n43883, n43884, n43885,
    n43886, n43887, n43888, n43889, n43890, n43891, n43892, n43893, n43894,
    n43895, n43896, n43897, n43898, n43899, n43900, n43901, n43902, n43903,
    n43904, n43905, n43906, n43907, n43908, n43909, n43910, n43911, n43912,
    n43913, n43914, n43915, n43916, n43917, n43918, n43919, n43920, n43921,
    n43922, n43923, n43924, n43925, n43926, n43927, n43928, n43929, n43930,
    n43931, n43932, n43933, n43934, n43935, n43936, n43937, n43938, n43939,
    n43940, n43941, n43942, n43943, n43944, n43945, n43946, n43947, n43948,
    n43949, n43950, n43951, n43952, n43953, n43954, n43955, n43956, n43957,
    n43958, n43959, n43960, n43961, n43962, n43963, n43964, n43965, n43966,
    n43967, n43968, n43970, n43971, n43972, n43973, n43974, n43975, n43976,
    n43977, n43979, n43980, n43981, n43982, n43983, n43984, n43985, n43986,
    n43987, n43988, n43989, n43990, n43991, n43992, n43994, n43995, n43996,
    n43997, n43998, n43999, n44000, n44001, n44002, n44003, n44004, n44005,
    n44006, n44007, n44008, n44009, n44010, n44011, n44012, n44013, n44014,
    n44015, n44016, n44017, n44018, n44019, n44020, n44021, n44022, n44023,
    n44024, n44025, n44026, n44027, n44028, n44029, n44030, n44031, n44032,
    n44033, n44035, n44036, n44037, n44038, n44039, n44040, n44041, n44042,
    n44043, n44044, n44045, n44046, n44047, n44048, n44049, n44050, n44051,
    n44052, n44053, n44054, n44055, n44056, n44057, n44058, n44059, n44060,
    n44061, n44062, n44063, n44064, n44065, n44066, n44067, n44068, n44069,
    n44070, n44071, n44072, n44073, n44074, n44075, n44076, n44077, n44078,
    n44079, n44080, n44081, n44082, n44083, n44084, n44085, n44086, n44087,
    n44088, n44089, n44090, n44091, n44092, n44093, n44094, n44095, n44096,
    n44097, n44098, n44099, n44100, n44101, n44102, n44103, n44104, n44105,
    n44106, n44107, n44108, n44109, n44110, n44111, n44112, n44113, n44114,
    n44115, n44116, n44117, n44118, n44119, n44120, n44121, n44122, n44123,
    n44124, n44125, n44126, n44127, n44128, n44129, n44130, n44131, n44132,
    n44133, n44134, n44135, n44136, n44137, n44138, n44139, n44140, n44141,
    n44142, n44143, n44144, n44145, n44146, n44147, n44148, n44149, n44150,
    n44151, n44152, n44153, n44154, n44155, n44156, n44157, n44158, n44159,
    n44160, n44161, n44162, n44163, n44164, n44165, n44166, n44167, n44168,
    n44169, n44170, n44171, n44172, n44173, n44174, n44175, n44176, n44177,
    n44178, n44179, n44180, n44181, n44182, n44183, n44184, n44185, n44186,
    n44187, n44188, n44189, n44190, n44191, n44192, n44193, n44194, n44195,
    n44196, n44197, n44198, n44199, n44200, n44201, n44202, n44203, n44204,
    n44205, n44206, n44207, n44208, n44209, n44210, n44211, n44212, n44213,
    n44214, n44215, n44216, n44217, n44218, n44219, n44220, n44221, n44222,
    n44223, n44224, n44225, n44226, n44227, n44228, n44229, n44230, n44231,
    n44232, n44233, n44234, n44235, n44236, n44237, n44238, n44239, n44240,
    n44241, n44242, n44243, n44244, n44245, n44246, n44247, n44248, n44249,
    n44250, n44251, n44252, n44253, n44254, n44255, n44256, n44257, n44258,
    n44259, n44260, n44261, n44262, n44263, n44264, n44265, n44266, n44267,
    n44268, n44269, n44270, n44271, n44272, n44273, n44274, n44275, n44276,
    n44277, n44278, n44279, n44280, n44281, n44282, n44283, n44284, n44285,
    n44286, n44287, n44288, n44289, n44290, n44291, n44292, n44293, n44294,
    n44295, n44296, n44297, n44298, n44299, n44300, n44301, n44302, n44303,
    n44304, n44305, n44306, n44307, n44308, n44309, n44310, n44311, n44312,
    n44313, n44314, n44315, n44316, n44317, n44318, n44319, n44320, n44321,
    n44322, n44323, n44324, n44325, n44326, n44327, n44328, n44329, n44330,
    n44331, n44332, n44333, n44334, n44335, n44336, n44337, n44338, n44339,
    n44340, n44341, n44342, n44343, n44344, n44345, n44346, n44347, n44348,
    n44349, n44350, n44351, n44352, n44353, n44354, n44355, n44356, n44357,
    n44358, n44359, n44360, n44361, n44362, n44363, n44364, n44365, n44366,
    n44367, n44368, n44369, n44370, n44371, n44372, n44373, n44374, n44375,
    n44376, n44377, n44378, n44379, n44380, n44381, n44382, n44383, n44384,
    n44385, n44386, n44387, n44388, n44389, n44390, n44391, n44392, n44393,
    n44394, n44395, n44396, n44397, n44398, n44399, n44400, n44401, n44402,
    n44403, n44404, n44405, n44406, n44407, n44408, n44409, n44410, n44411,
    n44412, n44413, n44414, n44415, n44416, n44417, n44418, n44419, n44420,
    n44421, n44422, n44423, n44424, n44425, n44426, n44427, n44428, n44429,
    n44430, n44431, n44432, n44433, n44434, n44435, n44436, n44437, n44438,
    n44439, n44440, n44441, n44442, n44443, n44444, n44445, n44446, n44447,
    n44448, n44449, n44450, n44451, n44452, n44453, n44454, n44455, n44456,
    n44457, n44458, n44459, n44460, n44461, n44462, n44463, n44464, n44465,
    n44466, n44467, n44468, n44469, n44470, n44471, n44472, n44473, n44474,
    n44475, n44476, n44477, n44478, n44479, n44480, n44481, n44482, n44483,
    n44484, n44485, n44486, n44487, n44488, n44489, n44490, n44491, n44492,
    n44493, n44494, n44495, n44496, n44497, n44498, n44499, n44500, n44501,
    n44502, n44503, n44504, n44505, n44506, n44507, n44508, n44509, n44510,
    n44511, n44512, n44513, n44514, n44515, n44516, n44517, n44518, n44519,
    n44520, n44521, n44522, n44523, n44524, n44525, n44526, n44527, n44528,
    n44529, n44530, n44531, n44532, n44533, n44534, n44535, n44536, n44537,
    n44538, n44539, n44540, n44541, n44542, n44543, n44544, n44545, n44546,
    n44547, n44548, n44549, n44550, n44551, n44552, n44553, n44554, n44555,
    n44556, n44557, n44558, n44559, n44560, n44561, n44562, n44563, n44564,
    n44565, n44566, n44567, n44568, n44569, n44570, n44571, n44572, n44573,
    n44574, n44575, n44576, n44577, n44578, n44579, n44580, n44581, n44582,
    n44583, n44584, n44585, n44586, n44587, n44588, n44589, n44590, n44591,
    n44592, n44593, n44594, n44595, n44596, n44597, n44598, n44599, n44600,
    n44601, n44602, n44603, n44604, n44605, n44606, n44607, n44608, n44609,
    n44610, n44611, n44612, n44613, n44614, n44615, n44616, n44617, n44618,
    n44619, n44620, n44621, n44622, n44623, n44624, n44625, n44626, n44627,
    n44628, n44629, n44630, n44631, n44632, n44633, n44634, n44635, n44636,
    n44637, n44638, n44639, n44640, n44641, n44642, n44643, n44644, n44645,
    n44646, n44647, n44648, n44649, n44650, n44651, n44652, n44653, n44654,
    n44655, n44656, n44657, n44658, n44659, n44660, n44661, n44662, n44663,
    n44664, n44665, n44666, n44667, n44668, n44669, n44670, n44671, n44672,
    n44673, n44674, n44675, n44676, n44677, n44678, n44679, n44680, n44681,
    n44682, n44683, n44684, n44685, n44686, n44687, n44688, n44689, n44690,
    n44691, n44692, n44693, n44694, n44695, n44696, n44697, n44698, n44699,
    n44700, n44701, n44702, n44703, n44704, n44705, n44706, n44707, n44708,
    n44709, n44710, n44711, n44712, n44713, n44714, n44715, n44716, n44717,
    n44718, n44719, n44720, n44721, n44722, n44723, n44724, n44725, n44726,
    n44727, n44728, n44729, n44730, n44731, n44732, n44733, n44734, n44735,
    n44736, n44737, n44738, n44739, n44740, n44741, n44742, n44743, n44744,
    n44745, n44746, n44747, n44748, n44749, n44750, n44751, n44752, n44753,
    n44754, n44755, n44756, n44757, n44758, n44759, n44760, n44761, n44762,
    n44763, n44764, n44765, n44766, n44767, n44768, n44769, n44770, n44771,
    n44772, n44773, n44774, n44775, n44776, n44777, n44778, n44779, n44780,
    n44781, n44782, n44783, n44784, n44785, n44786, n44787, n44788, n44789,
    n44790, n44791, n44792, n44793, n44794, n44795, n44796, n44797, n44798,
    n44799, n44800, n44801, n44802, n44803, n44804, n44805, n44806, n44807,
    n44808, n44809, n44810, n44811, n44812, n44813, n44814, n44815, n44816,
    n44817, n44818, n44819, n44820, n44821, n44822, n44823, n44824, n44825,
    n44826, n44827, n44828, n44829, n44830, n44831, n44832, n44833, n44834,
    n44835, n44836, n44837, n44838, n44839, n44840, n44841, n44842, n44843,
    n44844, n44845, n44846, n44847, n44848, n44849, n44850, n44851, n44852,
    n44853, n44854, n44855, n44856, n44857, n44858, n44859, n44860, n44861,
    n44862, n44863, n44864, n44865, n44866, n44867, n44868, n44869, n44870,
    n44871, n44872, n44873, n44874, n44875, n44876, n44877, n44878, n44879,
    n44880, n44881, n44882, n44883, n44884, n44885, n44886, n44887, n44888,
    n44889, n44890, n44891, n44892, n44893, n44894, n44895, n44896, n44897,
    n44898, n44899, n44900, n44901, n44902, n44903, n44904, n44905, n44906,
    n44907, n44908, n44909, n44910, n44911, n44912, n44913, n44914, n44915,
    n44916, n44917, n44918, n44919, n44920, n44921, n44922, n44923, n44924,
    n44925, n44926, n44927, n44928, n44929, n44930, n44931, n44932, n44933,
    n44934, n44935, n44936, n44937, n44938, n44939, n44940, n44941, n44942,
    n44943, n44944, n44945, n44946, n44947, n44948, n44949, n44950, n44951,
    n44952, n44953, n44954, n44955, n44956, n44957, n44958, n44959, n44960,
    n44961, n44962, n44963, n44964, n44965, n44966, n44967, n44968, n44969,
    n44970, n44971, n44972, n44973, n44974, n44975, n44976, n44977, n44978,
    n44979, n44980, n44981, n44982, n44983, n44984, n44985, n44986, n44987,
    n44988, n44989, n44990, n44991, n44992, n44993, n44994, n44995, n44996,
    n44997, n44998, n44999, n45000, n45001, n45002, n45003, n45004, n45005,
    n45006, n45007, n45008, n45009, n45010, n45011, n45012, n45013, n45014,
    n45015, n45016, n45017, n45018, n45019, n45020, n45021, n45022, n45023,
    n45024, n45025, n45026, n45027, n45028, n45029, n45030, n45031, n45032,
    n45033, n45034, n45035, n45036, n45037, n45038, n45039, n45040, n45041,
    n45042, n45043, n45044, n45045, n45046, n45047, n45048, n45049, n45050,
    n45051, n45052, n45053, n45054, n45055, n45056, n45057, n45058, n45059,
    n45060, n45061, n45062, n45063, n45064, n45065, n45066, n45067, n45068,
    n45069, n45070, n45071, n45072, n45073, n45074, n45075, n45076, n45077,
    n45078, n45079, n45080, n45081, n45082, n45083, n45084, n45085, n45086,
    n45087, n45088, n45089, n45090, n45091, n45092, n45093, n45094, n45095,
    n45096, n45097, n45098, n45099, n45100, n45101, n45102, n45103, n45104,
    n45105, n45106, n45107, n45108, n45109, n45110, n45111, n45112, n45113,
    n45114, n45115, n45116, n45117, n45118, n45119, n45120, n45121, n45122,
    n45123, n45124, n45125, n45126, n45127, n45128, n45129, n45130, n45131,
    n45132, n45133, n45134, n45135, n45136, n45137, n45138, n45139, n45140,
    n45141, n45142, n45143, n45144, n45145, n45146, n45147, n45148, n45149,
    n45150, n45151, n45152, n45153, n45154, n45155, n45156, n45157, n45158,
    n45159, n45160, n45161, n45162, n45163, n45164, n45165, n45166, n45167,
    n45168, n45169, n45170, n45171, n45172, n45173, n45174, n45175, n45176,
    n45177, n45178, n45179, n45180, n45181, n45182, n45183, n45184, n45185,
    n45186, n45187, n45188, n45189, n45190, n45191, n45192, n45193, n45194,
    n45195, n45196, n45197, n45198, n45199, n45200, n45201, n45202, n45203,
    n45204, n45205, n45206, n45207, n45208, n45209, n45210, n45211, n45212,
    n45213, n45214, n45215, n45216, n45217, n45218, n45219, n45220, n45221,
    n45222, n45223, n45224, n45225, n45226, n45227, n45228, n45229, n45230,
    n45231, n45232, n45233, n45234, n45235, n45236, n45237, n45238, n45239,
    n45240, n45241, n45242, n45243, n45244, n45245, n45246, n45247, n45248,
    n45249, n45250, n45251, n45252, n45253, n45254, n45255, n45256, n45257,
    n45258, n45259, n45260, n45261, n45262, n45263, n45264, n45265, n45266,
    n45267, n45268, n45269, n45270, n45271, n45272, n45273, n45274, n45275,
    n45276, n45277, n45278, n45279, n45280, n45281, n45282, n45283, n45284,
    n45285, n45286, n45287, n45288, n45289, n45290, n45291, n45292, n45293,
    n45294, n45295, n45296, n45297, n45298, n45299, n45300, n45301, n45302,
    n45303, n45304, n45305, n45306, n45307, n45308, n45309, n45310, n45311,
    n45312, n45313, n45314, n45315, n45316, n45317, n45318, n45319, n45320,
    n45321, n45322, n45323, n45324, n45325, n45326, n45327, n45328, n45329,
    n45330, n45331, n45332, n45333, n45334, n45335, n45336, n45337, n45338,
    n45339, n45340, n45341, n45342, n45343, n45344, n45345, n45346, n45347,
    n45348, n45349, n45350, n45351, n45352, n45353, n45354, n45355, n45356,
    n45357, n45358, n45359, n45360, n45361, n45362, n45363, n45364, n45365,
    n45366, n45367, n45368, n45369, n45370, n45371, n45372, n45373, n45374,
    n45375, n45376, n45377, n45378, n45379, n45380, n45381, n45382, n45383,
    n45384, n45385, n45386, n45387, n45388, n45389, n45390, n45391, n45392,
    n45393, n45394, n45395, n45396, n45397, n45398, n45399, n45400, n45401,
    n45402, n45403, n45404, n45405, n45406, n45407, n45408, n45409, n45410,
    n45411, n45412, n45413, n45414, n45415, n45416, n45417, n45418, n45419,
    n45420, n45421, n45422, n45423, n45424, n45425, n45426, n45427, n45428,
    n45429, n45430, n45431, n45432, n45433, n45434, n45435, n45436, n45437,
    n45438, n45439, n45440, n45441, n45442, n45443, n45444, n45445, n45446,
    n45447, n45448, n45449, n45450, n45451, n45452, n45453, n45454, n45455,
    n45456, n45457, n45458, n45459, n45460, n45461, n45462, n45463, n45464,
    n45465, n45466, n45467, n45468, n45469, n45470, n45471, n45472, n45473,
    n45474, n45475, n45476, n45477, n45478, n45479, n45480, n45481, n45482,
    n45483, n45484, n45485, n45486, n45487, n45488, n45489, n45490, n45491,
    n45492, n45493, n45494, n45495, n45496, n45497, n45498, n45499, n45500,
    n45501, n45502, n45503, n45504, n45505, n45506, n45507, n45508, n45509,
    n45510, n45511, n45512, n45513, n45514, n45515, n45516, n45517, n45518,
    n45519, n45520, n45521, n45522, n45523, n45524, n45525, n45526, n45527,
    n45528, n45529, n45530, n45531, n45532, n45533, n45534, n45535, n45536,
    n45537, n45538, n45539, n45540, n45541, n45542, n45543, n45544, n45545,
    n45546, n45547, n45548, n45549, n45550, n45551, n45552, n45553, n45554,
    n45555, n45556, n45557, n45558, n45559, n45560, n45561, n45562, n45563,
    n45564, n45565, n45566, n45567, n45568, n45569, n45570, n45571, n45572,
    n45573, n45574, n45575, n45576, n45577, n45578, n45579, n45580, n45581,
    n45582, n45583, n45584, n45585, n45586, n45587, n45588, n45589, n45590,
    n45591, n45592, n45593, n45594, n45595, n45596, n45597, n45598, n45599,
    n45600, n45601, n45602, n45603, n45604, n45605, n45606, n45607, n45608,
    n45609, n45610, n45611, n45612, n45613, n45614, n45615, n45616, n45617,
    n45618, n45619, n45620, n45621, n45622, n45623, n45624, n45625, n45626,
    n45627, n45628, n45629, n45630, n45631, n45632, n45633, n45634, n45635,
    n45636, n45637, n45638, n45639, n45640, n45641, n45642, n45643, n45644,
    n45645, n45646, n45647, n45648, n45649, n45650, n45651, n45652, n45653,
    n45654, n45655, n45656, n45657, n45658, n45659, n45660, n45661, n45662,
    n45663, n45664, n45665, n45666, n45667, n45668, n45669, n45670, n45671,
    n45672, n45673, n45674, n45675, n45676, n45677, n45678, n45679, n45680,
    n45681, n45682, n45683, n45684, n45685, n45686, n45687, n45688, n45689,
    n45690, n45691, n45692, n45693, n45694, n45695, n45696, n45697, n45698,
    n45699, n45700, n45701, n45702, n45703, n45704, n45705, n45706, n45707,
    n45708, n45709, n45710, n45711, n45712, n45713, n45714, n45715, n45716,
    n45717, n45718, n45719, n45720, n45721, n45722, n45723, n45724, n45725,
    n45726, n45727, n45728, n45729, n45730, n45731, n45732, n45733, n45734,
    n45735, n45736, n45737, n45738, n45739, n45740, n45741, n45742, n45743,
    n45744, n45745, n45746, n45747, n45748, n45749, n45750, n45751, n45752,
    n45753, n45754, n45755, n45756, n45757, n45758, n45759, n45760, n45761,
    n45762, n45763, n45764, n45765, n45766, n45767, n45768, n45769, n45770,
    n45771, n45772, n45773, n45774, n45775, n45776, n45777, n45778, n45779,
    n45780, n45781, n45782, n45783, n45784, n45785, n45786, n45787, n45788,
    n45789, n45790, n45791, n45792, n45793, n45794, n45795, n45796, n45797,
    n45798, n45799, n45800, n45801, n45802, n45803, n45804, n45805, n45806,
    n45807, n45808, n45809, n45810, n45811, n45812, n45813, n45814, n45815,
    n45816, n45817, n45818, n45819, n45820, n45821, n45822, n45823, n45824,
    n45825, n45826, n45827, n45828, n45829, n45830, n45831, n45832, n45833,
    n45834, n45835, n45836, n45837, n45838, n45839, n45840, n45841, n45842,
    n45843, n45844, n45845, n45846, n45847, n45848, n45849, n45850, n45851,
    n45852, n45853, n45854, n45855, n45856, n45857, n45858, n45859, n45860,
    n45861, n45862, n45863, n45864, n45865, n45866, n45867, n45868, n45869,
    n45870, n45871, n45872, n45873, n45874, n45875, n45876, n45877, n45878,
    n45879, n45880, n45881, n45882, n45883, n45884, n45885, n45886, n45887,
    n45888, n45889, n45890, n45891, n45892, n45893, n45894, n45895, n45896,
    n45897, n45898, n45899, n45900, n45901, n45902, n45903, n45904, n45905,
    n45906, n45907, n45908, n45909, n45910, n45911, n45912, n45913, n45914,
    n45915, n45916, n45917, n45918, n45919, n45920, n45921, n45922, n45923,
    n45924, n45925, n45926, n45927, n45928, n45929, n45930, n45931, n45932,
    n45933, n45934, n45935, n45936, n45937, n45938, n45939, n45940, n45941,
    n45942, n45943, n45944, n45945, n45946, n45947, n45948, n45949, n45950,
    n45951, n45952, n45953, n45954, n45955, n45956, n45957, n45958, n45959,
    n45960, n45961, n45962, n45963, n45964, n45965, n45966, n45967, n45968,
    n45969, n45970, n45971, n45972, n45973, n45974, n45975, n45976, n45977,
    n45978, n45979, n45980, n45981, n45982, n45983, n45984, n45985, n45986,
    n45987, n45988, n45989, n45990, n45991, n45992, n45993, n45994, n45995,
    n45996, n45997, n45998, n45999, n46000, n46001, n46002, n46003, n46004,
    n46005, n46006, n46007, n46008, n46009, n46010, n46011, n46012, n46013,
    n46014, n46015, n46016, n46017, n46018, n46019, n46020, n46021, n46022,
    n46023, n46024, n46025, n46026, n46027, n46028, n46029, n46030, n46031,
    n46032, n46033, n46034, n46035, n46036, n46037, n46038, n46039, n46040,
    n46041, n46042, n46043, n46044, n46045, n46046, n46047, n46048, n46049,
    n46050, n46051, n46052, n46053, n46054, n46055, n46056, n46057, n46058,
    n46059, n46060, n46061, n46062, n46063, n46064, n46065, n46066, n46067,
    n46068, n46069, n46070, n46071, n46072, n46073, n46074, n46075, n46076,
    n46077, n46078, n46079, n46080, n46081, n46082, n46083, n46084, n46085,
    n46086, n46087, n46088, n46089, n46090, n46091, n46092, n46093, n46094,
    n46095, n46096, n46097, n46098, n46099, n46100, n46101, n46102, n46103,
    n46104, n46105, n46106, n46107, n46108, n46109, n46110, n46111, n46112,
    n46113, n46114, n46115, n46116, n46117, n46118, n46119, n46120, n46121,
    n46122, n46123, n46124, n46125, n46126, n46127, n46128, n46129, n46130,
    n46131, n46132, n46133, n46134, n46135, n46136, n46137, n46138, n46139,
    n46140, n46141, n46142, n46143, n46144, n46145, n46146, n46147, n46148,
    n46149, n46150, n46151, n46152, n46153, n46154, n46155, n46156, n46157,
    n46158, n46159, n46160, n46161, n46162, n46163, n46164, n46165, n46166,
    n46167, n46168, n46169, n46170, n46171, n46172, n46173, n46174, n46175,
    n46176, n46177, n46178, n46179, n46180, n46181, n46182, n46183, n46184,
    n46185, n46186, n46187, n46188, n46189, n46190, n46191, n46192, n46193,
    n46194, n46195, n46196, n46197, n46198, n46199, n46200, n46201, n46202,
    n46203, n46204, n46205, n46206, n46207, n46208, n46209, n46210, n46211,
    n46212, n46213, n46214, n46215, n46216, n46217, n46218, n46219, n46220,
    n46221, n46222, n46223, n46224, n46225, n46226, n46227, n46228, n46229,
    n46230, n46231, n46232, n46233, n46234, n46235, n46236, n46237, n46238,
    n46239, n46240, n46241, n46242, n46243, n46244, n46245, n46246, n46247,
    n46248, n46249, n46250, n46251, n46252, n46253, n46254, n46255, n46256,
    n46257, n46258, n46259, n46260, n46261, n46262, n46263, n46264, n46265,
    n46266, n46267, n46268, n46269, n46270, n46271, n46272, n46273, n46274,
    n46275, n46276, n46277, n46278, n46279, n46280, n46281, n46282, n46283,
    n46284, n46285, n46286, n46287, n46288, n46289, n46290, n46291, n46292,
    n46293, n46294, n46295, n46296, n46297, n46298, n46299, n46300, n46301,
    n46302, n46303, n46304, n46305, n46306, n46307, n46308, n46309, n46310,
    n46311, n46312, n46313, n46314, n46315, n46316, n46317, n46318, n46319,
    n46320, n46321, n46322, n46323, n46324, n46325, n46326, n46327, n46328,
    n46329, n46330, n46331, n46332, n46333, n46334, n46335, n46336, n46337,
    n46338, n46339, n46340, n46341, n46342, n46343, n46344, n46345, n46346,
    n46347, n46348, n46349, n46350, n46351, n46352, n46353, n46354, n46355,
    n46356, n46357, n46358, n46359, n46360, n46361, n46362, n46363, n46364,
    n46365, n46366, n46367, n46368, n46369, n46370, n46371, n46372, n46373,
    n46374, n46375, n46376, n46377, n46378, n46379, n46380, n46381, n46382,
    n46383, n46384, n46385, n46386, n46387, n46388, n46389, n46390, n46391,
    n46392, n46393, n46394, n46395, n46396, n46397, n46398, n46399, n46400,
    n46401, n46402, n46403, n46404, n46405, n46406, n46407, n46408, n46409,
    n46410, n46411, n46412, n46413, n46414, n46415, n46416, n46417, n46418,
    n46419, n46420, n46421, n46422, n46423, n46424, n46425, n46426, n46427,
    n46428, n46429, n46430, n46431, n46432, n46433, n46434, n46435, n46436,
    n46437, n46438, n46439, n46440, n46441, n46442, n46443, n46444, n46445,
    n46446, n46447, n46448, n46449, n46450, n46451, n46452, n46453, n46454,
    n46455, n46456, n46457, n46458, n46459, n46460, n46461, n46462, n46463,
    n46464, n46465, n46466, n46467, n46468, n46469, n46470, n46471, n46472,
    n46473, n46474, n46475, n46476, n46477, n46478, n46479, n46480, n46481,
    n46482, n46483, n46484, n46485, n46486, n46487, n46488, n46489, n46490,
    n46491, n46492, n46493, n46494, n46495, n46496, n46497, n46498, n46499,
    n46500, n46501, n46502, n46503, n46504, n46505, n46506, n46507, n46508,
    n46509, n46510, n46511, n46512, n46513, n46514, n46515, n46516, n46517,
    n46518, n46519, n46520, n46521, n46522, n46523, n46524, n46525, n46526,
    n46527, n46528, n46529, n46530, n46531, n46532, n46533, n46534, n46535,
    n46536, n46537, n46538, n46539, n46540, n46541, n46542, n46543, n46544,
    n46545, n46546, n46547, n46548, n46549, n46550, n46551, n46552, n46553,
    n46554, n46555, n46556, n46557, n46558, n46559, n46560, n46561, n46562,
    n46563, n46564, n46565, n46566, n46567, n46568, n46569, n46570, n46571,
    n46572, n46573, n46574, n46575, n46576, n46577, n46578, n46579, n46580,
    n46581, n46582, n46583, n46584, n46585, n46586, n46587, n46588, n46589,
    n46590, n46591, n46592, n46593, n46594, n46595, n46596, n46597, n46598,
    n46599, n46600, n46601, n46602, n46603, n46604, n46605, n46606, n46607,
    n46608, n46609, n46610, n46611, n46612, n46613, n46614, n46615, n46616,
    n46617, n46618, n46619, n46620, n46621, n46622, n46623, n46624, n46625,
    n46626, n46627, n46628, n46629, n46630, n46631, n46632, n46633, n46634,
    n46635, n46636, n46637, n46638, n46639, n46640, n46641, n46642, n46643,
    n46644, n46645, n46646, n46647, n46648, n46649, n46650, n46651, n46652,
    n46653, n46654, n46655, n46656, n46657, n46658, n46659, n46660, n46661,
    n46662, n46663, n46664, n46665, n46666, n46667, n46668, n46669, n46670,
    n46671, n46672, n46673, n46674, n46675, n46676, n46677, n46678, n46679,
    n46680, n46681, n46682, n46683, n46684, n46685, n46686, n46687, n46688,
    n46689, n46690, n46691, n46692, n46693, n46694, n46695, n46696, n46697,
    n46698, n46699, n46700, n46701, n46702, n46703, n46704, n46705, n46706,
    n46707, n46708, n46709, n46710, n46711, n46712, n46713, n46714, n46715,
    n46716, n46717, n46718, n46719, n46720, n46721, n46722, n46723, n46724,
    n46725, n46726, n46727, n46728, n46729, n46730, n46731, n46732, n46733,
    n46734, n46735, n46736, n46737, n46738, n46739, n46740, n46741, n46742,
    n46743, n46744, n46745, n46746, n46747, n46748, n46749, n46750, n46751,
    n46752, n46753, n46754, n46755, n46756, n46757, n46758, n46759, n46760,
    n46761, n46762, n46763, n46764, n46765, n46766, n46767, n46768, n46769,
    n46770, n46771, n46772, n46773, n46774, n46775, n46776, n46777, n46778,
    n46779, n46780, n46781, n46782, n46783, n46784, n46785, n46786, n46787,
    n46788, n46789, n46790, n46791, n46792, n46793, n46794, n46795, n46796,
    n46797, n46798, n46799, n46800, n46801, n46802, n46803, n46804, n46805,
    n46806, n46807, n46808, n46809, n46810, n46811, n46812, n46813, n46814,
    n46815, n46816, n46817, n46818, n46819, n46820, n46821, n46822, n46823,
    n46824, n46825, n46826, n46827, n46828, n46829, n46830, n46831, n46832,
    n46833, n46834, n46835, n46836, n46837, n46838, n46839, n46840, n46841,
    n46842, n46843, n46844, n46845, n46846, n46847, n46848, n46849, n46850,
    n46851, n46852, n46853, n46854, n46855, n46856, n46857, n46858, n46859,
    n46860, n46861, n46862, n46863, n46864, n46865, n46866, n46867, n46868,
    n46869, n46870, n46871, n46872, n46873, n46874, n46875, n46876, n46877,
    n46878, n46879, n46880, n46881, n46882, n46883, n46884, n46885, n46886,
    n46887, n46888, n46889, n46890, n46891, n46892, n46893, n46894, n46895,
    n46896, n46897, n46898, n46899, n46900, n46901, n46902, n46903, n46904,
    n46905, n46906, n46907, n46908, n46909, n46910, n46911, n46912, n46913,
    n46914, n46915, n46916, n46917, n46918, n46919, n46920, n46921, n46922,
    n46923, n46924, n46925, n46926, n46927, n46928, n46929, n46930, n46931,
    n46932, n46933, n46934, n46935, n46936, n46937, n46938, n46939, n46940,
    n46941, n46942, n46943, n46944, n46945, n46946, n46947, n46948, n46949,
    n46950, n46951, n46952, n46953, n46954, n46955, n46956, n46957, n46958,
    n46959, n46960, n46961, n46962, n46963, n46964, n46965, n46966, n46967,
    n46968, n46969, n46970, n46971, n46972, n46973, n46974, n46975, n46976,
    n46977, n46978, n46979, n46980, n46981, n46982, n46983, n46984, n46985,
    n46986, n46987, n46988, n46989, n46990, n46991, n46992, n46993, n46994,
    n46995, n46996, n46997, n46998, n46999, n47000, n47001, n47002, n47003,
    n47004, n47005, n47006, n47007, n47008, n47009, n47010, n47011, n47012,
    n47013, n47014, n47015, n47016, n47017, n47018, n47019, n47020, n47021,
    n47022, n47023, n47024, n47025, n47026, n47027, n47028, n47029, n47030,
    n47031, n47032, n47033, n47034, n47035, n47036, n47037, n47038, n47039,
    n47040, n47041, n47042, n47043, n47044, n47045, n47046, n47047, n47048,
    n47049, n47050, n47051, n47052, n47053, n47054, n47055, n47056, n47057,
    n47058, n47059, n47060, n47061, n47062, n47063, n47064, n47065, n47066,
    n47067, n47068, n47069, n47070, n47071, n47072, n47073, n47074, n47075,
    n47076, n47077, n47078, n47079, n47080, n47081, n47082, n47083, n47084,
    n47085, n47086, n47087, n47088, n47089, n47090, n47091, n47092, n47093,
    n47094, n47095, n47096, n47097, n47098, n47099, n47100, n47101, n47102,
    n47103, n47104, n47105, n47106, n47107, n47108, n47109, n47110, n47111,
    n47112, n47113, n47114, n47115, n47116, n47117, n47118, n47119, n47120,
    n47121, n47122, n47123, n47124, n47125, n47126, n47127, n47128, n47129,
    n47130, n47131, n47132, n47133, n47134, n47135, n47136, n47137, n47138,
    n47139, n47140, n47141, n47142, n47143, n47144, n47145, n47146, n47147,
    n47148, n47149, n47150, n47151, n47152, n47153, n47154, n47155, n47156,
    n47157, n47158, n47159, n47160, n47161, n47162, n47163, n47164, n47165,
    n47166, n47167, n47168, n47169, n47170, n47171, n47172, n47173, n47174,
    n47175, n47176, n47177, n47178, n47179, n47180, n47181, n47182, n47183,
    n47184, n47185, n47186, n47187, n47188, n47189, n47190, n47191, n47192,
    n47193, n47194, n47195, n47196, n47197, n47198, n47199, n47200, n47201,
    n47202, n47203, n47204, n47205, n47206, n47207, n47208, n47209, n47210,
    n47211, n47212, n47213, n47214, n47215, n47216, n47217, n47218, n47219,
    n47220, n47221, n47222, n47223, n47224, n47225, n47226, n47227, n47228,
    n47229, n47230, n47231, n47232, n47233, n47234, n47235, n47236, n47237,
    n47238, n47239, n47240, n47241, n47242, n47243, n47244, n47245, n47246,
    n47247, n47248, n47249, n47250, n47251, n47252, n47253, n47254, n47255,
    n47256, n47257, n47258, n47259, n47260, n47261, n47262, n47263, n47264,
    n47265, n47266, n47267, n47268, n47269, n47270, n47271, n47272, n47273,
    n47274, n47275, n47276, n47277, n47278, n47279, n47280, n47281, n47282,
    n47283, n47284, n47285, n47286, n47287, n47288, n47289, n47290, n47291,
    n47292, n47293, n47294, n47295, n47296, n47297, n47298, n47299, n47300,
    n47301, n47302, n47303, n47304, n47305, n47306, n47307, n47308, n47309,
    n47310, n47311, n47312, n47313, n47314, n47315, n47316, n47317, n47318,
    n47319, n47320, n47321, n47322, n47323, n47324, n47325, n47326, n47327,
    n47328, n47329, n47330, n47331, n47332, n47333, n47334, n47335, n47336,
    n47337, n47338, n47339, n47340, n47341, n47342, n47343, n47344, n47345,
    n47346, n47347, n47348, n47349, n47350, n47351, n47352, n47353, n47354,
    n47355, n47356, n47357, n47358, n47359, n47360, n47361, n47362, n47363,
    n47364, n47365, n47366, n47367, n47368, n47369, n47370, n47371, n47372,
    n47373, n47374, n47375, n47376, n47377, n47378, n47379, n47380, n47381,
    n47382, n47383, n47384, n47385, n47386, n47387, n47388, n47389, n47390,
    n47391, n47392, n47393, n47394, n47395, n47396, n47397, n47398, n47399,
    n47400, n47401, n47402, n47403, n47404, n47405, n47406, n47407, n47408,
    n47409, n47410, n47411, n47412, n47413, n47414, n47415, n47416, n47417,
    n47418, n47419, n47420, n47421, n47422, n47423, n47424, n47425, n47426,
    n47427, n47428, n47429, n47430, n47431, n47432, n47433, n47434, n47435,
    n47436, n47437, n47438, n47439, n47440, n47441, n47442, n47443, n47444,
    n47445, n47446, n47447, n47448, n47449, n47450, n47451, n47452, n47453,
    n47454, n47455, n47456, n47457, n47458, n47459, n47460, n47461, n47462,
    n47463, n47464, n47465, n47466, n47467, n47468, n47469, n47470, n47471,
    n47472, n47473, n47474, n47475, n47476, n47477, n47478, n47479, n47480,
    n47481, n47482, n47483, n47484, n47485, n47486, n47487, n47488, n47489,
    n47490, n47491, n47492, n47493, n47494, n47495, n47496, n47497, n47498,
    n47499, n47500, n47501, n47502, n47503, n47504, n47505, n47506, n47507,
    n47508, n47509, n47510, n47511, n47512, n47513, n47514, n47515, n47516,
    n47517, n47518, n47519, n47520, n47521, n47522, n47523, n47524, n47525,
    n47526, n47527, n47528, n47529, n47530, n47531, n47532, n47533, n47534,
    n47535, n47536, n47537, n47538, n47539, n47540, n47541, n47542, n47543,
    n47544, n47545, n47546, n47547, n47548, n47549, n47550, n47551, n47552,
    n47553, n47554, n47555, n47556, n47557, n47558, n47559, n47560, n47561,
    n47562, n47563, n47564, n47565, n47566, n47567, n47568, n47569, n47570,
    n47571, n47572, n47573, n47574, n47575, n47576, n47577, n47578, n47579,
    n47580, n47581, n47582, n47583, n47584, n47585, n47586, n47587, n47588,
    n47589, n47590, n47591, n47592, n47593, n47594, n47595, n47596, n47597,
    n47598, n47599, n47600, n47601, n47602, n47603, n47604, n47605, n47606,
    n47607, n47608, n47609, n47610, n47611, n47612, n47613, n47614, n47615,
    n47616, n47617, n47618, n47619, n47620, n47621, n47622, n47623, n47624,
    n47625, n47626, n47627, n47628, n47629, n47630, n47631, n47632, n47633,
    n47634, n47635, n47636, n47637, n47638, n47639, n47640, n47641, n47642,
    n47643, n47644, n47645, n47646, n47647, n47648, n47649, n47650, n47651,
    n47652, n47653, n47654, n47655, n47656, n47657, n47658, n47659, n47660,
    n47661, n47662, n47663, n47664, n47665, n47666, n47667, n47668, n47669,
    n47670, n47671, n47672, n47673, n47674, n47675, n47676, n47677, n47678,
    n47679, n47680, n47681, n47682, n47683, n47684, n47685, n47686, n47687,
    n47688, n47689, n47690, n47691, n47692, n47693, n47694, n47695, n47696,
    n47697, n47698, n47699, n47700, n47701, n47702, n47703, n47704, n47705,
    n47706, n47707, n47708, n47709, n47710, n47711, n47712, n47713, n47714,
    n47715, n47716, n47717, n47718, n47719, n47720, n47721, n47722, n47723,
    n47724, n47725, n47726, n47727, n47728, n47729, n47730, n47731, n47732,
    n47733, n47734, n47735, n47736, n47737, n47738, n47739, n47740, n47741,
    n47742, n47743, n47744, n47745, n47746, n47747, n47748, n47749, n47750,
    n47751, n47752, n47753, n47754, n47755, n47756, n47757, n47758, n47759,
    n47760, n47761, n47762, n47763, n47764, n47765, n47766, n47767, n47768,
    n47769, n47770, n47771, n47772, n47773, n47774, n47775, n47776, n47777,
    n47778, n47779, n47780, n47781, n47782, n47783, n47784, n47785, n47786,
    n47787, n47788, n47789, n47790, n47791, n47792, n47793, n47794, n47795,
    n47796, n47797, n47798, n47799, n47800, n47801, n47802, n47803, n47804,
    n47805, n47806, n47807, n47808, n47809, n47810, n47811, n47812, n47813,
    n47814, n47815, n47816, n47817, n47818, n47819, n47820, n47821, n47822,
    n47823, n47824, n47825, n47826, n47827, n47828, n47829, n47830, n47831,
    n47832, n47833, n47834, n47835, n47836, n47837, n47838, n47839, n47840,
    n47841, n47842, n47843, n47844, n47845, n47846, n47847, n47848, n47849,
    n47850, n47851, n47852, n47853, n47854, n47855, n47856, n47857, n47858,
    n47859, n47860, n47861, n47862, n47863, n47864, n47865, n47866, n47867,
    n47868, n47869, n47870, n47871, n47872, n47873, n47874, n47875, n47876,
    n47877, n47878, n47879, n47880, n47881, n47882, n47883, n47884, n47885,
    n47886, n47887, n47888, n47889, n47890, n47891, n47892, n47893, n47894,
    n47895, n47896, n47897, n47898, n47899, n47900, n47901, n47902, n47903,
    n47904, n47905, n47906, n47907, n47908, n47909, n47910, n47911, n47912,
    n47913, n47914, n47915, n47916, n47917, n47918, n47919, n47920, n47921,
    n47922, n47923, n47924, n47925, n47926, n47927, n47928, n47929, n47930,
    n47931, n47932, n47933, n47934, n47935, n47936, n47937, n47938, n47939,
    n47940, n47941, n47942, n47943, n47944, n47945, n47946, n47947, n47948,
    n47949, n47950, n47951, n47952, n47953, n47954, n47955, n47956, n47957,
    n47958, n47959, n47960, n47961, n47962, n47963, n47964, n47965, n47966,
    n47967, n47968, n47969, n47970, n47971, n47972, n47973, n47974, n47975,
    n47976, n47977, n47978, n47979, n47980, n47981, n47982, n47983, n47984,
    n47985, n47986, n47987, n47988, n47989, n47990, n47991, n47992, n47993,
    n47994, n47995, n47996, n47997, n47998, n47999, n48000, n48001, n48002,
    n48003, n48004, n48005, n48006, n48007, n48008, n48009, n48010, n48011,
    n48012, n48013, n48014, n48015, n48016, n48017, n48018, n48019, n48020,
    n48021, n48022, n48023, n48024, n48025, n48026, n48027, n48028, n48029,
    n48030, n48031, n48032, n48033, n48034, n48035, n48036, n48037, n48038,
    n48039, n48040, n48041, n48042, n48043, n48044, n48045, n48046, n48047,
    n48048, n48049, n48050, n48051, n48052, n48053, n48054, n48055, n48056,
    n48057, n48058, n48059, n48060, n48061, n48062, n48063, n48064, n48065,
    n48066, n48067, n48068, n48069, n48070, n48071, n48072, n48073, n48074,
    n48075, n48076, n48077, n48078, n48079, n48080, n48081, n48082, n48083,
    n48084, n48085, n48086, n48087, n48088, n48089, n48090, n48091, n48092,
    n48093, n48094, n48095, n48096, n48097, n48098, n48099, n48100, n48101,
    n48102, n48103, n48104, n48105, n48106, n48107, n48108, n48109, n48110,
    n48111, n48112, n48113, n48114, n48115, n48116, n48117, n48118, n48119,
    n48120, n48121, n48122, n48123, n48124, n48125, n48126, n48127, n48128,
    n48129, n48130, n48131, n48132, n48133, n48134, n48135, n48136, n48137,
    n48138, n48139, n48140, n48141, n48142, n48143, n48144, n48145, n48146,
    n48147, n48148, n48149, n48150, n48151, n48152, n48153, n48154, n48155,
    n48156, n48157, n48158, n48159, n48160, n48161, n48162, n48163, n48164,
    n48165, n48166, n48167, n48168, n48169, n48170, n48171, n48172, n48173,
    n48174, n48175, n48176, n48177, n48178, n48179, n48180, n48181, n48182,
    n48183, n48184, n48185, n48186, n48187, n48188, n48189, n48190, n48191,
    n48192, n48193, n48194, n48195, n48196, n48197, n48198, n48199, n48200,
    n48201, n48202, n48203, n48204, n48205, n48206, n48207, n48208, n48209,
    n48210, n48211, n48212, n48213, n48214, n48215, n48216, n48217, n48218,
    n48219, n48220, n48221, n48222, n48223, n48224, n48225, n48226, n48227,
    n48228, n48229, n48230, n48231, n48232, n48233, n48234, n48235, n48236,
    n48237, n48238, n48239, n48240, n48241, n48242, n48243, n48244, n48245,
    n48246, n48247, n48248, n48249, n48250, n48251, n48252, n48253, n48254,
    n48255, n48256, n48257, n48258, n48259, n48260, n48261, n48262, n48263,
    n48264, n48265, n48266, n48267, n48268, n48269, n48270, n48271, n48272,
    n48273, n48274, n48275, n48276, n48277, n48278, n48279, n48280, n48281,
    n48282, n48283, n48284, n48285, n48286, n48287, n48288, n48289, n48290,
    n48291, n48292, n48293, n48294, n48295, n48296, n48297, n48298, n48299,
    n48300, n48301, n48302, n48303, n48304, n48305, n48306, n48307, n48308,
    n48309, n48310, n48311, n48312, n48313, n48314, n48315, n48316, n48317,
    n48318, n48319, n48320, n48321, n48322, n48323, n48324, n48325, n48326,
    n48327, n48328, n48329, n48330, n48331, n48332, n48333, n48334, n48335,
    n48336, n48337, n48338, n48339, n48340, n48341, n48342, n48343, n48344,
    n48345, n48346, n48347, n48348, n48349, n48350, n48351, n48352, n48353,
    n48354, n48355, n48356, n48357, n48358, n48359, n48360, n48361, n48362,
    n48363, n48364, n48365, n48366, n48367, n48368, n48369, n48370, n48371,
    n48372, n48373, n48374, n48375, n48376, n48377, n48378, n48379, n48380,
    n48381, n48382, n48383, n48384, n48385, n48386, n48387, n48388, n48389,
    n48390, n48391, n48392, n48393, n48394, n48395, n48396, n48397, n48398,
    n48399, n48400, n48401, n48402, n48403, n48404, n48405, n48406, n48407,
    n48408, n48409, n48410, n48411, n48412, n48413, n48414, n48415, n48416,
    n48417, n48418, n48419, n48420, n48421, n48422, n48423, n48424, n48425,
    n48426, n48427, n48428, n48429, n48430, n48431, n48432, n48433, n48434,
    n48435, n48436, n48437, n48438, n48439, n48440, n48441, n48442, n48443,
    n48444, n48445, n48446, n48447, n48448, n48449, n48450, n48451, n48452,
    n48453, n48454, n48455, n48456, n48457, n48458, n48459, n48460, n48461,
    n48462, n48463, n48464, n48465, n48466, n48467, n48468, n48469, n48470,
    n48471, n48472, n48473, n48474, n48475, n48476, n48477, n48478, n48479,
    n48480, n48481, n48482, n48483, n48484, n48485, n48486, n48487, n48488,
    n48489, n48490, n48491, n48492, n48493, n48494, n48495, n48496, n48497,
    n48498, n48499, n48500, n48501, n48502, n48503, n48504, n48505, n48506,
    n48507, n48508, n48509, n48510, n48511, n48512, n48513, n48514, n48515,
    n48516, n48517, n48518, n48519, n48520, n48521, n48522, n48523, n48524,
    n48525, n48526, n48527, n48528, n48529, n48530, n48531, n48532, n48533,
    n48534, n48535, n48536, n48537, n48538, n48539, n48540, n48541, n48542,
    n48543, n48544, n48545, n48546, n48547, n48548, n48549, n48550, n48551,
    n48552, n48553, n48554, n48555, n48556, n48557, n48558, n48559, n48560,
    n48561, n48562, n48563, n48564, n48565, n48566, n48567, n48568, n48569,
    n48570, n48571, n48572, n48573, n48574, n48575, n48576, n48577, n48578,
    n48579, n48580, n48581, n48582, n48583, n48584, n48585, n48586, n48587,
    n48588, n48589, n48590, n48591, n48592, n48593, n48594, n48595, n48596,
    n48597, n48598, n48599, n48600, n48601, n48602, n48603, n48604, n48605,
    n48606, n48607, n48608, n48609, n48610, n48611, n48612, n48613, n48614,
    n48615, n48616, n48617, n48618, n48619, n48620, n48621, n48622, n48623,
    n48624, n48625, n48626, n48627, n48628, n48629, n48630, n48631, n48632,
    n48633, n48634, n48635, n48636, n48637, n48638, n48639, n48640, n48641,
    n48642, n48643, n48644, n48645, n48646, n48647, n48648, n48649, n48650,
    n48651, n48652, n48653, n48654, n48655, n48656, n48657, n48658, n48659,
    n48660, n48661, n48662, n48663, n48664, n48665, n48666, n48667, n48668,
    n48669, n48670, n48671, n48672, n48673, n48674, n48675, n48676, n48677,
    n48678, n48679, n48680, n48681, n48682, n48683, n48684, n48685, n48686,
    n48687, n48688, n48689, n48690, n48691, n48692, n48693, n48694, n48695,
    n48696, n48697, n48698, n48699, n48700, n48701, n48702, n48703, n48704,
    n48705, n48706, n48707, n48708, n48709, n48710, n48711, n48712, n48713,
    n48714, n48715, n48716, n48717, n48718, n48719, n48720, n48721, n48722,
    n48723, n48724, n48725, n48726, n48727, n48728, n48729, n48730, n48731,
    n48732, n48733, n48734, n48735, n48736, n48737, n48738, n48739, n48740,
    n48741, n48742, n48743, n48744, n48745, n48746, n48747, n48748, n48749,
    n48750, n48751, n48752, n48753, n48754, n48755, n48756, n48757, n48758,
    n48759, n48760, n48761, n48762, n48763, n48764, n48765, n48766, n48767,
    n48768, n48769, n48770, n48771, n48772, n48773, n48774, n48775, n48776,
    n48777, n48778, n48779, n48780, n48781, n48782, n48783, n48784, n48785,
    n48786, n48787, n48788, n48789, n48790, n48791, n48792, n48793, n48794,
    n48795, n48796, n48797, n48798, n48799, n48800, n48801, n48802, n48803,
    n48804, n48805, n48806, n48807, n48808, n48809, n48810, n48811, n48812,
    n48813, n48814, n48815, n48816, n48817, n48818, n48819, n48820, n48821,
    n48822, n48823, n48824, n48825, n48826, n48827, n48828, n48829, n48830,
    n48831, n48832, n48833, n48834, n48835, n48836, n48837, n48838, n48839,
    n48840, n48841, n48842, n48843, n48844, n48845, n48846, n48847, n48848,
    n48849, n48850, n48851, n48852, n48853, n48854, n48855, n48856, n48857,
    n48858, n48859, n48860, n48861, n48862, n48863, n48864, n48865, n48866,
    n48867, n48868, n48869, n48870, n48871, n48872, n48873, n48874, n48875,
    n48876, n48877, n48878, n48879, n48880, n48881, n48882, n48883, n48884,
    n48885, n48886, n48887, n48888, n48889, n48890, n48891, n48892, n48893,
    n48894, n48895, n48896, n48897, n48898, n48899, n48900, n48901, n48902,
    n48903, n48904, n48905, n48906, n48907, n48908, n48909, n48910, n48911,
    n48912, n48913, n48914, n48915, n48916, n48917, n48918, n48919, n48920,
    n48921, n48922, n48923, n48924, n48925, n48926, n48927, n48928, n48929,
    n48930, n48931, n48932, n48933, n48934, n48935, n48936, n48937, n48938,
    n48939, n48940, n48941, n48942, n48943, n48944, n48945, n48946, n48947,
    n48948, n48949, n48950, n48951, n48952, n48953, n48954, n48955, n48956,
    n48957, n48958, n48959, n48960, n48961, n48962, n48963, n48964, n48965,
    n48966, n48967, n48968, n48969, n48970, n48971, n48972, n48973, n48974,
    n48975, n48976, n48977, n48978, n48979, n48980, n48981, n48982, n48983,
    n48984, n48985, n48986, n48987, n48988, n48989, n48990, n48991, n48992,
    n48993, n48994, n48995, n48996, n48997, n48998, n48999, n49000, n49001,
    n49002, n49003, n49004, n49005, n49006, n49007, n49008, n49009, n49010,
    n49011, n49012, n49013, n49014, n49015, n49016, n49017, n49018, n49019,
    n49020, n49021, n49022, n49023, n49024, n49025, n49026, n49027, n49028,
    n49029, n49030, n49031, n49032, n49033, n49034, n49035, n49036, n49037,
    n49038, n49039, n49040, n49041, n49042, n49043, n49044, n49045, n49046,
    n49047, n49048, n49049, n49050, n49051, n49052, n49053, n49054, n49055,
    n49056, n49057, n49058, n49059, n49060, n49061, n49062, n49063, n49064,
    n49065, n49066, n49067, n49068, n49069, n49070, n49071, n49072, n49073,
    n49074, n49075, n49076, n49077, n49078, n49079, n49080, n49081, n49082,
    n49083, n49084, n49085, n49086, n49087, n49088, n49089, n49090, n49091,
    n49092, n49093, n49094, n49095, n49096, n49097, n49098, n49099, n49100,
    n49101, n49102, n49103, n49104, n49105, n49106, n49107, n49108, n49109,
    n49110, n49111, n49112, n49113, n49114, n49115, n49116, n49117, n49118,
    n49119, n49120, n49121, n49122, n49123, n49124, n49125, n49126, n49127,
    n49128, n49129, n49130, n49131, n49132, n49133, n49134, n49135, n49136,
    n49137, n49138, n49139, n49140, n49141, n49142, n49143, n49144, n49145,
    n49146, n49147, n49148, n49149, n49150, n49151, n49152, n49153, n49154,
    n49155, n49156, n49157, n49158, n49159, n49160, n49161, n49162, n49163,
    n49164, n49165, n49166, n49167, n49168, n49169, n49170, n49171, n49172,
    n49173, n49174, n49175, n49176, n49177, n49178, n49179, n49180, n49181,
    n49182, n49183, n49184, n49185, n49186, n49187, n49188, n49189, n49190,
    n49191, n49192, n49193, n49194, n49195, n49196, n49197, n49198, n49199,
    n49200, n49201, n49202, n49203, n49204, n49205, n49206, n49207, n49208,
    n49209, n49210, n49211, n49212, n49213, n49214, n49215, n49216, n49217,
    n49218, n49219, n49220, n49221, n49222, n49223, n49224, n49225, n49226,
    n49227, n49228, n49229, n49230, n49231, n49232, n49233, n49234, n49235,
    n49236, n49237, n49238, n49239, n49240, n49241, n49242, n49243, n49244,
    n49245, n49246, n49247, n49248, n49249, n49250, n49251, n49252, n49253,
    n49254, n49255, n49256, n49257, n49258, n49259, n49260, n49261, n49262,
    n49263, n49264, n49265, n49266, n49267, n49268, n49269, n49270, n49271,
    n49272, n49273, n49274, n49275, n49276, n49277, n49278, n49279, n49280,
    n49281, n49282, n49283, n49284, n49285, n49286, n49287, n49288, n49289,
    n49290, n49291, n49292, n49293, n49294, n49295, n49296, n49297, n49298,
    n49299, n49300, n49301, n49302, n49303, n49304, n49305, n49306, n49307,
    n49308, n49309, n49310, n49311, n49312, n49313, n49314, n49315, n49316,
    n49317, n49318, n49319, n49320, n49321, n49322, n49323, n49324, n49325,
    n49326, n49327, n49328, n49329, n49330, n49331, n49332, n49333, n49334,
    n49335, n49336, n49337, n49338, n49339, n49340, n49341, n49342, n49343,
    n49344, n49345, n49346, n49347, n49348, n49349, n49350, n49351, n49352,
    n49353, n49354, n49355, n49356, n49357, n49358, n49359, n49360, n49361,
    n49362, n49363, n49364, n49365, n49366, n49367, n49368, n49369, n49370,
    n49371, n49372, n49373, n49374, n49375, n49376, n49377, n49378, n49379,
    n49380, n49381, n49382, n49383, n49384, n49385, n49386, n49387, n49388,
    n49389, n49390, n49391, n49392, n49393, n49394, n49395, n49396, n49397,
    n49398, n49399, n49400, n49401, n49402, n49403, n49404, n49405, n49406,
    n49407, n49408, n49409, n49410, n49411, n49412, n49413, n49414, n49415,
    n49416, n49417, n49418, n49419, n49420, n49421, n49422, n49423, n49424,
    n49425, n49426, n49427, n49428, n49429, n49430, n49431, n49432, n49433,
    n49434, n49435, n49436, n49437, n49438, n49439, n49440, n49441, n49442,
    n49443, n49444, n49445, n49446, n49447, n49448, n49449, n49450, n49451,
    n49452, n49453, n49454, n49455, n49456, n49457, n49458, n49459, n49460,
    n49461, n49462, n49463, n49464, n49465, n49466, n49467, n49468, n49469,
    n49470, n49471, n49472, n49473, n49474, n49475, n49476, n49477, n49478,
    n49479, n49480, n49481, n49482, n49483, n49484, n49485, n49486, n49487,
    n49488, n49489, n49490, n49491, n49492, n49493, n49494, n49495, n49496,
    n49497, n49498, n49499, n49500, n49501, n49502, n49503, n49504, n49505,
    n49506, n49507, n49508, n49509, n49510, n49511, n49512, n49513, n49514,
    n49515, n49516, n49517, n49518, n49519, n49520, n49521, n49522, n49523,
    n49524, n49525, n49526, n49527, n49528, n49529, n49530, n49531, n49532,
    n49533, n49534, n49535, n49536, n49537, n49538, n49539, n49540, n49541,
    n49542, n49543, n49544, n49545, n49546, n49547, n49548, n49549, n49550,
    n49551, n49552, n49553, n49554, n49555, n49556, n49557, n49558, n49559,
    n49560, n49561, n49562, n49563, n49564, n49565, n49566, n49567, n49568,
    n49569, n49570, n49571, n49572, n49573, n49574, n49575, n49576, n49577,
    n49578, n49579, n49580, n49581, n49582, n49583, n49584, n49585, n49586,
    n49587, n49588, n49589, n49590, n49591, n49592, n49593, n49594, n49595,
    n49596, n49597, n49598, n49599, n49600, n49601, n49602, n49603, n49604,
    n49605, n49606, n49607, n49608, n49609, n49610, n49611, n49612, n49613,
    n49614, n49615, n49616, n49617, n49618, n49619, n49620, n49621, n49622,
    n49623, n49624, n49625, n49626, n49627, n49628, n49629, n49630, n49631,
    n49632, n49633, n49634, n49635, n49636, n49637, n49638, n49639, n49640,
    n49641, n49642, n49643, n49644, n49645, n49646, n49647, n49648, n49649,
    n49650, n49651, n49652, n49653, n49654, n49655, n49656, n49657, n49658,
    n49659, n49660, n49661, n49662, n49663, n49664, n49665, n49666, n49667,
    n49668, n49669, n49670, n49671, n49672, n49673, n49674, n49675, n49676,
    n49677, n49678, n49679, n49680, n49681, n49682, n49683, n49684, n49685,
    n49686, n49687, n49688, n49689, n49690, n49691, n49692, n49693, n49694,
    n49695, n49696, n49697, n49698, n49699, n49700, n49701, n49702, n49703,
    n49704, n49705, n49706, n49707, n49708, n49709, n49710, n49711, n49712,
    n49713, n49714, n49715, n49716, n49717, n49718, n49719, n49720, n49721,
    n49722, n49723, n49724, n49725, n49726, n49727, n49728, n49729, n49730,
    n49731, n49732, n49733, n49734, n49735, n49736, n49737, n49738, n49739,
    n49740, n49741, n49742, n49743, n49744, n49745, n49746, n49747, n49748,
    n49749, n49750, n49751, n49752, n49753, n49754, n49755, n49756, n49757,
    n49758, n49759, n49760, n49761, n49762, n49763, n49764, n49765, n49766,
    n49767, n49768, n49769, n49770, n49771, n49772, n49773, n49774, n49775,
    n49776, n49777, n49778, n49779, n49780, n49781, n49782, n49783, n49784,
    n49785, n49786, n49787, n49788, n49789, n49790, n49791, n49792, n49793,
    n49794, n49795, n49796, n49797, n49798, n49799, n49800, n49801, n49802,
    n49803, n49804, n49805, n49806, n49807, n49808, n49809, n49810, n49811,
    n49812, n49813, n49814, n49815, n49816, n49817, n49818, n49819, n49820,
    n49821, n49822, n49823, n49824, n49825, n49826, n49827, n49828, n49829,
    n49830, n49831, n49832, n49833, n49834, n49835, n49836, n49837, n49838,
    n49839, n49840, n49841, n49842, n49843, n49844, n49845, n49846, n49847,
    n49848, n49849, n49850, n49851, n49852, n49853, n49854, n49855, n49856,
    n49857, n49858, n49859, n49860, n49861, n49862, n49863, n49864, n49865,
    n49866, n49867, n49868, n49869, n49870, n49871, n49872, n49873, n49874,
    n49875, n49876, n49877, n49878, n49879, n49880, n49881, n49882, n49883,
    n49884, n49885, n49886, n49887, n49888, n49889, n49890, n49891, n49892,
    n49893, n49894, n49895, n49896, n49897, n49898, n49899, n49900, n49901,
    n49902, n49903, n49904, n49905, n49906, n49907, n49908, n49909, n49910,
    n49911, n49912, n49913, n49914, n49915, n49916, n49917, n49918, n49919,
    n49920, n49921, n49922, n49923, n49924, n49925, n49926, n49927, n49928,
    n49929, n49930, n49931, n49932, n49933, n49934, n49935, n49936, n49937,
    n49938, n49939, n49940, n49941, n49942, n49943, n49944, n49945, n49946,
    n49947, n49948, n49949, n49950, n49951, n49952, n49953, n49954, n49955,
    n49956, n49957, n49958, n49959, n49960, n49961, n49962, n49963, n49964,
    n49965, n49966, n49967, n49968, n49969, n49970, n49971, n49972, n49973,
    n49974, n49975, n49976, n49977, n49978, n49979, n49980, n49981, n49982,
    n49983, n49984, n49985, n49986, n49987, n49988, n49989, n49990, n49991,
    n49992, n49993, n49994, n49995, n49996, n49997, n49998, n49999, n50000,
    n50001, n50002, n50003, n50004, n50005, n50006, n50007, n50008, n50009,
    n50010, n50011, n50012, n50013, n50014, n50015, n50016, n50017, n50018,
    n50019, n50020, n50021, n50022, n50023, n50024, n50025, n50026, n50027,
    n50028, n50029, n50030, n50031, n50032, n50033, n50034, n50035, n50036,
    n50037, n50038, n50039, n50040, n50041, n50042, n50043, n50044, n50045,
    n50046, n50047, n50048, n50049, n50050, n50051, n50052, n50053, n50054,
    n50055, n50056, n50057, n50058, n50059, n50060, n50061, n50062, n50063,
    n50064, n50065, n50066, n50067, n50068, n50069, n50070, n50071, n50072,
    n50073, n50074, n50075, n50076, n50077, n50078, n50079, n50080, n50081,
    n50082, n50083, n50084, n50085, n50086, n50087, n50088, n50089, n50090,
    n50091, n50092, n50093, n50094, n50095, n50096, n50097, n50098, n50099,
    n50100, n50101, n50102, n50103, n50104, n50105, n50106, n50107, n50108,
    n50109, n50110, n50111, n50112, n50113, n50114, n50115, n50116, n50117,
    n50118, n50119, n50120, n50121, n50122, n50123, n50124, n50125, n50126,
    n50127, n50128, n50129, n50130, n50131, n50132, n50133, n50134, n50135,
    n50136, n50137, n50138, n50139, n50140, n50141, n50142, n50143, n50144,
    n50145, n50146, n50147, n50148, n50149, n50150, n50151, n50152, n50153,
    n50154, n50155, n50156, n50157, n50158, n50159, n50160, n50161, n50162,
    n50163, n50164, n50165, n50166, n50167, n50168, n50169, n50170, n50171,
    n50172, n50173, n50174, n50175, n50176, n50177, n50178, n50179, n50180,
    n50181, n50182, n50183, n50184, n50185, n50186, n50187, n50188, n50189,
    n50191, n50192, n50193, n50194, n50195, n50196, n50197, n50198, n50199,
    n50200, n50201, n50202, n50203, n50204, n50205, n50206, n50207, n50208,
    n50209, n50210, n50211, n50212, n50213, n50214, n50215, n50216, n50217,
    n50218, n50219, n50220, n50221, n50222, n50223, n50224, n50225, n50226,
    n50227, n50228, n50229, n50230, n50231, n50232, n50233, n50234, n50235,
    n50236, n50237, n50238, n50240, n50241, n50242, n50243, n50244, n50245,
    n50246, n50247, n50248, n50249, n50250, n50251, n50252, n50253, n50254,
    n50255, n50256, n50257, n50258, n50259, n50260, n50261, n50262, n50263,
    n50264, n50265, n50266, n50267, n50268, n50269, n50270, n50271, n50272,
    n50273, n50274, n50275, n50276, n50277, n50278, n50279, n50280, n50282,
    n50283, n50284, n50285, n50286, n50287, n50288, n50289, n50290, n50291,
    n50292, n50293, n50294, n50295, n50296, n50297, n50298, n50299, n50300,
    n50301, n50302, n50303, n50304, n50305, n50306, n50307, n50308, n50309,
    n50310, n50311, n50312, n50313, n50314, n50315, n50316, n50317, n50318,
    n50319, n50320, n50321, n50322, n50323, n50324, n50325, n50326, n50328,
    n50329, n50330, n50331, n50332, n50333, n50334, n50335, n50336, n50337,
    n50338, n50339, n50340, n50341, n50342, n50343, n50344, n50345, n50346,
    n50347, n50348, n50349, n50350, n50351, n50352, n50353, n50354, n50355,
    n50356, n50357, n50358, n50359, n50360, n50361, n50362, n50363, n50364,
    n50365, n50366, n50367, n50369, n50370, n50371, n50372, n50373, n50374,
    n50375, n50376, n50377, n50378, n50379, n50380, n50381, n50382, n50383,
    n50384, n50385, n50386, n50387, n50388, n50389, n50390, n50391, n50392,
    n50393, n50394, n50395, n50396, n50397, n50398, n50399, n50400, n50401,
    n50402, n50403, n50404, n50405, n50406, n50407, n50408, n50409, n50410,
    n50411, n50412, n50413, n50414, n50415, n50417, n50418, n50419, n50420,
    n50421, n50422, n50423, n50424, n50425, n50426, n50427, n50428, n50429,
    n50430, n50431, n50432, n50433, n50434, n50435, n50436, n50437, n50438,
    n50439, n50440, n50441, n50442, n50443, n50444, n50445, n50446, n50447,
    n50448, n50449, n50450, n50451, n50452, n50453, n50455, n50456, n50457,
    n50458, n50459, n50460, n50461, n50462, n50463, n50464, n50465, n50466,
    n50467, n50468, n50469, n50470, n50471, n50472, n50473, n50474, n50475,
    n50476, n50477, n50478, n50479, n50480, n50481, n50482, n50483, n50484,
    n50485, n50486, n50487, n50488, n50489, n50490, n50491, n50492, n50494,
    n50495, n50496, n50497, n50498, n50499, n50500, n50501, n50502, n50503,
    n50504, n50505, n50506, n50507, n50508, n50509, n50510, n50511, n50512,
    n50513, n50514, n50515, n50516, n50517, n50518, n50519, n50521, n50522,
    n50523, n50524, n50525, n50526, n50527, n50528, n50530, n50531, n50532,
    n50533, n50534, n50535, n50536, n50537, n50539, n50540, n50541, n50542,
    n50543, n50544, n50545, n50546, n50548, n50549, n50550, n50551, n50552,
    n50553, n50554, n50555, n50557, n50558, n50559, n50560, n50561, n50562,
    n50563, n50564, n50566, n50567, n50568, n50569, n50570, n50571, n50572,
    n50573, n50575, n50576, n50577, n50578, n50579, n50580, n50581, n50582,
    n50584, n50585, n50586, n50587, n50588, n50589, n50590, n50591, n50592,
    n50593, n50594, n50595, n50596, n50597, n50598, n50599, n50600, n50601,
    n50602, n50603, n50604, n50605, n50606, n50607, n50608, n50610, n50611,
    n50612, n50613, n50614, n50615, n50616, n50617, n50619, n50620, n50621,
    n50622, n50623, n50624, n50625, n50626, n50628, n50629, n50630, n50631,
    n50632, n50633, n50634, n50635, n50637, n50638, n50639, n50640, n50641,
    n50642, n50643, n50644, n50646, n50647, n50648, n50649, n50650, n50651,
    n50652, n50653, n50655, n50656, n50657, n50658, n50659, n50660, n50661,
    n50662, n50664, n50665, n50666, n50667, n50668, n50669, n50670, n50671,
    n50673, n50674, n50675, n50676, n50677, n50678, n50679, n50680, n50681,
    n50682, n50683, n50684, n50685, n50686, n50687, n50688, n50689, n50690,
    n50691, n50692, n50693, n50694, n50695, n50696, n50697, n50699, n50700,
    n50701, n50702, n50703, n50704, n50705, n50706, n50708, n50709, n50710,
    n50711, n50712, n50713, n50714, n50715, n50717, n50718, n50719, n50720,
    n50721, n50722, n50723, n50724, n50726, n50727, n50728, n50729, n50730,
    n50731, n50732, n50733, n50735, n50736, n50737, n50738, n50739, n50740,
    n50741, n50742, n50744, n50745, n50746, n50747, n50748, n50749, n50750,
    n50751, n50753, n50754, n50755, n50756, n50757, n50758, n50759, n50760,
    n50762, n50763, n50764, n50765, n50766, n50767, n50768, n50769, n50770,
    n50771, n50772, n50773, n50774, n50775, n50776, n50777, n50778, n50779,
    n50780, n50781, n50782, n50783, n50784, n50785, n50786, n50787, n50789,
    n50790, n50791, n50792, n50793, n50794, n50795, n50796, n50798, n50799,
    n50800, n50801, n50802, n50803, n50804, n50805, n50807, n50808, n50809,
    n50810, n50811, n50812, n50813, n50814, n50816, n50817, n50818, n50819,
    n50820, n50821, n50822, n50823, n50825, n50826, n50827, n50828, n50829,
    n50830, n50831, n50832, n50834, n50835, n50836, n50837, n50838, n50839,
    n50840, n50841, n50843, n50844, n50845, n50846, n50847, n50848, n50849,
    n50850, n50852, n50853, n50854, n50855, n50856, n50857, n50858, n50859,
    n50860, n50861, n50862, n50863, n50864, n50865, n50866, n50867, n50868,
    n50869, n50870, n50871, n50872, n50873, n50874, n50875, n50877, n50878,
    n50879, n50880, n50881, n50882, n50883, n50884, n50886, n50887, n50888,
    n50889, n50890, n50891, n50892, n50893, n50895, n50896, n50897, n50898,
    n50899, n50900, n50901, n50902, n50904, n50905, n50906, n50907, n50908,
    n50909, n50910, n50911, n50913, n50914, n50915, n50916, n50917, n50918,
    n50919, n50920, n50922, n50923, n50924, n50925, n50926, n50927, n50928,
    n50929, n50931, n50932, n50933, n50934, n50935, n50936, n50937, n50938,
    n50940, n50941, n50942, n50943, n50944, n50945, n50946, n50947, n50948,
    n50949, n50950, n50951, n50952, n50953, n50954, n50955, n50956, n50957,
    n50958, n50959, n50960, n50961, n50962, n50964, n50965, n50966, n50967,
    n50968, n50969, n50970, n50971, n50973, n50974, n50975, n50976, n50977,
    n50978, n50979, n50980, n50982, n50983, n50984, n50985, n50986, n50987,
    n50988, n50989, n50991, n50992, n50993, n50994, n50995, n50996, n50997,
    n50998, n51000, n51001, n51002, n51003, n51004, n51005, n51006, n51007,
    n51009, n51010, n51011, n51012, n51013, n51014, n51015, n51016, n51018,
    n51019, n51020, n51021, n51022, n51023, n51024, n51025, n51027, n51028,
    n51029, n51030, n51031, n51032, n51033, n51034, n51035, n51036, n51037,
    n51038, n51039, n51040, n51041, n51042, n51043, n51044, n51045, n51046,
    n51047, n51048, n51050, n51051, n51052, n51053, n51054, n51055, n51056,
    n51057, n51059, n51060, n51061, n51062, n51063, n51064, n51065, n51066,
    n51068, n51069, n51070, n51071, n51072, n51073, n51074, n51075, n51077,
    n51078, n51079, n51080, n51081, n51082, n51083, n51084, n51086, n51087,
    n51088, n51089, n51090, n51091, n51092, n51093, n51095, n51096, n51097,
    n51098, n51099, n51100, n51101, n51102, n51104, n51105, n51106, n51107,
    n51108, n51109, n51110, n51111, n51113, n51114, n51115, n51116, n51117,
    n51118, n51119, n51120, n51121, n51122, n51123, n51124, n51125, n51126,
    n51127, n51128, n51129, n51130, n51131, n51132, n51133, n51135, n51136,
    n51137, n51138, n51139, n51140, n51141, n51142, n51144, n51145, n51146,
    n51147, n51148, n51149, n51150, n51151, n51153, n51154, n51155, n51156,
    n51157, n51158, n51159, n51160, n51162, n51163, n51164, n51165, n51166,
    n51167, n51168, n51169, n51171, n51172, n51173, n51174, n51175, n51176,
    n51177, n51178, n51180, n51181, n51182, n51183, n51184, n51185, n51186,
    n51187, n51189, n51190, n51191, n51192, n51193, n51194, n51195, n51196,
    n51198, n51199, n51200, n51201, n51202, n51203, n51204, n51205, n51206,
    n51207, n51208, n51209, n51210, n51211, n51212, n51213, n51214, n51215,
    n51216, n51217, n51218, n51219, n51220, n51221, n51223, n51224, n51225,
    n51226, n51227, n51228, n51229, n51230, n51232, n51233, n51234, n51235,
    n51236, n51237, n51238, n51239, n51241, n51242, n51243, n51244, n51245,
    n51246, n51247, n51248, n51250, n51251, n51252, n51253, n51254, n51255,
    n51256, n51257, n51259, n51260, n51261, n51262, n51263, n51264, n51265,
    n51266, n51268, n51269, n51270, n51271, n51272, n51273, n51274, n51275,
    n51277, n51278, n51279, n51280, n51281, n51282, n51283, n51284, n51286,
    n51287, n51288, n51289, n51290, n51291, n51292, n51293, n51294, n51295,
    n51296, n51297, n51298, n51299, n51300, n51301, n51302, n51303, n51304,
    n51305, n51306, n51307, n51308, n51309, n51311, n51312, n51313, n51314,
    n51315, n51316, n51317, n51318, n51320, n51321, n51322, n51323, n51324,
    n51325, n51326, n51327, n51329, n51330, n51331, n51332, n51333, n51334,
    n51335, n51336, n51338, n51339, n51340, n51341, n51342, n51343, n51344,
    n51345, n51347, n51348, n51349, n51350, n51351, n51352, n51353, n51354,
    n51356, n51357, n51358, n51359, n51360, n51361, n51362, n51363, n51365,
    n51366, n51367, n51368, n51369, n51370, n51371, n51372, n51374, n51375,
    n51376, n51377, n51378, n51379, n51380, n51381, n51382, n51383, n51384,
    n51385, n51386, n51387, n51388, n51389, n51390, n51391, n51392, n51393,
    n51394, n51395, n51397, n51398, n51399, n51400, n51401, n51402, n51403,
    n51404, n51406, n51407, n51408, n51409, n51410, n51411, n51412, n51413,
    n51415, n51416, n51417, n51418, n51419, n51420, n51421, n51422, n51424,
    n51425, n51426, n51427, n51428, n51429, n51430, n51431, n51433, n51434,
    n51435, n51436, n51437, n51438, n51439, n51440, n51442, n51443, n51444,
    n51445, n51446, n51447, n51448, n51449, n51451, n51452, n51453, n51454,
    n51455, n51456, n51457, n51458, n51460, n51461, n51462, n51463, n51464,
    n51465, n51466, n51467, n51468, n51469, n51470, n51471, n51472, n51473,
    n51474, n51475, n51476, n51477, n51478, n51479, n51480, n51481, n51482,
    n51483, n51484, n51486, n51487, n51488, n51489, n51490, n51491, n51492,
    n51493, n51495, n51496, n51497, n51498, n51499, n51500, n51501, n51502,
    n51504, n51505, n51506, n51507, n51508, n51509, n51510, n51511, n51513,
    n51514, n51515, n51516, n51517, n51518, n51519, n51520, n51522, n51523,
    n51524, n51525, n51526, n51527, n51528, n51529, n51531, n51532, n51533,
    n51534, n51535, n51536, n51537, n51538, n51540, n51541, n51542, n51543,
    n51544, n51545, n51546, n51547, n51549, n51550, n51551, n51552, n51553,
    n51554, n51555, n51556, n51557, n51558, n51559, n51560, n51561, n51562,
    n51563, n51564, n51565, n51566, n51567, n51568, n51569, n51571, n51572,
    n51573, n51574, n51575, n51576, n51577, n51578, n51580, n51581, n51582,
    n51583, n51584, n51585, n51586, n51587, n51589, n51590, n51591, n51592,
    n51593, n51594, n51595, n51596, n51598, n51599, n51600, n51601, n51602,
    n51603, n51604, n51605, n51607, n51608, n51609, n51610, n51611, n51612,
    n51613, n51614, n51616, n51617, n51618, n51619, n51620, n51621, n51622,
    n51623, n51625, n51626, n51627, n51628, n51629, n51630, n51631, n51632,
    n51634, n51635, n51636, n51637, n51638, n51639, n51640, n51641, n51642,
    n51643, n51644, n51645, n51646, n51647, n51648, n51649, n51650, n51651,
    n51652, n51653, n51654, n51656, n51657, n51658, n51659, n51660, n51661,
    n51662, n51663, n51665, n51666, n51667, n51668, n51669, n51670, n51671,
    n51672, n51674, n51675, n51676, n51677, n51678, n51679, n51680, n51681,
    n51683, n51684, n51685, n51686, n51687, n51688, n51689, n51690, n51692,
    n51693, n51694, n51695, n51696, n51697, n51698, n51699, n51701, n51702,
    n51703, n51704, n51705, n51706, n51707, n51708, n51710, n51711, n51712,
    n51713, n51714, n51715, n51716, n51717, n51719, n51720, n51721, n51722,
    n51723, n51724, n51725, n51726, n51727, n51728, n51729, n51730, n51731,
    n51732, n51733, n51734, n51735, n51736, n51737, n51738, n51740, n51741,
    n51742, n51743, n51744, n51745, n51746, n51747, n51749, n51750, n51751,
    n51752, n51753, n51754, n51755, n51756, n51758, n51759, n51760, n51761,
    n51762, n51763, n51764, n51765, n51767, n51768, n51769, n51770, n51771,
    n51772, n51773, n51774, n51776, n51777, n51778, n51779, n51780, n51781,
    n51782, n51783, n51785, n51786, n51787, n51788, n51789, n51790, n51791,
    n51792, n51794, n51795, n51796, n51797, n51798, n51799, n51800, n51801,
    n51803, n51804, n51805, n51806, n51807, n51808, n51809, n51810, n51811,
    n51812, n51814, n51815, n51816, n51817, n51818, n51819, n51821, n51822,
    n51823, n51824, n51825, n51826, n51827, n51828, n51830, n51831, n51832,
    n51833, n51834, n51835, n51836, n51838, n51839, n51840, n51841, n51842,
    n51843, n51844, n51846, n51847, n51848, n51849, n51851, n51852, n51853,
    n51854, n51855, n51856, n51857, n51858, n51859, n51860, n51861, n51862,
    n51863, n51865, n51866, n51867, n51868, n51869, n51870, n51871, n51872,
    n51873, n51874, n51875, n51876, n51877, n51879, n51880, n51881, n51882,
    n51883, n51884, n51885, n51886, n51887, n51888, n51889, n51890, n51892,
    n51893, n51894, n51895, n51896, n51898, n51899, n51900, n51901, n51902,
    n51903, n51904, n51905, n51906, n51907, n51908, n51909, n51910, n51911,
    n51912, n51913, n51914, n51915, n51916, n51917, n51918, n51919, n51920,
    n51921, n51922, n51923, n51924, n51925, n51926, n51927, n51928, n51929,
    n51930, n51931, n51932, n51933, n51934, n51935, n51936, n51937, n51938,
    n51939, n51940, n51941, n51942, n51943, n51944, n51945, n51946, n51947,
    n51948, n51949, n51950, n51951, n51952, n51953, n51954, n51955, n51956,
    n51957, n51958, n51959, n51960, n51961, n51962, n51963, n51964, n51965,
    n51966, n51967, n51968, n51969, n51970, n51971, n51972, n51973, n51974,
    n51975, n51976, n51977, n51978, n51979, n51980, n51981, n51982, n51983,
    n51984, n51985, n51986, n51987, n51988, n51989, n51990, n51991, n51992,
    n51993, n51994, n51995, n51996, n51997, n51998, n51999, n52000, n52001,
    n52002, n52003, n52004, n52005, n52006, n52007, n52008, n52009, n52010,
    n52011, n52012, n52013, n52014, n52015, n52016, n52017, n52018, n52019,
    n52020, n52021, n52022, n52023, n52024, n52025, n52026, n52027, n52028,
    n52029, n52030, n52031, n52032, n52033, n52034, n52035, n52036, n52037,
    n52038, n52039, n52040, n52041, n52042, n52043, n52044, n52045, n52046,
    n52047, n52048, n52049, n52050, n52051, n52052, n52053, n52054, n52055,
    n52056, n52057, n52058, n52059, n52060, n52061, n52062, n52063, n52064,
    n52065, n52066, n52067, n52068, n52069, n52070, n52071, n52072, n52074,
    n52075, n52076, n52077, n52078, n52079, n52080, n52081, n52082, n52083,
    n52084, n52085, n52086, n52087, n52088, n52089, n52090, n52091, n52092,
    n52093, n52094, n52095, n52096, n52097, n52098, n52099, n52100, n52101,
    n52102, n52103, n52104, n52105, n52106, n52107, n52108, n52109, n52110,
    n52111, n52112, n52113, n52114, n52115, n52116, n52117, n52118, n52119,
    n52120, n52121, n52122, n52123, n52124, n52125, n52126, n52127, n52128,
    n52129, n52130, n52131, n52132, n52133, n52134, n52135, n52136, n52137,
    n52138, n52139, n52140, n52141, n52142, n52143, n52144, n52145, n52146,
    n52147, n52148, n52149, n52150, n52151, n52152, n52153, n52154, n52155,
    n52156, n52157, n52158, n52159, n52160, n52161, n52162, n52163, n52164,
    n52165, n52166, n52167, n52168, n52169, n52170, n52171, n52172, n52173,
    n52174, n52175, n52176, n52177, n52178, n52179, n52181, n52182, n52183,
    n52184, n52185, n52186, n52187, n52188, n52189, n52190, n52191, n52192,
    n52193, n52194, n52195, n52196, n52197, n52198, n52199, n52200, n52201,
    n52202, n52203, n52204, n52205, n52206, n52207, n52208, n52209, n52210,
    n52211, n52212, n52213, n52214, n52215, n52216, n52217, n52218, n52219,
    n52220, n52221, n52222, n52223, n52224, n52225, n52226, n52227, n52228,
    n52229, n52230, n52231, n52232, n52233, n52234, n52235, n52236, n52237,
    n52238, n52239, n52240, n52241, n52242, n52243, n52244, n52245, n52246,
    n52247, n52248, n52249, n52250, n52251, n52252, n52253, n52254, n52255,
    n52256, n52257, n52258, n52259, n52260, n52261, n52262, n52263, n52264,
    n52265, n52266, n52267, n52268, n52269, n52270, n52271, n52272, n52273,
    n52274, n52275, n52276, n52277, n52278, n52279, n52280, n52281, n52282,
    n52283, n52284, n52285, n52286, n52287, n52288, n52289, n52290, n52291,
    n52292, n52293, n52294, n52295, n52296, n52297, n52298, n52299, n52300,
    n52301, n52303, n52304, n52305, n52306, n52307, n52308, n52309, n52310,
    n52311, n52312, n52313, n52314, n52315, n52316, n52317, n52318, n52319,
    n52320, n52321, n52322, n52323, n52324, n52325, n52326, n52327, n52328,
    n52329, n52330, n52331, n52332, n52333, n52334, n52335, n52336, n52337,
    n52338, n52339, n52340, n52341, n52342, n52343, n52344, n52345, n52346,
    n52347, n52348, n52349, n52350, n52351, n52352, n52353, n52354, n52355,
    n52356, n52357, n52358, n52359, n52360, n52361, n52362, n52363, n52364,
    n52365, n52366, n52367, n52368, n52369, n52370, n52371, n52372, n52373,
    n52374, n52375, n52376, n52377, n52378, n52379, n52380, n52381, n52382,
    n52383, n52384, n52385, n52386, n52387, n52388, n52389, n52390, n52391,
    n52392, n52393, n52394, n52395, n52396, n52397, n52398, n52399, n52400,
    n52401, n52402, n52403, n52404, n52405, n52406, n52407, n52408, n52409,
    n52410, n52411, n52412, n52413, n52414, n52415, n52416, n52417, n52418,
    n52419, n52420, n52421, n52422, n52423, n52424, n52425, n52426, n52427,
    n52428, n52429, n52430, n52431, n52432, n52434, n52435, n52436, n52437,
    n52438, n52439, n52440, n52441, n52442, n52443, n52444, n52445, n52446,
    n52447, n52448, n52449, n52450, n52451, n52452, n52453, n52454, n52455,
    n52456, n52457, n52458, n52459, n52460, n52461, n52462, n52463, n52464,
    n52465, n52466, n52467, n52468, n52469, n52470, n52471, n52472, n52473,
    n52474, n52475, n52476, n52477, n52478, n52479, n52480, n52481, n52482,
    n52483, n52484, n52485, n52486, n52487, n52488, n52489, n52490, n52491,
    n52492, n52493, n52494, n52495, n52496, n52497, n52498, n52499, n52500,
    n52501, n52502, n52503, n52504, n52505, n52506, n52507, n52508, n52509,
    n52510, n52511, n52512, n52513, n52514, n52515, n52516, n52517, n52518,
    n52519, n52520, n52521, n52522, n52523, n52524, n52525, n52526, n52527,
    n52528, n52529, n52530, n52531, n52532, n52533, n52534, n52535, n52536,
    n52537, n52538, n52539, n52540, n52541, n52542, n52543, n52544, n52545,
    n52546, n52547, n52548, n52549, n52550, n52551, n52552, n52553, n52554,
    n52555, n52556, n52557, n52558, n52559, n52560, n52561, n52562, n52563,
    n52564, n52565, n52566, n52567, n52568, n52570, n52571, n52572, n52573,
    n52574, n52575, n52576, n52577, n52578, n52579, n52580, n52581, n52582,
    n52583, n52584, n52585, n52586, n52587, n52588, n52589, n52590, n52591,
    n52592, n52593, n52594, n52595, n52596, n52597, n52598, n52599, n52600,
    n52601, n52602, n52603, n52604, n52605, n52606, n52607, n52608, n52609,
    n52610, n52611, n52612, n52613, n52614, n52615, n52616, n52617, n52618,
    n52619, n52620, n52621, n52622, n52623, n52624, n52625, n52626, n52627,
    n52628, n52629, n52630, n52631, n52632, n52633, n52634, n52635, n52636,
    n52637, n52638, n52639, n52640, n52641, n52642, n52643, n52644, n52645,
    n52646, n52647, n52648, n52649, n52650, n52651, n52652, n52653, n52654,
    n52655, n52656, n52657, n52658, n52659, n52660, n52661, n52662, n52663,
    n52664, n52665, n52666, n52667, n52668, n52669, n52670, n52671, n52672,
    n52673, n52674, n52675, n52676, n52677, n52678, n52679, n52680, n52681,
    n52682, n52683, n52684, n52685, n52686, n52687, n52688, n52689, n52690,
    n52691, n52692, n52693, n52694, n52695, n52696, n52697, n52698, n52699,
    n52700, n52701, n52703, n52704, n52705, n52706, n52707, n52708, n52709,
    n52710, n52711, n52712, n52713, n52714, n52715, n52716, n52717, n52718,
    n52719, n52720, n52721, n52722, n52723, n52724, n52725, n52726, n52727,
    n52728, n52729, n52730, n52731, n52732, n52733, n52734, n52735, n52736,
    n52737, n52738, n52739, n52740, n52741, n52742, n52743, n52744, n52745,
    n52746, n52747, n52748, n52749, n52750, n52751, n52752, n52753, n52754,
    n52755, n52756, n52757, n52758, n52759, n52760, n52761, n52762, n52763,
    n52764, n52765, n52766, n52767, n52768, n52769, n52770, n52771, n52772,
    n52773, n52774, n52775, n52776, n52777, n52778, n52779, n52780, n52781,
    n52782, n52783, n52784, n52785, n52786, n52787, n52788, n52789, n52790,
    n52791, n52792, n52793, n52794, n52795, n52796, n52797, n52798, n52799,
    n52800, n52801, n52802, n52803, n52804, n52805, n52806, n52807, n52808,
    n52809, n52810, n52811, n52812, n52813, n52814, n52815, n52816, n52817,
    n52818, n52819, n52820, n52821, n52822, n52823, n52824, n52825, n52826,
    n52827, n52828, n52829, n52830, n52831, n52832, n52833, n52835, n52836,
    n52837, n52838, n52839, n52840, n52841, n52842, n52843, n52844, n52845,
    n52846, n52847, n52848, n52849, n52850, n52851, n52852, n52853, n52854,
    n52855, n52856, n52857, n52858, n52859, n52860, n52861, n52862, n52863,
    n52864, n52865, n52866, n52867, n52868, n52869, n52870, n52871, n52872,
    n52873, n52874, n52875, n52876, n52877, n52878, n52879, n52880, n52881,
    n52882, n52883, n52884, n52885, n52886, n52887, n52888, n52889, n52890,
    n52891, n52892, n52893, n52894, n52895, n52896, n52897, n52898, n52899,
    n52900, n52901, n52902, n52903, n52904, n52905, n52906, n52907, n52908,
    n52909, n52910, n52911, n52912, n52913, n52914, n52915, n52916, n52917,
    n52918, n52919, n52920, n52921, n52922, n52923, n52924, n52925, n52926,
    n52927, n52928, n52929, n52930, n52931, n52932, n52933, n52934, n52935,
    n52936, n52937, n52939, n52940, n52941, n52942, n52943, n52944, n52945,
    n52946, n52947, n52948, n52949, n52950, n52951, n52952, n52953, n52954,
    n52955, n52956, n52957, n52958, n52959, n52960, n52961, n52962, n52963,
    n52964, n52965, n52966, n52967, n52968, n52969, n52970, n52971, n52972,
    n52973, n52974, n52975, n52976, n52977, n52978, n52979, n52980, n52981,
    n52982, n52983, n52984, n52985, n52986, n52987, n52988, n52989, n52990,
    n52991, n52992, n52993, n52994, n52995, n52996, n52997, n52998, n52999,
    n53000, n53001, n53002, n53003, n53004, n53005, n53006, n53007, n53008,
    n53009, n53010, n53011, n53012, n53013, n53014, n53015, n53016, n53017,
    n53018, n53019, n53020, n53021, n53022, n53023, n53024, n53025, n53026,
    n53027, n53029, n53030, n53031, n53032, n53033, n53034, n53035, n53036,
    n53037, n53038, n53039, n53040, n53041, n53042, n53043, n53044, n53045,
    n53046, n53047, n53048, n53049, n53050, n53051, n53052, n53053, n53054,
    n53055, n53056, n53057, n53058, n53059, n53060, n53061, n53062, n53063,
    n53064, n53065, n53066, n53067, n53068, n53069, n53070, n53071, n53072,
    n53073, n53074, n53075, n53076, n53077, n53078, n53079, n53080, n53081,
    n53082, n53083, n53084, n53085, n53086, n53087, n53088, n53089, n53090,
    n53091, n53092, n53093, n53094, n53095, n53096, n53097, n53098, n53099,
    n53100, n53101, n53102, n53103, n53104, n53105, n53106, n53107, n53108,
    n53109, n53110, n53112, n53113, n53114, n53115, n53116, n53117, n53118,
    n53119, n53120, n53121, n53122, n53123, n53124, n53125, n53126, n53127,
    n53128, n53129, n53130, n53131, n53132, n53133, n53134, n53135, n53136,
    n53137, n53138, n53139, n53140, n53141, n53142, n53143, n53144, n53145,
    n53146, n53147, n53148, n53149, n53150, n53151, n53152, n53153, n53154,
    n53155, n53156, n53157, n53158, n53159, n53160, n53161, n53162, n53163,
    n53164, n53165, n53166, n53167, n53168, n53169, n53170, n53171, n53172,
    n53173, n53174, n53175, n53176, n53177, n53178, n53179, n53180, n53181,
    n53182, n53183, n53184, n53185, n53186, n53188, n53189, n53190, n53191,
    n53192, n53193, n53194, n53195, n53196, n53197, n53198, n53199, n53200,
    n53201, n53202, n53203, n53204, n53205, n53206, n53207, n53208, n53209,
    n53210, n53211, n53212, n53213, n53214, n53215, n53216, n53217, n53218,
    n53219, n53220, n53221, n53222, n53223, n53224, n53225, n53226, n53227,
    n53228, n53229, n53230, n53231, n53232, n53233, n53234, n53235, n53236,
    n53237, n53238, n53239, n53240, n53241, n53242, n53243, n53244, n53245,
    n53246, n53247, n53248, n53249, n53250, n53251, n53252, n53253, n53254,
    n53255, n53256, n53257, n53258, n53260, n53261, n53262, n53263, n53264,
    n53265, n53266, n53267, n53268, n53269, n53270, n53271, n53272, n53273,
    n53274, n53275, n53276, n53277, n53278, n53279, n53280, n53281, n53282,
    n53283, n53284, n53285, n53286, n53287, n53288, n53289, n53290, n53291,
    n53292, n53293, n53294, n53295, n53296, n53297, n53298, n53299, n53300,
    n53301, n53302, n53303, n53304, n53305, n53306, n53307, n53308, n53309,
    n53310, n53311, n53312, n53313, n53314, n53315, n53316, n53317, n53318,
    n53319, n53320, n53321, n53322, n53323, n53324, n53325, n53326, n53327,
    n53328, n53329, n53330, n53331, n53332, n53333, n53334, n53335, n53336,
    n53337, n53339, n53340, n53341, n53342, n53343, n53344, n53345, n53346,
    n53347, n53348, n53349, n53350, n53351, n53352, n53353, n53354, n53355,
    n53356, n53357, n53358, n53359, n53360, n53361, n53362, n53363, n53364,
    n53365, n53366, n53367, n53368, n53369, n53370, n53371, n53372, n53373,
    n53374, n53375, n53376, n53377, n53378, n53379, n53380, n53381, n53382,
    n53383, n53384, n53385, n53386, n53387, n53388, n53389, n53390, n53391,
    n53392, n53393, n53394, n53395, n53396, n53397, n53398, n53399, n53400,
    n53401, n53402, n53403, n53404, n53405, n53406, n53407, n53408, n53409,
    n53410, n53411, n53412, n53414, n53415, n53416, n53417, n53418, n53419,
    n53420, n53421, n53422, n53423, n53424, n53425, n53426, n53427, n53428,
    n53429, n53430, n53431, n53432, n53433, n53434, n53435, n53436, n53437,
    n53438, n53439, n53440, n53441, n53442, n53443, n53444, n53445, n53446,
    n53447, n53448, n53449, n53450, n53451, n53452, n53453, n53454, n53455,
    n53456, n53457, n53458, n53459, n53460, n53461, n53462, n53463, n53464,
    n53465, n53466, n53467, n53468, n53469, n53470, n53471, n53472, n53473,
    n53474, n53475, n53476, n53477, n53478, n53479, n53480, n53481, n53482,
    n53483, n53484, n53485, n53487, n53488, n53489, n53490, n53491, n53492,
    n53493, n53494, n53495, n53496, n53497, n53498, n53499, n53500, n53501,
    n53502, n53503, n53504, n53505, n53506, n53507, n53508, n53509, n53510,
    n53511, n53512, n53513, n53514, n53515, n53516, n53517, n53518, n53519,
    n53520, n53521, n53522, n53523, n53524, n53525, n53526, n53527, n53528,
    n53529, n53530, n53531, n53532, n53533, n53534, n53535, n53536, n53537,
    n53538, n53539, n53540, n53541, n53542, n53543, n53544, n53545, n53546,
    n53547, n53548, n53549, n53550, n53551, n53552, n53553, n53554, n53555,
    n53556, n53557, n53558, n53559, n53560, n53561, n53562, n53563, n53565,
    n53566, n53567, n53568, n53569, n53570, n53571, n53572, n53573, n53574,
    n53575, n53576, n53577, n53578, n53579, n53580, n53581, n53582, n53583,
    n53584, n53585, n53586, n53587, n53588, n53589, n53590, n53591, n53592,
    n53593, n53594, n53595, n53596, n53597, n53598, n53599, n53600, n53601,
    n53602, n53603, n53604, n53605, n53606, n53607, n53608, n53609, n53610,
    n53611, n53612, n53613, n53614, n53615, n53616, n53617, n53618, n53619,
    n53620, n53621, n53622, n53623, n53624, n53625, n53626, n53627, n53628,
    n53629, n53630, n53631, n53632, n53633, n53634, n53635, n53637, n53638,
    n53639, n53640, n53641, n53642, n53643, n53644, n53645, n53646, n53647,
    n53648, n53649, n53650, n53651, n53652, n53653, n53654, n53655, n53656,
    n53657, n53658, n53659, n53660, n53661, n53662, n53663, n53664, n53665,
    n53666, n53667, n53668, n53669, n53670, n53671, n53672, n53673, n53674,
    n53675, n53676, n53677, n53678, n53679, n53680, n53681, n53682, n53683,
    n53684, n53685, n53686, n53687, n53688, n53689, n53690, n53691, n53692,
    n53693, n53694, n53695, n53696, n53697, n53698, n53699, n53700, n53701,
    n53702, n53703, n53704, n53705, n53706, n53707, n53708, n53709, n53710,
    n53711, n53712, n53713, n53714, n53716, n53717, n53718, n53719, n53720,
    n53721, n53722, n53723, n53724, n53725, n53726, n53727, n53728, n53729,
    n53730, n53731, n53732, n53733, n53734, n53735, n53736, n53737, n53738,
    n53739, n53740, n53741, n53742, n53743, n53744, n53745, n53746, n53747,
    n53748, n53749, n53750, n53751, n53752, n53753, n53754, n53755, n53756,
    n53757, n53758, n53759, n53760, n53761, n53762, n53763, n53764, n53765,
    n53766, n53767, n53768, n53769, n53770, n53771, n53772, n53773, n53774,
    n53775, n53776, n53777, n53778, n53779, n53780, n53781, n53782, n53783,
    n53784, n53785, n53787, n53788, n53789, n53790, n53791, n53792, n53793,
    n53794, n53795, n53796, n53797, n53798, n53799, n53800, n53801, n53802,
    n53803, n53804, n53805, n53806, n53807, n53808, n53809, n53810, n53811,
    n53812, n53813, n53814, n53815, n53816, n53817, n53818, n53819, n53820,
    n53821, n53822, n53823, n53824, n53825, n53826, n53827, n53828, n53829,
    n53830, n53831, n53832, n53833, n53834, n53835, n53836, n53837, n53838,
    n53839, n53840, n53841, n53842, n53843, n53844, n53845, n53846, n53847,
    n53848, n53849, n53850, n53851, n53852, n53853, n53854, n53855, n53856,
    n53857, n53858, n53859, n53860, n53861, n53862, n53863, n53864, n53865,
    n53867, n53868, n53869, n53870, n53871, n53872, n53873, n53874, n53875,
    n53876, n53877, n53878, n53879, n53880, n53881, n53882, n53883, n53884,
    n53885, n53886, n53887, n53888, n53889, n53890, n53891, n53892, n53893,
    n53894, n53895, n53896, n53897, n53898, n53899, n53900, n53901, n53902,
    n53903, n53904, n53905, n53906, n53907, n53908, n53909, n53910, n53911,
    n53912, n53913, n53914, n53915, n53916, n53917, n53918, n53919, n53920,
    n53921, n53922, n53923, n53924, n53925, n53926, n53927, n53928, n53929,
    n53930, n53931, n53932, n53933, n53934, n53935, n53936, n53937, n53938,
    n53939, n53940, n53941, n53943, n53944, n53945, n53946, n53947, n53948,
    n53949, n53950, n53951, n53952, n53953, n53954, n53955, n53956, n53957,
    n53958, n53959, n53960, n53961, n53962, n53963, n53964, n53965, n53966,
    n53967, n53968, n53969, n53970, n53971, n53972, n53973, n53974, n53975,
    n53976, n53977, n53978, n53979, n53980, n53981, n53982, n53983, n53984,
    n53985, n53986, n53987, n53988, n53989, n53990, n53991, n53992, n53993,
    n53994, n53995, n53996, n53997, n53998, n53999, n54000, n54001, n54002,
    n54003, n54004, n54005, n54006, n54007, n54008, n54009, n54010, n54011,
    n54012, n54013, n54014, n54016, n54017, n54018, n54019, n54020, n54021,
    n54022, n54023, n54024, n54025, n54026, n54027, n54028, n54029, n54030,
    n54031, n54032, n54033, n54034, n54035, n54036, n54037, n54038, n54039,
    n54040, n54041, n54042, n54043, n54044, n54045, n54046, n54047, n54048,
    n54049, n54050, n54051, n54052, n54053, n54054, n54055, n54056, n54057,
    n54058, n54059, n54060, n54061, n54062, n54063, n54064, n54065, n54066,
    n54067, n54068, n54069, n54070, n54071, n54072, n54073, n54074, n54075,
    n54076, n54077, n54078, n54079, n54080, n54081, n54082, n54083, n54084,
    n54085, n54086, n54087, n54088, n54089, n54090, n54091, n54093, n54094,
    n54095, n54096, n54097, n54098, n54099, n54100, n54101, n54102, n54103,
    n54104, n54105, n54106, n54107, n54108, n54109, n54110, n54111, n54112,
    n54113, n54114, n54115, n54116, n54117, n54118, n54119, n54120, n54121,
    n54122, n54123, n54124, n54125, n54126, n54127, n54128, n54129, n54130,
    n54131, n54132, n54133, n54134, n54135, n54136, n54137, n54138, n54139,
    n54140, n54141, n54142, n54143, n54144, n54145, n54146, n54147, n54148,
    n54149, n54150, n54151, n54152, n54153, n54154, n54155, n54156, n54157,
    n54158, n54159, n54160, n54161, n54162, n54163, n54164, n54165, n54166,
    n54167, n54168, n54169, n54170, n54172, n54173, n54174, n54175, n54176,
    n54177, n54178, n54179, n54180, n54181, n54182, n54183, n54184, n54185,
    n54186, n54187, n54188, n54189, n54190, n54191, n54192, n54193, n54194,
    n54195, n54196, n54197, n54198, n54199, n54200, n54201, n54202, n54203,
    n54204, n54205, n54206, n54207, n54208, n54209, n54210, n54211, n54212,
    n54213, n54214, n54215, n54216, n54217, n54218, n54219, n54220, n54221,
    n54222, n54223, n54224, n54225, n54226, n54227, n54228, n54229, n54230,
    n54231, n54232, n54233, n54234, n54235, n54236, n54237, n54238, n54239,
    n54240, n54241, n54242, n54243, n54244, n54246, n54247, n54248, n54249,
    n54250, n54251, n54252, n54253, n54254, n54255, n54256, n54257, n54258,
    n54259, n54260, n54261, n54262, n54263, n54264, n54265, n54266, n54267,
    n54268, n54269, n54270, n54271, n54272, n54273, n54274, n54275, n54276,
    n54277, n54278, n54279, n54280, n54281, n54282, n54283, n54284, n54285,
    n54286, n54287, n54288, n54289, n54290, n54291, n54292, n54293, n54294,
    n54295, n54296, n54297, n54298, n54299, n54300, n54301, n54302, n54303,
    n54304, n54305, n54306, n54307, n54308, n54309, n54310, n54311, n54312,
    n54313, n54314, n54315, n54316, n54317, n54318, n54319, n54320, n54321,
    n54322, n54323, n54324, n54326, n54327, n54328, n54329, n54330, n54331,
    n54332, n54333, n54334, n54335, n54336, n54337, n54338, n54339, n54340,
    n54341, n54342, n54343, n54344, n54345, n54346, n54347, n54348, n54349,
    n54350, n54351, n54352, n54353, n54354, n54355, n54356, n54357, n54358,
    n54359, n54360, n54361, n54362, n54363, n54364, n54365, n54366, n54367,
    n54368, n54369, n54370, n54371, n54372, n54373, n54374, n54375, n54376,
    n54377, n54378, n54379, n54380, n54381, n54382, n54383, n54384, n54385,
    n54386, n54387, n54388, n54389, n54390, n54391, n54392, n54393, n54394,
    n54395, n54396, n54397, n54398, n54399, n54401, n54402, n54403, n54404,
    n54405, n54406, n54407, n54408, n54409, n54410, n54411, n54412, n54413,
    n54414, n54415, n54416, n54417, n54418, n54419, n54420, n54421, n54422,
    n54423, n54424, n54425, n54426, n54427, n54428, n54429, n54430, n54431,
    n54432, n54433, n54434, n54435, n54436, n54437, n54438, n54439, n54440,
    n54441, n54442, n54443, n54444, n54445, n54446, n54447, n54448, n54449,
    n54450, n54451, n54452, n54453, n54454, n54455, n54456, n54457, n54458,
    n54459, n54460, n54461, n54462, n54463, n54464, n54465, n54466, n54467,
    n54468, n54469, n54470, n54472, n54473, n54474, n54475, n54476, n54477,
    n54478, n54479, n54480, n54481, n54482, n54483, n54484, n54485, n54486,
    n54487, n54488, n54489, n54490, n54491, n54492, n54493, n54494, n54495,
    n54496, n54497, n54498, n54499, n54500, n54501, n54502, n54503, n54504,
    n54505, n54506, n54507, n54508, n54509, n54510, n54511, n54512, n54513,
    n54514, n54515, n54516, n54517, n54518, n54519, n54520, n54521, n54522,
    n54523, n54524, n54525, n54526, n54527, n54528, n54529, n54530, n54531,
    n54532, n54533, n54534, n54535, n54536, n54537, n54538, n54539, n54540,
    n54541, n54542, n54543, n54544, n54545, n54546, n54547, n54548, n54549,
    n54550, n54551, n54552, n54553, n54554, n54555, n54557, n54558, n54559,
    n54560, n54561, n54562, n54563, n54564, n54565, n54566, n54567, n54568,
    n54569, n54570, n54571, n54572, n54573, n54574, n54575, n54576, n54577,
    n54578, n54579, n54580, n54581, n54582, n54583, n54584, n54585, n54586,
    n54587, n54588, n54589, n54590, n54591, n54592, n54593, n54594, n54595,
    n54596, n54597, n54598, n54599, n54600, n54601, n54602, n54603, n54604,
    n54605, n54606, n54607, n54608, n54609, n54610, n54611, n54612, n54613,
    n54614, n54615, n54616, n54617, n54618, n54619, n54620, n54621, n54622,
    n54623, n54624, n54625, n54626, n54628, n54629, n54630, n54631, n54632,
    n54633, n54634, n54635, n54636, n54637, n54638, n54639, n54640, n54641,
    n54642, n54643, n54644, n54645, n54646, n54647, n54648, n54649, n54650,
    n54651, n54652, n54653, n54654, n54655, n54656, n54657, n54658, n54659,
    n54660, n54661, n54662, n54663, n54664, n54665, n54666, n54667, n54668,
    n54669, n54670, n54671, n54672, n54673, n54674, n54675, n54676, n54677,
    n54678, n54679, n54680, n54681, n54682, n54683, n54684, n54685, n54686,
    n54687, n54688, n54689, n54690, n54691, n54692, n54693, n54694, n54695,
    n54696, n54697, n54698, n54700, n54701, n54702, n54703, n54704, n54705,
    n54706, n54707, n54708, n54709, n54710, n54711, n54712, n54713, n54714,
    n54715, n54716, n54717, n54718, n54719, n54720, n54721, n54722, n54723,
    n54724, n54725, n54726, n54727, n54728, n54729, n54730, n54731, n54732,
    n54733, n54734, n54735, n54736, n54737, n54738, n54739, n54740, n54741,
    n54742, n54743, n54744, n54745, n54746, n54747, n54748, n54749, n54750,
    n54751, n54752, n54753, n54754, n54755, n54756, n54757, n54758, n54759,
    n54760, n54761, n54762, n54763, n54764, n54765, n54766, n54767, n54768,
    n54769, n54770, n54771, n54772, n54773, n54774, n54775, n54776, n54777,
    n54778, n54779, n54780, n54781, n54783, n54784, n54785, n54786, n54787,
    n54788, n54789, n54790, n54791, n54792, n54793, n54794, n54795, n54796,
    n54797, n54798, n54799, n54800, n54801, n54802, n54803, n54804, n54805,
    n54806, n54807, n54808, n54809, n54810, n54811, n54812, n54813, n54814,
    n54816, n54817, n54818, n54819, n54820, n54821, n54822, n54823, n54824,
    n54825, n54826, n54827, n54828, n54829, n54831, n54832, n54833, n54834,
    n54835, n54836, n54837, n54838, n54839, n54840, n54841, n54842, n54843,
    n54844, n54845, n54846, n54847, n54849, n54850, n54851, n54852, n54853,
    n54854, n54855, n54856, n54857, n54858, n54859, n54860, n54861, n54862,
    n54863, n54864, n54865, n54866, n54867, n54868, n54869, n54871, n54872,
    n54873, n54874, n54875, n54876, n54877, n54878, n54879, n54880, n54881,
    n54882, n54883, n54884, n54885, n54886, n54887, n54888, n54889, n54890,
    n54891, n54892, n54894, n54895, n54896, n54897, n54898, n54899, n54900,
    n54901, n54902, n54903, n54904, n54905, n54906, n54907, n54908, n54909,
    n54910, n54911, n54912, n54913, n54914, n54915, n54917, n54918, n54919,
    n54920, n54921, n54922, n54923, n54924, n54925, n54926, n54927, n54928,
    n54929, n54930, n54931, n54932, n54933, n54934, n54935, n54936, n54937,
    n54938, n54940, n54941, n54942, n54943, n54944, n54945, n54946, n54947,
    n54948, n54949, n54950, n54951, n54952, n54953, n54954, n54955, n54956,
    n54957, n54958, n54959, n54960, n54961, n54963, n54964, n54965, n54966,
    n54967, n54968, n54969, n54970, n54971, n54972, n54973, n54974, n54975,
    n54976, n54977, n54978, n54979, n54980, n54981, n54982, n54983, n54984,
    n54986, n54987, n54988, n54989, n54990, n54991, n54992, n54993, n54994,
    n54995, n54996, n54997, n54998, n54999, n55000, n55001, n55002, n55003,
    n55004, n55005, n55006, n55007, n55009, n55010, n55011, n55012, n55013,
    n55014, n55015, n55016, n55017, n55018, n55019, n55020, n55021, n55022,
    n55023, n55024, n55025, n55026, n55027, n55028, n55029, n55030, n55032,
    n55033, n55034, n55035, n55036, n55037, n55038, n55039, n55040, n55041,
    n55042, n55043, n55044, n55045, n55046, n55047, n55048, n55049, n55050,
    n55051, n55052, n55053, n55055, n55056, n55057, n55058, n55059, n55060,
    n55061, n55062, n55063, n55064, n55065, n55066, n55067, n55068, n55069,
    n55070, n55071, n55072, n55073, n55074, n55075, n55076, n55078, n55079,
    n55080, n55081, n55082, n55083, n55084, n55085, n55086, n55087, n55088,
    n55089, n55090, n55091, n55092, n55093, n55094, n55095, n55096, n55097,
    n55098, n55099, n55101, n55102, n55103, n55104, n55105, n55106, n55107,
    n55108, n55109, n55110, n55111, n55112, n55113, n55114, n55115, n55116,
    n55117, n55118, n55119, n55120, n55121, n55122, n55124, n55125, n55126,
    n55127, n55128, n55129, n55130, n55131, n55132, n55133, n55134, n55135,
    n55136, n55137, n55138, n55139, n55140, n55141, n55142, n55143, n55144,
    n55145, n55147, n55148, n55149, n55150, n55151, n55152, n55153, n55154,
    n55155, n55156, n55157, n55158, n55159, n55160, n55161, n55162, n55163,
    n55164, n55165, n55166, n55167, n55168, n55170, n55171, n55172, n55173,
    n55174, n55175, n55176, n55177, n55178, n55179, n55180, n55181, n55182,
    n55183, n55184, n55185, n55186, n55187, n55188, n55189, n55190, n55191,
    n55193, n55194, n55195, n55196, n55197, n55198, n55199, n55200, n55201,
    n55202, n55203, n55204, n55205, n55206, n55207, n55208, n55209, n55210,
    n55211, n55212, n55213, n55214, n55216, n55217, n55218, n55219, n55220,
    n55221, n55222, n55223, n55224, n55225, n55226, n55227, n55228, n55229,
    n55230, n55231, n55232, n55233, n55234, n55235, n55236, n55237, n55239,
    n55240, n55241, n55242, n55243, n55244, n55245, n55246, n55247, n55248,
    n55249, n55250, n55251, n55252, n55253, n55254, n55255, n55256, n55257,
    n55258, n55259, n55260, n55262, n55263, n55264, n55265, n55266, n55267,
    n55268, n55269, n55270, n55271, n55272, n55273, n55274, n55275, n55276,
    n55277, n55278, n55279, n55280, n55281, n55282, n55283, n55285, n55286,
    n55287, n55288, n55289, n55290, n55291, n55292, n55293, n55294, n55295,
    n55296, n55297, n55298, n55299, n55300, n55301, n55302, n55303, n55304,
    n55305, n55306, n55308, n55309, n55310, n55311, n55312, n55313, n55314,
    n55315, n55316, n55317, n55318, n55319, n55320, n55321, n55322, n55323,
    n55324, n55325, n55326, n55327, n55328, n55329, n55331, n55332, n55333,
    n55334, n55335, n55336, n55337, n55338, n55339, n55340, n55341, n55342,
    n55343, n55344, n55345, n55346, n55347, n55348, n55349, n55350, n55351,
    n55352, n55354, n55355, n55356, n55357, n55358, n55359, n55360, n55361,
    n55362, n55363, n55364, n55365, n55366, n55367, n55368, n55369, n55370,
    n55371, n55372, n55373, n55374, n55375, n55377, n55378, n55379, n55380,
    n55381, n55382, n55383, n55384, n55385, n55386, n55387, n55388, n55389,
    n55390, n55391, n55392, n55393, n55394, n55395, n55396, n55397, n55398,
    n55400, n55401, n55402, n55403, n55404, n55405, n55406, n55407, n55408,
    n55409, n55410, n55411, n55412, n55413, n55414, n55415, n55416, n55417,
    n55418, n55419, n55420, n55421, n55423, n55424, n55425, n55426, n55427,
    n55428, n55429, n55430, n55431, n55432, n55433, n55434, n55435, n55436,
    n55437, n55438, n55439, n55440, n55441, n55442, n55443, n55444, n55446,
    n55447, n55448, n55449, n55450, n55451, n55452, n55453, n55454, n55455,
    n55456, n55457, n55458, n55459, n55460, n55461, n55462, n55463, n55464,
    n55465, n55466, n55467, n55469, n55470, n55471, n55472, n55473, n55474,
    n55475, n55476, n55477, n55478, n55479, n55480, n55481, n55482, n55483,
    n55484, n55485, n55486, n55487, n55488, n55489, n55490, n55492, n55493,
    n55494, n55495, n55496, n55497, n55498, n55499, n55500, n55501, n55502,
    n55503, n55504, n55505, n55506, n55507, n55508, n55509, n55510, n55511,
    n55512, n55513, n55515, n55516, n55517, n55518, n55519, n55520, n55521,
    n55522, n55523, n55524, n55525, n55526, n55527, n55528, n55529, n55530,
    n55531, n55532, n55533, n55534, n55536, n55537, n55538, n55539, n55540,
    n55541, n55542, n55543, n55544, n55545, n55546, n55547, n55548, n55549,
    n55550, n55552, n55553, n55554, n55555, n55556, n55557, n55558, n55559,
    n55560, n55561, n55562, n55563, n55564, n55566, n55567, n55568, n55569,
    n55570, n55571, n55572, n55573, n55574, n55575, n55576, n55577, n55578,
    n55579, n55580, n55582, n55583, n55584, n55585, n55586, n55587, n55588,
    n55589, n55590, n55591, n55592, n55593, n55594, n55595, n55597, n55598,
    n55599, n55600, n55601, n55602, n55603, n55604, n55605, n55606, n55607,
    n55608, n55609, n55610, n55611, n55613, n55614, n55615, n55616, n55617,
    n55618, n55619, n55620, n55621, n55622, n55623, n55625, n55626, n55627,
    n55628, n55629, n55630, n55631, n55632, n55633, n55634, n55635, n55636,
    n55637, n55638, n55639, n55640, n55642, n55643, n55644, n55645, n55647,
    n55648, n55649, n55650, n55652, n55653, n55654, n55655, n55657, n55658,
    n55659, n55660, n55662, n55663, n55664, n55665, n55667, n55668, n55669,
    n55670, n55672, n55673, n55674, n55675, n55677, n55678, n55679, n55680,
    n55682, n55683, n55684, n55686, n55687, n55688, n55690, n55691, n55692,
    n55694, n55695, n55696, n55698, n55699, n55700, n55702, n55703, n55704,
    n55706, n55707, n55708, n55710, n55711, n55712, n55714, n55715, n55716,
    n55718, n55719, n55720, n55722, n55723, n55724, n55726, n55727, n55728,
    n55730, n55731, n55732, n55734, n55735, n55736, n55738, n55739, n55740,
    n55742, n55743, n55744, n55745, n55746, n55747, n55748, n55749, n55750,
    n55751, n55753, n55754, n55755, n55756, n55758, n55759, n55760, n55761,
    n55763, n55764, n55765, n55766, n55768, n55769, n55770, n55771, n55773,
    n55774, n55775, n55776, n55778, n55779, n55780, n55781, n55783, n55784,
    n55785, n55786, n55788, n55789, n55790, n55791, n55793, n55794, n55795,
    n55796, n55798, n55799, n55800, n55801, n55803, n55804, n55805, n55806,
    n55808, n55809, n55810, n55811, n55813, n55814, n55815, n55816, n55818,
    n55819, n55820, n55821, n55823, n55824, n55825, n55826, n55828, n55829,
    n55830, n55831, n55832, n55834, n55835, n55836, n55837, n55839, n55840,
    n55841, n55842, n55844, n55845, n55846, n55847, n55849, n55850, n55851,
    n55852, n55854, n55855, n55856, n55857, n55859, n55860, n55861, n55862,
    n55864, n55865, n55866, n55867, n55869, n55870, n55871, n55872, n55874,
    n55875, n55876, n55877, n55879, n55880, n55881, n55882, n55884, n55885,
    n55886, n55887, n55889, n55890, n55891, n55892, n55894, n55895, n55896,
    n55897, n55899, n55900, n55901, n55902, n55905, n55906, n55907, n55908,
    n55909, n55910, n55911, n55912, n55913, n55914, n55915, n55916, n55918,
    n55919, n55920, n55921, n55922, n55923, n55924, n55925, n55926, n55928,
    n55929, n55930, n55931, n55932, n55933, n55934, n55935, n55936, n55937,
    n55939, n55940, n55941, n55942, n55943, n55944, n55945, n55946, n55947,
    n55948, n55950, n55951, n55952, n55953, n55954, n55955, n55956, n55957,
    n55958, n55959, n55961, n55962, n55963, n55964, n55965, n55966, n55967,
    n55968, n55969, n55970, n55972, n55973, n55974, n55975, n55976, n55977,
    n55978, n55979, n55980, n55981, n55983, n55984, n55985, n55986, n55987,
    n55988, n55989, n55990, n55991, n55992, n55994, n55995, n55996, n55997,
    n55998, n55999, n56000, n56001, n56002, n56003, n56004, n56005, n56006,
    n56007, n56008, n56009, n56010, n56011, n56012, n56013, n56014, n56015,
    n56016, n56017, n56018, n56019, n56020, n56021, n56022, n56023, n56024,
    n56025, n56026, n56027, n56028, n56029, n56030, n56031, n56032, n56033,
    n56034, n56035, n56036, n56037, n56038, n56039, n56040, n56041, n56042,
    n56043, n56044, n56045, n56046, n56047, n56048, n56049, n56050, n56051,
    n56052, n56053, n56054, n56055, n56057, n56058, n56059, n56060, n56061,
    n56062, n56063, n56064, n56065, n56066, n56067, n56068, n56069, n56070,
    n56071, n56072, n56073, n56074, n56075, n56076, n56077, n56078, n56079,
    n56080, n56081, n56082, n56083, n56084, n56085, n56086, n56087, n56088,
    n56089, n56090, n56091, n56092, n56093, n56094, n56095, n56096, n56097,
    n56099, n56100, n56101, n56102, n56103, n56104, n56105, n56106, n56107,
    n56108, n56109, n56110, n56111, n56112, n56113, n56114, n56115, n56116,
    n56117, n56118, n56119, n56120, n56121, n56122, n56123, n56124, n56125,
    n56126, n56127, n56128, n56129, n56130, n56131, n56132, n56133, n56134,
    n56135, n56136, n56137, n56138, n56139, n56141, n56142, n56143, n56144,
    n56145, n56146, n56147, n56148, n56149, n56150, n56151, n56152, n56153,
    n56154, n56155, n56156, n56157, n56158, n56159, n56160, n56161, n56162,
    n56163, n56164, n56165, n56166, n56167, n56168, n56169, n56170, n56171,
    n56172, n56173, n56174, n56175, n56176, n56177, n56178, n56179, n56180,
    n56181, n56183, n56184, n56185, n56186, n56187, n56188, n56189, n56190,
    n56191, n56192, n56193, n56194, n56195, n56196, n56197, n56198, n56199,
    n56200, n56201, n56202, n56203, n56204, n56205, n56206, n56207, n56208,
    n56209, n56210, n56211, n56212, n56213, n56214, n56215, n56216, n56217,
    n56218, n56219, n56220, n56221, n56222, n56223, n56225, n56226, n56227,
    n56228, n56229, n56230, n56231, n56232, n56233, n56234, n56235, n56236,
    n56237, n56238, n56239, n56240, n56241, n56242, n56243, n56244, n56245,
    n56246, n56247, n56248, n56249, n56250, n56251, n56252, n56253, n56254,
    n56255, n56256, n56257, n56258, n56259, n56260, n56261, n56262, n56263,
    n56264, n56265, n56267, n56268, n56269, n56270, n56271, n56272, n56273,
    n56274, n56275, n56276, n56277, n56278, n56279, n56280, n56281, n56282,
    n56283, n56284, n56285, n56286, n56287, n56288, n56289, n56290, n56291,
    n56292, n56293, n56294, n56295, n56296, n56297, n56298, n56299, n56300,
    n56301, n56302, n56303, n56304, n56305, n56306, n56307, n56309, n56310,
    n56311, n56312, n56313, n56314, n56315, n56316, n56317, n56318, n56319,
    n56320, n56321, n56322, n56323, n56324, n56325, n56326, n56327, n56328,
    n56329, n56330, n56331, n56332, n56333, n56334, n56335, n56336, n56337,
    n56338, n56339, n56340, n56341, n56342, n56343, n56344, n56345, n56346,
    n56347, n56348, n56349, n56351, n56352, n56353, n56354, n56355, n56356,
    n56357, n56358, n56359, n56360, n56361, n56362, n56363, n56364, n56365,
    n56366, n56367, n56368, n56369, n56370, n56371, n56372, n56373, n56374,
    n56375, n56376, n56377, n56378, n56379, n56380, n56381, n56382, n56383,
    n56384, n56385, n56386, n56387, n56388, n56389, n56390, n56391, n56392,
    n56393, n56394, n56395, n56396, n56397, n56398, n56399, n56400, n56401,
    n56402, n56403, n56404, n56405, n56406, n56407, n56408, n56409, n56410,
    n56411, n56412, n56413, n56414, n56415, n56416, n56417, n56418, n56419,
    n56420, n56422, n56423, n56424, n56425, n56426, n56427, n56428, n56429,
    n56430, n56431, n56432, n56433, n56434, n56435, n56436, n56437, n56438,
    n56439, n56440, n56441, n56442, n56443, n56444, n56445, n56446, n56447,
    n56448, n56449, n56450, n56451, n56452, n56453, n56454, n56455, n56456,
    n56457, n56458, n56459, n56460, n56461, n56462, n56463, n56464, n56466,
    n56467, n56468, n56469, n56470, n56471, n56472, n56473, n56474, n56475,
    n56476, n56477, n56478, n56479, n56480, n56481, n56482, n56483, n56484,
    n56485, n56486, n56487, n56488, n56489, n56490, n56491, n56492, n56493,
    n56494, n56495, n56496, n56497, n56498, n56499, n56500, n56501, n56502,
    n56503, n56504, n56505, n56506, n56507, n56508, n56510, n56511, n56512,
    n56513, n56514, n56515, n56516, n56517, n56518, n56519, n56520, n56521,
    n56522, n56523, n56524, n56525, n56526, n56527, n56528, n56529, n56530,
    n56531, n56532, n56533, n56534, n56535, n56536, n56537, n56538, n56539,
    n56540, n56541, n56542, n56543, n56544, n56545, n56546, n56547, n56548,
    n56549, n56550, n56551, n56552, n56554, n56555, n56556, n56557, n56558,
    n56559, n56560, n56561, n56562, n56563, n56564, n56565, n56566, n56567,
    n56568, n56569, n56570, n56571, n56572, n56573, n56574, n56575, n56576,
    n56577, n56578, n56579, n56580, n56581, n56582, n56583, n56584, n56585,
    n56586, n56587, n56588, n56589, n56590, n56591, n56592, n56593, n56594,
    n56595, n56596, n56598, n56599, n56600, n56601, n56602, n56603, n56604,
    n56605, n56606, n56607, n56608, n56609, n56610, n56611, n56612, n56613,
    n56614, n56615, n56616, n56617, n56618, n56619, n56620, n56621, n56622,
    n56623, n56624, n56625, n56626, n56627, n56628, n56629, n56630, n56631,
    n56632, n56633, n56634, n56635, n56636, n56637, n56638, n56639, n56640,
    n56642, n56643, n56644, n56645, n56646, n56647, n56648, n56649, n56650,
    n56651, n56652, n56653, n56654, n56655, n56656, n56657, n56658, n56659,
    n56660, n56661, n56662, n56663, n56664, n56665, n56666, n56667, n56668,
    n56669, n56670, n56671, n56672, n56673, n56674, n56675, n56676, n56677,
    n56678, n56679, n56680, n56681, n56682, n56683, n56684, n56686, n56687,
    n56688, n56689, n56690, n56691, n56692, n56693, n56694, n56695, n56696,
    n56697, n56698, n56699, n56700, n56701, n56702, n56703, n56704, n56705,
    n56706, n56707, n56708, n56709, n56710, n56711, n56712, n56713, n56714,
    n56715, n56716, n56717, n56718, n56719, n56720, n56721, n56722, n56723,
    n56724, n56725, n56726, n56727, n56728, n56729, n56730, n56731, n56732,
    n56733, n56734, n56735, n56736, n56737, n56738, n56739, n56740, n56741,
    n56742, n56743, n56744, n56745, n56746, n56747, n56748, n56749, n56750,
    n56751, n56752, n56753, n56754, n56755, n56756, n56757, n56758, n56759,
    n56760, n56761, n56762, n56763, n56764, n56765, n56766, n56767, n56768,
    n56769, n56770, n56771, n56772, n56773, n56774, n56775, n56776, n56777,
    n56778, n56779, n56780, n56781, n56782, n56784, n56785, n56786, n56787,
    n56788, n56789, n56790, n56791, n56792, n56793, n56794, n56795, n56796,
    n56797, n56798, n56799, n56800, n56801, n56802, n56803, n56804, n56805,
    n56806, n56807, n56808, n56809, n56810, n56811, n56812, n56813, n56814,
    n56815, n56816, n56817, n56818, n56819, n56820, n56821, n56822, n56823,
    n56824, n56825, n56826, n56827, n56828, n56829, n56830, n56832, n56833,
    n56834, n56835, n56836, n56837, n56838, n56839, n56840, n56841, n56842,
    n56843, n56844, n56845, n56846, n56847, n56848, n56849, n56850, n56851,
    n56852, n56853, n56854, n56855, n56856, n56857, n56858, n56859, n56860,
    n56861, n56862, n56863, n56864, n56865, n56866, n56867, n56868, n56869,
    n56870, n56871, n56872, n56873, n56874, n56875, n56876, n56877, n56878,
    n56880, n56881, n56882, n56883, n56884, n56885, n56886, n56887, n56888,
    n56889, n56890, n56891, n56892, n56893, n56894, n56895, n56896, n56897,
    n56898, n56899, n56900, n56901, n56902, n56903, n56904, n56905, n56906,
    n56907, n56908, n56909, n56910, n56911, n56912, n56913, n56914, n56915,
    n56916, n56917, n56918, n56919, n56920, n56921, n56922, n56923, n56924,
    n56925, n56926, n56928, n56929, n56930, n56931, n56932, n56933, n56934,
    n56935, n56936, n56937, n56938, n56939, n56940, n56941, n56942, n56943,
    n56944, n56945, n56946, n56947, n56948, n56949, n56950, n56951, n56952,
    n56953, n56954, n56955, n56956, n56957, n56958, n56959, n56960, n56961,
    n56962, n56963, n56964, n56965, n56966, n56967, n56968, n56969, n56970,
    n56971, n56972, n56973, n56974, n56976, n56977, n56978, n56979, n56980,
    n56981, n56982, n56983, n56984, n56985, n56986, n56987, n56988, n56989,
    n56990, n56991, n56992, n56993, n56994, n56995, n56996, n56997, n56998,
    n56999, n57000, n57001, n57002, n57003, n57004, n57005, n57006, n57007,
    n57008, n57009, n57010, n57011, n57012, n57013, n57014, n57015, n57016,
    n57017, n57018, n57019, n57020, n57021, n57022, n57024, n57025, n57026,
    n57027, n57028, n57029, n57030, n57031, n57032, n57033, n57034, n57035,
    n57036, n57037, n57038, n57039, n57040, n57041, n57042, n57043, n57044,
    n57045, n57046, n57047, n57048, n57049, n57050, n57051, n57052, n57053,
    n57054, n57055, n57056, n57057, n57058, n57059, n57060, n57061, n57062,
    n57063, n57064, n57065, n57066, n57067, n57068, n57069, n57070, n57072,
    n57073, n57074, n57075, n57076, n57077, n57078, n57079, n57080, n57081,
    n57082, n57083, n57084, n57085, n57086, n57087, n57088, n57089, n57090,
    n57091, n57092, n57093, n57094, n57095, n57096, n57097, n57098, n57099,
    n57100, n57101, n57102, n57103, n57104, n57105, n57106, n57107, n57108,
    n57109, n57110, n57111, n57112, n57113, n57114, n57115, n57116, n57117,
    n57118, n57120, n57121, n57122, n57123, n57124, n57125, n57126, n57127,
    n57129, n57130, n57131, n57132, n57133, n57134, n57135, n57136, n57138,
    n57139, n57140, n57141, n57142, n57143, n57144, n57146, n57147, n57148,
    n57149, n57150, n57151, n57152, n57153, n57155, n57156, n57157, n57158,
    n57159, n57160, n57161, n57162, n57163, n57165, n57166, n57167, n57168,
    n57169, n57170, n57171, n57172, n57174, n57175, n57176, n57177, n57178,
    n57179, n57180, n57181, n57182, n57184, n57185, n57186, n57187, n57188,
    n57189, n57190, n57191, n57193, n57194, n57195, n57196, n57197, n57198,
    n57199, n57200, n57201, n57203, n57204, n57205, n57206, n57207, n57208,
    n57209, n57210, n57212, n57213, n57214, n57215, n57216, n57217, n57218,
    n57219, n57220, n57222, n57223, n57224, n57225, n57226, n57227, n57228,
    n57229, n57231, n57232, n57233, n57234, n57235, n57236, n57237, n57238,
    n57239, n57241, n57242, n57243, n57244, n57245, n57246, n57247, n57248,
    n57250, n57251, n57252, n57253, n57254, n57255, n57256, n57257, n57258,
    n57260, n57261, n57262, n57263, n57264, n57265, n57266, n57267, n57269,
    n57270, n57271, n57272, n57273, n57274, n57275, n57276, n57277, n57279,
    n57280, n57281, n57282, n57283, n57284, n57285, n57286, n57288, n57289,
    n57290, n57291, n57292, n57293, n57294, n57295, n57296, n57298, n57299,
    n57300, n57301, n57302, n57303, n57304, n57305, n57307, n57308, n57309,
    n57310, n57311, n57312, n57313, n57314, n57315, n57317, n57318, n57319,
    n57320, n57321, n57322, n57323, n57324, n57326, n57327, n57328, n57329,
    n57330, n57331, n57332, n57333, n57334, n57336, n57337, n57338, n57339,
    n57340, n57341, n57342, n57343, n57345, n57346, n57347, n57348, n57349,
    n57350, n57351, n57352, n57353, n57355, n57356, n57357, n57358, n57359,
    n57360, n57361, n57362, n57364, n57365, n57366, n57367, n57368, n57369,
    n57370, n57371, n57372, n57374, n57375, n57376, n57377, n57378, n57379,
    n57380, n57381, n57383, n57384, n57385, n57386, n57387, n57388, n57389,
    n57390, n57391, n57393, n57394, n57395, n57396, n57397, n57398, n57399,
    n57400, n57402, n57403, n57404, n57405, n57406, n57407, n57408, n57409,
    n57410, n57412, n57413, n57414, n57415, n57416, n57417, n57418, n57419,
    n57421, n57422, n57423, n57424, n57425, n57426, n57428, n57429, n57430,
    n57431, n57432, n57433, n57434, n57435, n57436, n57437, n57438, n57439,
    n57440, n57441, n57442, n57443, n57444, n57445, n57446, n57447, n57448,
    n57449, n57450, n57451, n57452, n57453, n57454, n57455, n57456, n57457,
    n57458, n57459, n57460, n57461, n57462, n57463, n57464, n57465, n57466,
    n57467, n57468, n57469, n57471, n57472, n57473, n57474, n57475, n57476,
    n57477, n57478, n57479, n57480, n57481, n57482, n57483, n57484, n57485,
    n57486, n57487, n57488, n57489, n57490, n57491, n57492, n57494, n57495,
    n57496, n57497, n57498, n57499, n57500, n57501, n57502, n57503, n57504,
    n57505, n57506, n57507, n57508, n57509, n57510, n57511, n57512, n57513,
    n57514, n57515, n57516, n57517, n57518, n57519, n57520, n57521, n57522,
    n57524, n57525, n57526, n57527, n57528, n57529, n57530, n57531, n57532,
    n57533, n57534, n57535, n57536, n57537, n57538, n57539, n57540, n57541,
    n57542, n57543, n57544, n57545, n57546, n57547, n57548, n57549, n57550,
    n57551, n57552, n57553, n57555, n57556, n57557, n57558, n57559, n57560,
    n57561, n57562, n57563, n57564, n57565, n57566, n57567, n57568, n57569,
    n57570, n57571, n57572, n57573, n57574, n57575, n57576, n57577, n57578,
    n57579, n57580, n57581, n57582, n57583, n57584, n57585, n57586, n57587,
    n57588, n57589, n57590, n57592, n57593, n57594, n57595, n57596, n57597,
    n57598, n57599, n57600, n57601, n57602, n57603, n57604, n57605, n57606,
    n57607, n57608, n57609, n57610, n57611, n57612, n57613, n57614, n57615,
    n57616, n57617, n57618, n57619, n57620, n57621, n57623, n57624, n57625,
    n57626, n57627, n57628, n57629, n57630, n57631, n57632, n57633, n57634,
    n57635, n57636, n57637, n57638, n57639, n57640, n57641, n57642, n57643,
    n57644, n57645, n57646, n57647, n57648, n57649, n57651, n57652, n57653,
    n57654, n57655, n57656, n57657, n57658, n57659, n57660, n57661, n57662,
    n57663, n57664, n57665, n57666, n57667, n57668, n57669, n57670, n57671,
    n57672, n57673, n57674, n57675, n57677, n57678, n57679, n57680, n57681,
    n57682, n57683, n57684, n57685, n57686, n57687, n57688, n57689, n57690,
    n57691, n57692, n57693, n57694, n57695, n57696, n57697, n57698, n57699,
    n57700, n57701, n57702, n57703, n57705, n57706, n57707, n57708, n57709,
    n57710, n57711, n57712, n57713, n57714, n57715, n57716, n57717, n57718,
    n57719, n57720, n57721, n57722, n57723, n57724, n57725, n57726, n57727,
    n57728, n57729, n57731, n57732, n57733, n57734, n57735, n57736, n57737,
    n57738, n57739, n57740, n57741, n57742, n57743, n57744, n57745, n57746,
    n57747, n57748, n57749, n57750, n57751, n57752, n57753, n57754, n57755,
    n57756, n57757, n57759, n57760, n57761, n57762, n57763, n57764, n57765,
    n57766, n57767, n57768, n57769, n57770, n57771, n57772, n57773, n57774,
    n57775, n57776, n57777, n57778, n57779, n57780, n57781, n57782, n57783,
    n57785, n57786, n57787, n57788, n57789, n57790, n57791, n57792, n57793,
    n57794, n57795, n57796, n57797, n57798, n57799, n57800, n57801, n57802,
    n57803, n57804, n57805, n57806, n57807, n57808, n57809, n57810, n57811,
    n57813, n57814, n57815, n57816, n57817, n57818, n57819, n57820, n57821,
    n57822, n57823, n57824, n57825, n57826, n57827, n57828, n57829, n57830,
    n57831, n57832, n57833, n57834, n57835, n57836, n57837, n57839, n57840,
    n57841, n57842, n57843, n57844, n57845, n57846, n57847, n57848, n57849,
    n57850, n57851, n57852, n57853, n57854, n57855, n57856, n57857, n57858,
    n57859, n57860, n57861, n57862, n57863, n57864, n57865, n57867, n57868,
    n57869, n57870, n57871, n57872, n57873, n57874, n57875, n57876, n57877,
    n57878, n57879, n57880, n57881, n57882, n57883, n57884, n57885, n57886,
    n57887, n57888, n57889, n57890, n57891, n57893, n57894, n57895, n57896,
    n57897, n57898, n57899, n57900, n57901, n57902, n57903, n57904, n57905,
    n57906, n57907, n57908, n57909, n57910, n57911, n57912, n57913, n57914,
    n57915, n57916, n57917, n57918, n57919, n57921, n57922, n57923, n57924,
    n57925, n57926, n57927, n57928, n57929, n57930, n57931, n57932, n57933,
    n57934, n57935, n57936, n57937, n57938, n57939, n57940, n57941, n57942,
    n57943, n57944, n57945, n57947, n57948, n57949, n57950, n57951, n57952,
    n57953, n57954, n57955, n57956, n57957, n57958, n57959, n57960, n57961,
    n57962, n57963, n57964, n57965, n57966, n57967, n57968, n57969, n57970,
    n57971, n57972, n57973, n57975, n57976, n57977, n57978, n57979, n57980,
    n57981, n57982, n57983, n57984, n57985, n57986, n57987, n57988, n57989,
    n57990, n57991, n57992, n57993, n57994, n57995, n57996, n57997, n57998,
    n57999, n58001, n58002, n58003, n58004, n58005, n58006, n58007, n58008,
    n58009, n58010, n58011, n58012, n58013, n58014, n58015, n58016, n58017,
    n58018, n58019, n58020, n58021, n58022, n58023, n58024, n58025, n58026,
    n58028, n58029, n58030, n58031, n58032, n58033, n58034, n58035, n58036,
    n58037, n58038, n58039, n58040, n58041, n58042, n58043, n58044, n58045,
    n58046, n58047, n58048, n58049, n58050, n58051, n58053, n58054, n58055,
    n58056, n58057, n58058, n58059, n58060, n58061, n58062, n58063, n58064,
    n58065, n58066, n58067, n58068, n58069, n58070, n58071, n58072, n58073,
    n58074, n58075, n58076, n58077, n58078, n58080, n58081, n58082, n58083,
    n58084, n58085, n58086, n58087, n58088, n58089, n58090, n58091, n58092,
    n58093, n58094, n58095, n58096, n58097, n58098, n58099, n58100, n58101,
    n58102, n58103, n58105, n58106, n58107, n58108, n58109, n58110, n58111,
    n58112, n58113, n58114, n58115, n58116, n58117, n58118, n58119, n58120,
    n58121, n58122, n58123, n58124, n58125, n58126, n58127, n58128, n58129,
    n58130, n58132, n58133, n58134, n58135, n58136, n58137, n58138, n58139,
    n58140, n58141, n58142, n58143, n58144, n58145, n58146, n58147, n58148,
    n58149, n58150, n58151, n58152, n58153, n58154, n58155, n58157, n58158,
    n58159, n58160, n58161, n58162, n58163, n58164, n58165, n58166, n58167,
    n58168, n58169, n58170, n58171, n58172, n58173, n58174, n58175, n58176,
    n58177, n58178, n58179, n58180, n58181, n58182, n58184, n58185, n58186,
    n58187, n58188, n58189, n58190, n58191, n58192, n58193, n58194, n58195,
    n58196, n58197, n58198, n58199, n58200, n58201, n58202, n58203, n58204,
    n58205, n58206, n58207, n58209, n58210, n58211, n58212, n58213, n58214,
    n58215, n58216, n58217, n58218, n58219, n58220, n58221, n58222, n58223,
    n58224, n58225, n58226, n58227, n58228, n58229, n58230, n58231, n58232,
    n58233, n58234, n58236, n58237, n58238, n58239, n58240, n58241, n58242,
    n58243, n58244, n58245, n58246, n58247, n58248, n58249, n58250, n58251,
    n58252, n58253, n58254, n58255, n58256, n58257, n58258, n58259, n58261,
    n58262, n58263, n58264, n58265, n58266, n58267, n58268, n58269, n58270,
    n58271, n58272, n58273, n58274, n58275, n58276, n58277, n58278, n58279,
    n58280, n58281, n58282, n58283, n58284, n58286, n58287, n58288, n58289,
    n58290, n58291, n58292, n58293, n58294, n58295, n58296, n58297, n58298,
    n58299, n58300, n58301, n58302, n58303, n58304, n58305, n58306, n58307,
    n58308, n58309, n58311, n58312, n58313, n58314, n58315, n58316, n58317,
    n58318, n58319, n58320, n58321, n58322, n58323, n58324, n58325, n58326,
    n58327, n58328, n58329, n58330, n58331, n58332, n58333, n58334, n58335,
    n58336, n58337, n58338, n58339, n58340, n58341, n58342, n58343, n58344,
    n58345, n58346, n58347, n58348, n58350, n58351, n58352, n58353, n58354,
    n58355, n58356, n58357, n58359, n58360, n58361, n58363, n58364, n58365,
    n58367, n58368, n58370, n58371, n58372, n58374, n58375, n58377, n58378,
    n58379, n58380, n58382, n58383, n58384, n58385, n58386, n58387, n58388,
    n58389, n58390, n58391, n58392, n58393, n58394, n58395, n58396, n58398,
    n58399, n58400, n58402, n58403, n58405, n58406, n58407, n58409, n58411,
    n58412, n58413, n58414, n58415, n58417, n58418, n58419, n58421, n58422,
    n58423, n58425, n58426, n58428, n58429, n58431, n58432, n58434, n58435,
    n58436, n58437, n58438, n58439, n58441, n58442, n58443, n58444, n58446,
    n58447, n58448, n58449, n58451, n58452, n58453, n58454, n58456, n58457,
    n58458, n58459, n58461, n58462, n58463, n58464, n58466, n58467, n58468,
    n58469, n58471, n58472, n58473, n58474, n58476, n58477, n58478, n58479,
    n58481, n58482, n58483, n58484, n58486, n58487, n58488, n58489, n58491,
    n58492, n58493, n58494, n58496, n58497, n58498, n58499, n58501, n58502,
    n58503, n58504, n58506, n58507, n58508, n58509, n58511, n58512, n58513,
    n58514, n58516, n58517, n58518, n58519, n58521, n58522, n58523, n58524,
    n58526, n58527, n58528, n58529, n58531, n58532, n58533, n58534, n58536,
    n58537, n58538, n58539, n58541, n58542, n58543, n58544, n58546, n58547,
    n58548, n58549, n58551, n58552, n58553, n58554, n58556, n58557, n58558,
    n58559, n58561, n58562, n58563, n58564, n58566, n58567, n58568, n58569,
    n58571, n58572, n58573, n58574, n58576, n58577, n58578, n58579, n58581,
    n58582, n58583, n58584, n58586, n58587, n58588, n58589, n58590, n58591,
    n58592, n58593, n58594, n58595, n58596, n58597, n58598, n58599, n58600,
    n58601, n58602, n58603, n58604, n58605, n58606, n58607, n58608, n58609,
    n58610, n58611, n58612, n58613, n58615, n58616, n58617, n58618, n58619,
    n58620, n58621, n58622, n58623, n58624, n58625, n58626, n58627, n58629,
    n58630, n58631, n58632, n58633, n58634, n58635, n58636, n58637, n58639,
    n58640, n58641, n58642, n58643, n58644, n58646, n58647, n58679, n58680,
    n58681, n58682, n58683, n58684, n58685, n58686, n58687, n58688, n58689,
    n58690, n58691, n58692, n58693, n58694, n58695, n58696, n58697, n58698,
    n58699, n58700, n58701, n58702, n58703, n58704, n58705, n58706, n58707,
    n58708, n58709, n58710, n58711, n58712, n58713, n58714, n58715, n58716,
    n58717, n58718, n58719, n58720, n58721, n58722, n58723, n58724, n58725,
    n58726, n58727, n58728, n58729, n58730, n58731, n58732, n58733, n58734,
    n58735, n58736, n58737, n58738, n58739, n58740, n58741, n58742, n58743,
    n58744, n58745, n58746, n58747, n58748, n58749, n58750, n58751, n58752,
    n58753, n58754, n58755, n58756, n58757, n58758, n58759, n58760, n58761,
    n58762, n58763, n58764, n58765, n58766, n58767, n58768, n58769, n58770,
    n58771, n58772, n58773, n58774, n58775, n58776, n58777, n58778, n58779,
    n58780, n58781, n58782, n58783, n58784, n58785, n58786, n58787, n58788,
    n58789, n58790, n58791, n58792, n58793, n58794, n58795, n58796, n58797,
    n58798, n58799, n58800, n58801, n58802, n58803, n58804, n58805, n58806,
    n58807, n58808, n58809, n58810, n58811, n58812, n58813, n58814, n58815,
    n58816, n58817, n58818, n58819, n58820, n58821, n58822, n58823, n58824,
    n58825, n58826, n58827, n58828, n58829, n58830, n58831, n58832, n58833,
    n58834, n58835, n58836, n58837, n58838, n58839, n58840, n58841, n58842,
    n58843, n58844, n58845, n58846, n58847, n58848, n58849, n58850, n58851,
    n58852, n58853, n58854, n58855, n58856, n58857, n58858, n58859, n58860,
    n58861, n58862, n58863, n58864, n58865, n58866, n58867, n58868, n58869,
    n58870, n58871, n58872, n58873, n58874, n58875, n58876, n58877, n58878,
    n58879, n58880, n58881, n58882, n58883, n58884, n58885, n58886, n58887,
    n58888, n58889, n58890, n58891, n58892, n58893, n58894, n58895, n58896,
    n58897, n58898, n58899, n58900, n58901, n58902, n58903, n58904, n58905,
    n58906, n58907, n58908, n58909, n58910, n58911, n58912, n58913, n58914,
    n58915, n58916, n58917, n58918, n58919, n58920, n58921, n58922, n58923,
    n58924, n58925, n58926, n58927, n58928, n58929, n58930, n58931, n58932,
    n58933, n58934, n58935, n58936, n58937, n58938, n58939, n58940, n58941,
    n58942, n58943, n58944, n58945, n58946, n58947, n58948, n58949, n58950,
    n58951, n58952, n58953, n58954, n58955, n58956, n58957, n58958, n58959,
    n58960, n58961, n58962, n58963, n58964, n58965, n58966, n58967, n58968,
    n58969, n58970, n58971, n58972, n58973, n58974, n58975, n58976, n58977,
    n58978, n58979, n58980, n58981, n58982, n58983, n58984, n58985, n58986,
    n58987, n58988, n58989, n58990, n58991, n58992, n58993, n58994, n58995,
    n58996, n58997, n58998, n58999, n59000, n59001, n59002, n59003, n59004,
    n59005, n59006, n59007, n59008, n59009, n59010, n59011, n59012, n59013,
    n59014, n59015, n59016, n59017, n59018, n59019, n59020, n59021, n59022,
    n59023, n59024, n59025, n59026, n59027, n59028, n59029, n59030, n59031,
    n59032, n59033, n59034, n59035, n59036, n59037, n59038, n59039, n59040,
    n59041, n59042, n59043, n59044, n59045, n59046, n59047, n59048, n59049,
    n59050, n59051, n59052, n59053, n59054, n59055, n59056, n59057, n59058,
    n59059, n59060, n59061, n59062, n59063, n59064, n59065, n59066, n59067,
    n59068, n59069, n59070, n59071, n59072, n59073, n59074, n59075, n59076,
    n59077, n59078, n59079, n59080, n59081, n59082, n59083, n59084, n59085,
    n59086, n59087, n59088, n59089, n59090, n59091, n59092, n59093, n59094,
    n59095, n59096, n59097, n59098, n59099, n59100, n59101, n59102, n59103,
    n59104, n59105, n59106, n59107, n59108, n59109, n59110, n59111, n59112,
    n59113, n59114, n59115, n59116, n59117, n59118, n59119, n59120, n59121,
    n59122, n59123, n59124, n59125, n59126, n59127, n59128, n59129, n59130,
    n59131, n59132, n59133, n59134, n59135, n59136, n59137, n59138, n59139,
    n59140, n59141, n59142, n59143, n59144, n59145, n59146, n59147, n59148,
    n59149, n59150, n59151, n59152, n59153, n59154, n59155, n59156, n59157,
    n59158, n59159, n59160, n59161, n59162, n59163, n59164, n59165, n59166,
    n59167, n59168, n59169, n59170, n59171, n59172, n59173, n59174, n59175,
    n59176, n59177, n59178, n59179, n59180, n59181, n59182, n59183, n59184,
    n59185, n59186, n59187, n59188, n59189, n59190, n59191, n59192, n59193,
    n59194, n59195, n59196, n59197, n59198, n59199, n59200, n59201, n59202,
    n59203, n59204, n59205, n59206, n59207, n59208, n59209, n59210, n59211,
    n59212, n59213, n59214, n59215, n59216, n59217, n59218, n59219, n59220,
    n59221, n59222, n59223, n59224, n59225, n59226, n59227, n59228, n59229,
    n59230, n59231, n59232, n59233, n59234, n59235, n59236, n59237, n59238,
    n59239, n59240, n59241, n59242, n59243, n59244, n59245, n59246, n59247,
    n59248, n59249, n59250, n59251, n59252, n59253, n59254, n59255, n59256,
    n59257, n59258, n59259, n59260, n59261, n59262, n59263, n59264, n59265,
    n59266, n59267, n59268, n59269, n59270, n59271, n59272, n59273, n59274,
    n59275, n59276, n59277, n59278, n59279, n59280, n59281, n59282, n59283,
    n59284, n59285, n59286, n59287, n59288, n59289, n59290, n59291, n59292,
    n59293, n59294, n59295, n59296, n59297, n59298, n59299, n59300, n59301,
    n59302, n59303, n59304, n59305, n59306, n59307, n59308, n59309, n59310,
    n59312, n59313, n59314, n59315, n59316, n59317, n59318, n59319, n59321,
    n59322, n59323, n59324, n59325, n59326, n59327, n59328, n59329, n59330,
    n59331, n59332, n59333, n59334, n59336, n59337, n59338, n59339, n59340,
    n59341, n59342, n59343, n59344, n59345, n59346, n59347, n59348, n59349,
    n59350, n59351, n59352, n59353, n59354, n59355, n59356, n59357, n59358,
    n59359, n59360, n59361, n59362, n59363, n59364, n59365, n59366, n59367,
    n59368, n59369, n59370, n59371, n59372, n59373, n59374, n59375, n59377,
    n59378, n59379, n59380, n59381, n59382, n59383, n59384, n59385, n59386,
    n59387, n59388, n59389, n59390, n59391, n59392, n59393, n59394, n59395,
    n59396, n59397, n59398, n59399, n59400, n59401, n59402, n59403, n59404,
    n59405, n59406, n59407, n59408, n59409, n59410, n59411, n59412, n59413,
    n59414, n59415, n59416, n59417, n59418, n59419, n59420, n59421, n59422,
    n59423, n59424, n59425, n59426, n59427, n59428, n59429, n59430, n59431,
    n59432, n59433, n59434, n59435, n59436, n59437, n59438, n59439, n59440,
    n59441, n59442, n59443, n59444, n59445, n59446, n59447, n59448, n59449,
    n59450, n59451, n59452, n59454, n59455, n59456, n59457, n59458, n59459,
    n59460, n59461, n59462, n59463, n59464, n59465, n59467, n59468, n59469,
    n59470, n59471, n59472, n59473, n59474, n59475, n59476, n59477, n59478,
    n59480, n59481, n59482, n59483, n59484, n59485, n59486, n59487, n59488,
    n59489, n59490, n59491, n59493, n59494, n59495, n59496, n59497, n59498,
    n59499, n59500, n59501, n59502, n59503, n59504, n59506, n59507, n59508,
    n59509, n59510, n59511, n59512, n59513, n59514, n59515, n59516, n59517,
    n59519, n59520, n59521, n59522, n59523, n59524, n59525, n59526, n59527,
    n59528, n59529, n59530, n59532, n59533, n59534, n59535, n59536, n59537,
    n59538, n59539, n59540, n59541, n59542, n59543, n59545, n59546, n59547,
    n59548, n59549, n59550, n59551, n59552, n59553, n59554, n59555, n59556,
    n59557, n59558, n59559, n59560, n59561, n59562, n59563, n59564, n59565,
    n59566, n59567, n59568, n59569, n59571, n59572, n59573, n59574, n59575,
    n59576, n59577, n59578, n59580, n59581, n59582, n59583, n59584, n59585,
    n59586, n59587, n59589, n59590, n59591, n59592, n59593, n59594, n59595,
    n59596, n59598, n59599, n59600, n59601, n59602, n59603, n59604, n59605,
    n59607, n59608, n59609, n59610, n59611, n59612, n59613, n59614, n59616,
    n59617, n59618, n59619, n59620, n59621, n59622, n59623, n59625, n59626,
    n59627, n59628, n59629, n59630, n59631, n59632, n59634, n59635, n59636,
    n59637, n59638, n59639, n59640, n59641, n59642, n59643, n59644, n59645,
    n59646, n59647, n59648, n59649, n59650, n59651, n59652, n59653, n59654,
    n59655, n59656, n59657, n59659, n59660, n59661, n59662, n59663, n59664,
    n59665, n59666, n59668, n59669, n59670, n59671, n59672, n59673, n59674,
    n59675, n59677, n59678, n59679, n59680, n59681, n59682, n59683, n59684,
    n59686, n59687, n59688, n59689, n59690, n59691, n59692, n59693, n59695,
    n59696, n59697, n59698, n59699, n59700, n59701, n59702, n59704, n59705,
    n59706, n59707, n59708, n59709, n59710, n59711, n59713, n59714, n59715,
    n59716, n59717, n59718, n59719, n59720, n59722, n59723, n59724, n59725,
    n59726, n59727, n59728, n59729, n59730, n59731, n59732, n59733, n59734,
    n59735, n59736, n59737, n59738, n59739, n59740, n59741, n59742, n59743,
    n59744, n59745, n59747, n59748, n59749, n59750, n59751, n59752, n59753,
    n59754, n59756, n59757, n59758, n59759, n59760, n59761, n59762, n59763,
    n59765, n59766, n59767, n59768, n59769, n59770, n59771, n59772, n59774,
    n59775, n59776, n59777, n59778, n59779, n59780, n59781, n59783, n59784,
    n59785, n59786, n59787, n59788, n59789, n59790, n59792, n59793, n59794,
    n59795, n59796, n59797, n59798, n59799, n59801, n59802, n59803, n59804,
    n59805, n59806, n59807, n59808, n59810, n59811, n59812, n59813, n59814,
    n59815, n59816, n59817, n59818, n59819, n59820, n59821, n59822, n59823,
    n59824, n59825, n59826, n59827, n59828, n59829, n59830, n59831, n59832,
    n59833, n59834, n59836, n59837, n59838, n59839, n59840, n59841, n59842,
    n59843, n59845, n59846, n59847, n59848, n59849, n59850, n59851, n59852,
    n59854, n59855, n59856, n59857, n59858, n59859, n59860, n59861, n59863,
    n59864, n59865, n59866, n59867, n59868, n59869, n59870, n59872, n59873,
    n59874, n59875, n59876, n59877, n59878, n59879, n59881, n59882, n59883,
    n59884, n59885, n59886, n59887, n59888, n59890, n59891, n59892, n59893,
    n59894, n59895, n59896, n59897, n59899, n59900, n59901, n59902, n59903,
    n59904, n59905, n59906, n59907, n59908, n59909, n59910, n59911, n59912,
    n59913, n59914, n59915, n59916, n59917, n59918, n59919, n59920, n59921,
    n59923, n59924, n59925, n59926, n59927, n59928, n59929, n59930, n59932,
    n59933, n59934, n59935, n59936, n59937, n59938, n59939, n59941, n59942,
    n59943, n59944, n59945, n59946, n59947, n59948, n59950, n59951, n59952,
    n59953, n59954, n59955, n59956, n59957, n59959, n59960, n59961, n59962,
    n59963, n59964, n59965, n59966, n59968, n59969, n59970, n59971, n59972,
    n59973, n59974, n59975, n59977, n59978, n59979, n59980, n59981, n59982,
    n59983, n59984, n59986, n59987, n59988, n59989, n59990, n59991, n59992,
    n59993, n59994, n59995, n59996, n59997, n59998, n59999, n60000, n60001,
    n60002, n60003, n60004, n60005, n60006, n60007, n60009, n60010, n60011,
    n60012, n60013, n60014, n60015, n60016, n60018, n60019, n60020, n60021,
    n60022, n60023, n60024, n60025, n60027, n60028, n60029, n60030, n60031,
    n60032, n60033, n60034, n60036, n60037, n60038, n60039, n60040, n60041,
    n60042, n60043, n60045, n60046, n60047, n60048, n60049, n60050, n60051,
    n60052, n60054, n60055, n60056, n60057, n60058, n60059, n60060, n60061,
    n60063, n60064, n60065, n60066, n60067, n60068, n60069, n60070, n60072,
    n60073, n60074, n60075, n60076, n60077, n60078, n60079, n60080, n60081,
    n60082, n60083, n60084, n60085, n60086, n60087, n60088, n60089, n60090,
    n60091, n60092, n60094, n60095, n60096, n60097, n60098, n60099, n60100,
    n60101, n60103, n60104, n60105, n60106, n60107, n60108, n60109, n60110,
    n60112, n60113, n60114, n60115, n60116, n60117, n60118, n60119, n60121,
    n60122, n60123, n60124, n60125, n60126, n60127, n60128, n60130, n60131,
    n60132, n60133, n60134, n60135, n60136, n60137, n60139, n60140, n60141,
    n60142, n60143, n60144, n60145, n60146, n60148, n60149, n60150, n60151,
    n60152, n60153, n60154, n60155, n60157, n60158, n60159, n60160, n60161,
    n60162, n60163, n60164, n60165, n60166, n60167, n60168, n60169, n60170,
    n60171, n60172, n60173, n60174, n60175, n60176, n60178, n60179, n60180,
    n60181, n60182, n60183, n60184, n60185, n60187, n60188, n60189, n60190,
    n60191, n60192, n60193, n60194, n60196, n60197, n60198, n60199, n60200,
    n60201, n60202, n60203, n60205, n60206, n60207, n60208, n60209, n60210,
    n60211, n60212, n60214, n60215, n60216, n60217, n60218, n60219, n60220,
    n60221, n60223, n60224, n60225, n60226, n60227, n60228, n60229, n60230,
    n60232, n60233, n60234, n60235, n60236, n60237, n60238, n60239, n60241,
    n60242, n60243, n60244, n60245, n60246, n60247, n60248, n60249, n60250,
    n60251, n60252, n60253, n60254, n60255, n60256, n60257, n60258, n60259,
    n60260, n60261, n60262, n60263, n60265, n60266, n60267, n60268, n60269,
    n60270, n60271, n60272, n60274, n60275, n60276, n60277, n60278, n60279,
    n60280, n60281, n60283, n60284, n60285, n60286, n60287, n60288, n60289,
    n60290, n60292, n60293, n60294, n60295, n60296, n60297, n60298, n60299,
    n60301, n60302, n60303, n60304, n60305, n60306, n60307, n60308, n60310,
    n60311, n60312, n60313, n60314, n60315, n60316, n60317, n60319, n60320,
    n60321, n60322, n60323, n60324, n60325, n60326, n60328, n60329, n60330,
    n60331, n60332, n60333, n60334, n60335, n60336, n60337, n60338, n60339,
    n60340, n60341, n60342, n60343, n60344, n60345, n60346, n60347, n60348,
    n60349, n60350, n60352, n60353, n60354, n60355, n60356, n60357, n60358,
    n60359, n60361, n60362, n60363, n60364, n60365, n60366, n60367, n60368,
    n60370, n60371, n60372, n60373, n60374, n60375, n60376, n60377, n60379,
    n60380, n60381, n60382, n60383, n60384, n60385, n60386, n60388, n60389,
    n60390, n60391, n60392, n60393, n60394, n60395, n60397, n60398, n60399,
    n60400, n60401, n60402, n60403, n60404, n60406, n60407, n60408, n60409,
    n60410, n60411, n60412, n60413, n60415, n60416, n60417, n60418, n60419,
    n60420, n60421, n60422, n60423, n60424, n60425, n60426, n60427, n60428,
    n60429, n60430, n60431, n60432, n60433, n60434, n60435, n60437, n60438,
    n60439, n60440, n60441, n60442, n60443, n60444, n60446, n60447, n60448,
    n60449, n60450, n60451, n60452, n60453, n60455, n60456, n60457, n60458,
    n60459, n60460, n60461, n60462, n60464, n60465, n60466, n60467, n60468,
    n60469, n60470, n60471, n60473, n60474, n60475, n60476, n60477, n60478,
    n60479, n60480, n60482, n60483, n60484, n60485, n60486, n60487, n60488,
    n60489, n60491, n60492, n60493, n60494, n60495, n60496, n60497, n60498,
    n60500, n60501, n60502, n60503, n60504, n60505, n60506, n60507, n60508,
    n60509, n60510, n60511, n60512, n60513, n60514, n60515, n60516, n60517,
    n60518, n60519, n60520, n60521, n60522, n60523, n60525, n60526, n60527,
    n60528, n60529, n60530, n60531, n60532, n60534, n60535, n60536, n60537,
    n60538, n60539, n60540, n60541, n60543, n60544, n60545, n60546, n60547,
    n60548, n60549, n60550, n60552, n60553, n60554, n60555, n60556, n60557,
    n60558, n60559, n60561, n60562, n60563, n60564, n60565, n60566, n60567,
    n60568, n60570, n60571, n60572, n60573, n60574, n60575, n60576, n60577,
    n60579, n60580, n60581, n60582, n60583, n60584, n60585, n60586, n60588,
    n60589, n60590, n60591, n60592, n60593, n60594, n60595, n60596, n60597,
    n60598, n60599, n60600, n60601, n60602, n60603, n60604, n60605, n60606,
    n60607, n60609, n60610, n60611, n60612, n60613, n60614, n60615, n60616,
    n60618, n60619, n60620, n60621, n60622, n60623, n60624, n60625, n60627,
    n60628, n60629, n60630, n60631, n60632, n60633, n60634, n60636, n60637,
    n60638, n60639, n60640, n60641, n60642, n60643, n60645, n60646, n60647,
    n60648, n60649, n60650, n60651, n60652, n60654, n60655, n60656, n60657,
    n60658, n60659, n60660, n60661, n60663, n60664, n60665, n60666, n60667,
    n60668, n60669, n60670, n60672, n60673, n60674, n60675, n60676, n60677,
    n60678, n60679, n60680, n60681, n60682, n60683, n60684, n60685, n60686,
    n60687, n60688, n60689, n60690, n60691, n60693, n60694, n60695, n60696,
    n60697, n60698, n60699, n60700, n60702, n60703, n60704, n60705, n60706,
    n60707, n60708, n60709, n60711, n60712, n60713, n60714, n60715, n60716,
    n60717, n60718, n60720, n60721, n60722, n60723, n60724, n60725, n60726,
    n60727, n60729, n60730, n60731, n60732, n60733, n60734, n60735, n60736,
    n60738, n60739, n60740, n60741, n60742, n60743, n60744, n60745, n60747,
    n60748, n60749, n60750, n60751, n60752, n60753, n60754, n60756, n60757,
    n60758, n60759, n60760, n60761, n60762, n60763, n60764, n60765, n60766,
    n60767, n60768, n60769, n60770, n60771, n60772, n60773, n60774, n60776,
    n60777, n60778, n60779, n60780, n60781, n60782, n60783, n60785, n60786,
    n60787, n60788, n60789, n60790, n60791, n60792, n60794, n60795, n60796,
    n60797, n60798, n60799, n60800, n60801, n60803, n60804, n60805, n60806,
    n60807, n60808, n60809, n60810, n60812, n60813, n60814, n60815, n60816,
    n60817, n60818, n60819, n60821, n60822, n60823, n60824, n60825, n60826,
    n60827, n60828, n60830, n60831, n60832, n60833, n60834, n60835, n60836,
    n60837, n60839, n60840, n60841, n60842, n60843, n60844, n60845, n60846,
    n60847, n60848, n60850, n60851, n60852, n60853, n60854, n60855, n60857,
    n60858, n60859, n60860, n60861, n60862, n60863, n60864, n60866, n60867,
    n60868, n60869, n60870, n60871, n60872, n60874, n60875, n60876, n60877,
    n60878, n60879, n60880, n60882, n60883, n60884, n60885, n60887, n60888,
    n60889, n60890, n60891, n60892, n60893, n60894, n60895, n60896, n60897,
    n60898, n60899, n60901, n60902, n60903, n60904, n60905, n60906, n60907,
    n60908, n60909, n60910, n60911, n60912, n60913, n60915, n60916, n60917,
    n60918, n60919, n60920, n60921, n60922, n60923, n60924, n60925, n60926,
    n60928, n60929, n60930, n60931, n60932, n60934, n60935, n60936, n60937,
    n60938, n60939, n60940, n60941, n60942, n60943, n60944, n60945, n60946,
    n60947, n60948, n60949, n60950, n60951, n60952, n60953, n60954, n60955,
    n60956, n60957, n60958, n60959, n60960, n60961, n60962, n60963, n60964,
    n60965, n60966, n60967, n60968, n60969, n60970, n60971, n60972, n60973,
    n60974, n60975, n60976, n60977, n60978, n60979, n60980, n60981, n60982,
    n60983, n60984, n60985, n60986, n60987, n60988, n60989, n60990, n60991,
    n60992, n60993, n60994, n60995, n60996, n60997, n60998, n60999, n61000,
    n61001, n61002, n61003, n61004, n61005, n61006, n61007, n61008, n61009,
    n61010, n61011, n61012, n61013, n61014, n61015, n61016, n61017, n61018,
    n61019, n61020, n61021, n61022, n61023, n61024, n61025, n61026, n61027,
    n61028, n61029, n61030, n61031, n61032, n61033, n61034, n61035, n61036,
    n61037, n61038, n61039, n61040, n61041, n61042, n61043, n61044, n61045,
    n61046, n61047, n61048, n61049, n61050, n61051, n61052, n61053, n61054,
    n61055, n61056, n61057, n61058, n61059, n61060, n61061, n61062, n61063,
    n61064, n61065, n61066, n61067, n61068, n61069, n61070, n61071, n61072,
    n61073, n61074, n61075, n61076, n61077, n61078, n61079, n61080, n61081,
    n61082, n61083, n61084, n61085, n61086, n61087, n61088, n61089, n61090,
    n61091, n61092, n61093, n61094, n61095, n61096, n61097, n61098, n61099,
    n61100, n61101, n61102, n61103, n61104, n61105, n61106, n61107, n61108,
    n61110, n61111, n61112, n61113, n61114, n61115, n61116, n61117, n61118,
    n61119, n61120, n61121, n61122, n61123, n61124, n61125, n61126, n61127,
    n61128, n61129, n61130, n61131, n61132, n61133, n61134, n61135, n61136,
    n61137, n61138, n61139, n61140, n61141, n61142, n61143, n61144, n61145,
    n61146, n61147, n61148, n61149, n61150, n61151, n61152, n61153, n61154,
    n61155, n61156, n61157, n61158, n61159, n61160, n61161, n61162, n61163,
    n61164, n61165, n61166, n61167, n61168, n61169, n61170, n61171, n61172,
    n61173, n61174, n61175, n61176, n61177, n61178, n61179, n61180, n61181,
    n61182, n61183, n61184, n61185, n61186, n61187, n61188, n61189, n61190,
    n61191, n61192, n61193, n61194, n61195, n61196, n61197, n61198, n61199,
    n61200, n61201, n61202, n61203, n61204, n61205, n61206, n61207, n61208,
    n61209, n61210, n61211, n61212, n61213, n61214, n61215, n61216, n61218,
    n61219, n61220, n61221, n61222, n61223, n61224, n61225, n61226, n61227,
    n61228, n61229, n61230, n61231, n61232, n61233, n61234, n61235, n61236,
    n61237, n61238, n61239, n61240, n61241, n61242, n61243, n61244, n61245,
    n61246, n61247, n61248, n61249, n61250, n61251, n61252, n61253, n61254,
    n61255, n61256, n61257, n61258, n61259, n61260, n61261, n61262, n61263,
    n61264, n61265, n61266, n61267, n61268, n61269, n61270, n61271, n61272,
    n61273, n61274, n61275, n61276, n61277, n61278, n61279, n61280, n61281,
    n61282, n61283, n61284, n61285, n61286, n61287, n61288, n61289, n61290,
    n61291, n61292, n61293, n61294, n61295, n61296, n61297, n61298, n61299,
    n61300, n61301, n61302, n61303, n61304, n61305, n61306, n61307, n61308,
    n61309, n61310, n61311, n61312, n61313, n61314, n61315, n61316, n61317,
    n61318, n61319, n61320, n61321, n61322, n61323, n61324, n61325, n61326,
    n61327, n61328, n61329, n61330, n61331, n61332, n61333, n61334, n61335,
    n61336, n61337, n61339, n61340, n61341, n61342, n61343, n61344, n61345,
    n61346, n61347, n61348, n61349, n61350, n61351, n61352, n61353, n61354,
    n61355, n61356, n61357, n61358, n61359, n61360, n61361, n61362, n61363,
    n61364, n61365, n61366, n61367, n61368, n61369, n61370, n61371, n61372,
    n61373, n61374, n61375, n61376, n61377, n61378, n61379, n61380, n61381,
    n61382, n61383, n61384, n61385, n61386, n61387, n61388, n61389, n61390,
    n61391, n61392, n61393, n61394, n61395, n61396, n61397, n61398, n61399,
    n61400, n61401, n61402, n61403, n61404, n61405, n61406, n61407, n61408,
    n61409, n61410, n61411, n61412, n61413, n61414, n61415, n61416, n61417,
    n61418, n61419, n61420, n61421, n61422, n61423, n61424, n61425, n61426,
    n61427, n61428, n61429, n61430, n61431, n61432, n61433, n61434, n61435,
    n61436, n61437, n61438, n61439, n61440, n61441, n61442, n61443, n61444,
    n61445, n61446, n61447, n61448, n61449, n61450, n61451, n61452, n61453,
    n61454, n61455, n61456, n61457, n61458, n61459, n61460, n61461, n61462,
    n61463, n61464, n61465, n61466, n61467, n61468, n61470, n61471, n61472,
    n61473, n61474, n61475, n61476, n61477, n61478, n61479, n61480, n61481,
    n61482, n61483, n61484, n61485, n61486, n61487, n61488, n61489, n61490,
    n61491, n61492, n61493, n61494, n61495, n61496, n61497, n61498, n61499,
    n61500, n61501, n61502, n61503, n61504, n61505, n61506, n61507, n61508,
    n61509, n61510, n61511, n61512, n61513, n61514, n61515, n61516, n61517,
    n61518, n61519, n61520, n61521, n61522, n61523, n61524, n61525, n61526,
    n61527, n61528, n61529, n61530, n61531, n61532, n61533, n61534, n61535,
    n61536, n61537, n61538, n61539, n61540, n61541, n61542, n61543, n61544,
    n61545, n61546, n61547, n61548, n61549, n61550, n61551, n61552, n61553,
    n61554, n61555, n61556, n61557, n61558, n61559, n61560, n61561, n61562,
    n61563, n61564, n61565, n61566, n61567, n61568, n61569, n61570, n61571,
    n61572, n61573, n61574, n61575, n61576, n61577, n61578, n61579, n61580,
    n61581, n61582, n61583, n61584, n61585, n61586, n61587, n61588, n61589,
    n61590, n61591, n61592, n61593, n61594, n61595, n61596, n61597, n61598,
    n61599, n61600, n61601, n61602, n61603, n61604, n61606, n61607, n61608,
    n61609, n61610, n61611, n61612, n61613, n61614, n61615, n61616, n61617,
    n61618, n61619, n61620, n61621, n61622, n61623, n61624, n61625, n61626,
    n61627, n61628, n61629, n61630, n61631, n61632, n61633, n61634, n61635,
    n61636, n61637, n61638, n61639, n61640, n61641, n61642, n61643, n61644,
    n61645, n61646, n61647, n61648, n61649, n61650, n61651, n61652, n61653,
    n61654, n61655, n61656, n61657, n61658, n61659, n61660, n61661, n61662,
    n61663, n61664, n61665, n61666, n61667, n61668, n61669, n61670, n61671,
    n61672, n61673, n61674, n61675, n61676, n61677, n61678, n61679, n61680,
    n61681, n61682, n61683, n61684, n61685, n61686, n61687, n61688, n61689,
    n61690, n61691, n61692, n61693, n61694, n61695, n61696, n61697, n61698,
    n61699, n61700, n61701, n61702, n61703, n61704, n61705, n61706, n61707,
    n61708, n61709, n61710, n61711, n61712, n61713, n61714, n61715, n61716,
    n61717, n61718, n61719, n61720, n61721, n61722, n61723, n61724, n61725,
    n61726, n61727, n61728, n61729, n61730, n61731, n61732, n61733, n61734,
    n61735, n61736, n61737, n61739, n61740, n61741, n61742, n61743, n61744,
    n61745, n61746, n61747, n61748, n61749, n61750, n61751, n61752, n61753,
    n61754, n61755, n61756, n61757, n61758, n61759, n61760, n61761, n61762,
    n61763, n61764, n61765, n61766, n61767, n61768, n61769, n61770, n61771,
    n61772, n61773, n61774, n61775, n61776, n61777, n61778, n61779, n61780,
    n61781, n61782, n61783, n61784, n61785, n61786, n61787, n61788, n61789,
    n61790, n61791, n61792, n61793, n61794, n61795, n61796, n61797, n61798,
    n61799, n61800, n61801, n61802, n61803, n61804, n61805, n61806, n61807,
    n61808, n61809, n61810, n61811, n61812, n61813, n61814, n61815, n61816,
    n61817, n61818, n61819, n61820, n61821, n61822, n61823, n61824, n61825,
    n61826, n61827, n61828, n61829, n61830, n61831, n61832, n61833, n61834,
    n61835, n61836, n61837, n61838, n61839, n61840, n61841, n61842, n61843,
    n61844, n61845, n61846, n61847, n61848, n61849, n61850, n61851, n61852,
    n61853, n61854, n61855, n61856, n61857, n61858, n61859, n61860, n61861,
    n61862, n61863, n61864, n61865, n61866, n61867, n61868, n61870, n61871,
    n61872, n61873, n61874, n61875, n61876, n61877, n61878, n61879, n61880,
    n61881, n61882, n61883, n61884, n61885, n61886, n61887, n61888, n61889,
    n61890, n61891, n61892, n61893, n61894, n61895, n61896, n61897, n61898,
    n61899, n61900, n61901, n61902, n61903, n61904, n61905, n61906, n61907,
    n61908, n61909, n61910, n61911, n61912, n61913, n61914, n61915, n61916,
    n61917, n61918, n61919, n61920, n61921, n61922, n61923, n61924, n61925,
    n61926, n61927, n61928, n61929, n61930, n61931, n61932, n61933, n61934,
    n61935, n61936, n61937, n61938, n61939, n61940, n61941, n61942, n61943,
    n61944, n61945, n61946, n61947, n61948, n61949, n61950, n61951, n61952,
    n61953, n61954, n61955, n61956, n61957, n61958, n61959, n61960, n61961,
    n61962, n61963, n61964, n61965, n61966, n61968, n61969, n61970, n61971,
    n61972, n61973, n61974, n61975, n61976, n61977, n61978, n61979, n61980,
    n61981, n61982, n61983, n61984, n61985, n61986, n61987, n61988, n61989,
    n61990, n61991, n61992, n61993, n61994, n61995, n61996, n61997, n61998,
    n61999, n62000, n62001, n62002, n62003, n62004, n62005, n62006, n62007,
    n62008, n62009, n62010, n62011, n62012, n62013, n62014, n62015, n62016,
    n62017, n62018, n62019, n62020, n62021, n62022, n62023, n62024, n62025,
    n62026, n62027, n62028, n62029, n62030, n62031, n62032, n62033, n62034,
    n62035, n62036, n62037, n62038, n62039, n62040, n62041, n62042, n62043,
    n62044, n62045, n62046, n62047, n62048, n62049, n62050, n62051, n62052,
    n62053, n62054, n62055, n62056, n62058, n62059, n62060, n62061, n62062,
    n62063, n62064, n62065, n62066, n62067, n62068, n62069, n62070, n62071,
    n62072, n62073, n62074, n62075, n62076, n62077, n62078, n62079, n62080,
    n62081, n62082, n62083, n62084, n62085, n62086, n62087, n62088, n62089,
    n62090, n62091, n62092, n62093, n62094, n62095, n62096, n62097, n62098,
    n62099, n62100, n62101, n62102, n62103, n62104, n62105, n62106, n62107,
    n62108, n62109, n62110, n62111, n62112, n62113, n62114, n62115, n62116,
    n62117, n62118, n62119, n62120, n62121, n62122, n62123, n62124, n62125,
    n62126, n62127, n62128, n62129, n62130, n62131, n62132, n62133, n62134,
    n62135, n62136, n62137, n62138, n62139, n62141, n62142, n62143, n62144,
    n62145, n62146, n62147, n62148, n62149, n62150, n62151, n62152, n62153,
    n62154, n62155, n62156, n62157, n62158, n62159, n62160, n62161, n62162,
    n62163, n62164, n62165, n62166, n62167, n62168, n62169, n62170, n62171,
    n62172, n62173, n62174, n62175, n62176, n62177, n62178, n62179, n62180,
    n62181, n62182, n62183, n62184, n62185, n62186, n62187, n62188, n62189,
    n62190, n62191, n62192, n62193, n62194, n62195, n62196, n62197, n62198,
    n62199, n62200, n62201, n62202, n62203, n62204, n62205, n62206, n62207,
    n62208, n62209, n62210, n62211, n62212, n62213, n62214, n62215, n62217,
    n62218, n62219, n62220, n62221, n62222, n62223, n62224, n62225, n62226,
    n62227, n62228, n62229, n62230, n62231, n62232, n62233, n62234, n62235,
    n62236, n62237, n62238, n62239, n62240, n62241, n62242, n62243, n62244,
    n62245, n62246, n62247, n62248, n62249, n62250, n62251, n62252, n62253,
    n62254, n62255, n62256, n62257, n62258, n62259, n62260, n62261, n62262,
    n62263, n62264, n62265, n62266, n62267, n62268, n62269, n62270, n62271,
    n62272, n62273, n62274, n62275, n62276, n62277, n62278, n62279, n62280,
    n62281, n62282, n62283, n62284, n62285, n62286, n62287, n62289, n62290,
    n62291, n62292, n62293, n62294, n62295, n62296, n62297, n62298, n62299,
    n62300, n62301, n62302, n62303, n62304, n62305, n62306, n62307, n62308,
    n62309, n62310, n62311, n62312, n62313, n62314, n62315, n62316, n62317,
    n62318, n62319, n62320, n62321, n62322, n62323, n62324, n62325, n62326,
    n62327, n62328, n62329, n62330, n62331, n62332, n62333, n62334, n62335,
    n62336, n62337, n62338, n62339, n62340, n62341, n62342, n62343, n62344,
    n62345, n62346, n62347, n62348, n62349, n62350, n62351, n62352, n62353,
    n62354, n62355, n62356, n62357, n62358, n62359, n62360, n62361, n62362,
    n62363, n62364, n62365, n62367, n62368, n62369, n62370, n62371, n62372,
    n62373, n62374, n62375, n62376, n62377, n62378, n62379, n62380, n62381,
    n62382, n62383, n62384, n62385, n62386, n62387, n62388, n62389, n62390,
    n62391, n62392, n62393, n62394, n62395, n62396, n62397, n62398, n62399,
    n62400, n62401, n62402, n62403, n62404, n62405, n62406, n62407, n62408,
    n62409, n62410, n62411, n62412, n62413, n62414, n62415, n62416, n62417,
    n62418, n62419, n62420, n62421, n62422, n62423, n62424, n62425, n62426,
    n62427, n62428, n62429, n62430, n62431, n62432, n62433, n62434, n62435,
    n62436, n62437, n62438, n62439, n62440, n62442, n62443, n62444, n62445,
    n62446, n62447, n62448, n62449, n62450, n62451, n62452, n62453, n62454,
    n62455, n62456, n62457, n62458, n62459, n62460, n62461, n62462, n62463,
    n62464, n62465, n62466, n62467, n62468, n62469, n62470, n62471, n62472,
    n62473, n62474, n62475, n62476, n62477, n62478, n62479, n62480, n62481,
    n62482, n62483, n62484, n62485, n62486, n62487, n62488, n62489, n62490,
    n62491, n62492, n62493, n62494, n62495, n62496, n62497, n62498, n62499,
    n62500, n62501, n62502, n62503, n62504, n62505, n62506, n62507, n62508,
    n62509, n62510, n62511, n62512, n62513, n62515, n62516, n62517, n62518,
    n62519, n62520, n62521, n62522, n62523, n62524, n62525, n62526, n62527,
    n62528, n62529, n62530, n62531, n62532, n62533, n62534, n62535, n62536,
    n62537, n62538, n62539, n62540, n62541, n62542, n62543, n62544, n62545,
    n62546, n62547, n62548, n62549, n62550, n62551, n62552, n62553, n62554,
    n62555, n62556, n62557, n62558, n62559, n62560, n62561, n62562, n62563,
    n62564, n62565, n62566, n62567, n62568, n62569, n62570, n62571, n62572,
    n62573, n62574, n62575, n62576, n62577, n62578, n62579, n62580, n62581,
    n62582, n62583, n62584, n62585, n62586, n62587, n62588, n62589, n62590,
    n62591, n62593, n62594, n62595, n62596, n62597, n62598, n62599, n62600,
    n62601, n62602, n62603, n62604, n62605, n62606, n62607, n62608, n62609,
    n62610, n62611, n62612, n62613, n62614, n62615, n62616, n62617, n62618,
    n62619, n62620, n62621, n62622, n62623, n62624, n62625, n62626, n62627,
    n62628, n62629, n62630, n62631, n62632, n62633, n62634, n62635, n62636,
    n62637, n62638, n62639, n62640, n62641, n62642, n62643, n62644, n62645,
    n62646, n62647, n62648, n62649, n62650, n62651, n62652, n62653, n62654,
    n62655, n62656, n62657, n62658, n62659, n62660, n62661, n62662, n62663,
    n62665, n62666, n62667, n62668, n62669, n62670, n62671, n62672, n62673,
    n62674, n62675, n62676, n62677, n62678, n62679, n62680, n62681, n62682,
    n62683, n62684, n62685, n62686, n62687, n62688, n62689, n62690, n62691,
    n62692, n62693, n62694, n62695, n62696, n62697, n62698, n62699, n62700,
    n62701, n62702, n62703, n62704, n62705, n62706, n62707, n62708, n62709,
    n62710, n62711, n62712, n62713, n62714, n62715, n62716, n62717, n62718,
    n62719, n62720, n62721, n62722, n62723, n62724, n62725, n62726, n62727,
    n62728, n62729, n62730, n62731, n62732, n62733, n62734, n62735, n62736,
    n62737, n62738, n62739, n62740, n62741, n62742, n62744, n62745, n62746,
    n62747, n62748, n62749, n62750, n62751, n62752, n62753, n62754, n62755,
    n62756, n62757, n62758, n62759, n62760, n62761, n62762, n62763, n62764,
    n62765, n62766, n62767, n62768, n62769, n62770, n62771, n62772, n62773,
    n62774, n62775, n62776, n62777, n62778, n62779, n62780, n62781, n62782,
    n62783, n62784, n62785, n62786, n62787, n62788, n62789, n62790, n62791,
    n62792, n62793, n62794, n62795, n62796, n62797, n62798, n62799, n62800,
    n62801, n62802, n62803, n62804, n62805, n62806, n62807, n62808, n62809,
    n62810, n62811, n62812, n62813, n62815, n62816, n62817, n62818, n62819,
    n62820, n62821, n62822, n62823, n62824, n62825, n62826, n62827, n62828,
    n62829, n62830, n62831, n62832, n62833, n62834, n62835, n62836, n62837,
    n62838, n62839, n62840, n62841, n62842, n62843, n62844, n62845, n62846,
    n62847, n62848, n62849, n62850, n62851, n62852, n62853, n62854, n62855,
    n62856, n62857, n62858, n62859, n62860, n62861, n62862, n62863, n62864,
    n62865, n62866, n62867, n62868, n62869, n62870, n62871, n62872, n62873,
    n62874, n62875, n62876, n62877, n62878, n62879, n62880, n62881, n62882,
    n62883, n62884, n62885, n62886, n62887, n62888, n62889, n62890, n62891,
    n62893, n62894, n62895, n62896, n62897, n62898, n62899, n62900, n62901,
    n62902, n62903, n62904, n62905, n62906, n62907, n62908, n62909, n62910,
    n62911, n62912, n62913, n62914, n62915, n62916, n62917, n62918, n62919,
    n62920, n62921, n62922, n62923, n62924, n62925, n62926, n62927, n62928,
    n62929, n62930, n62931, n62932, n62933, n62934, n62935, n62936, n62937,
    n62938, n62939, n62940, n62941, n62942, n62943, n62944, n62945, n62946,
    n62947, n62948, n62949, n62950, n62951, n62952, n62953, n62954, n62955,
    n62956, n62957, n62958, n62959, n62960, n62961, n62962, n62963, n62964,
    n62965, n62966, n62967, n62969, n62970, n62971, n62972, n62973, n62974,
    n62975, n62976, n62977, n62978, n62979, n62980, n62981, n62982, n62983,
    n62984, n62985, n62986, n62987, n62988, n62989, n62990, n62991, n62992,
    n62993, n62994, n62995, n62996, n62997, n62998, n62999, n63000, n63001,
    n63002, n63003, n63004, n63005, n63006, n63007, n63008, n63009, n63010,
    n63011, n63012, n63013, n63014, n63015, n63016, n63017, n63018, n63019,
    n63020, n63021, n63022, n63023, n63024, n63025, n63026, n63027, n63028,
    n63029, n63030, n63031, n63032, n63033, n63034, n63035, n63036, n63037,
    n63038, n63039, n63040, n63042, n63043, n63044, n63045, n63046, n63047,
    n63048, n63049, n63050, n63051, n63052, n63053, n63054, n63055, n63056,
    n63057, n63058, n63059, n63060, n63061, n63062, n63063, n63064, n63065,
    n63066, n63067, n63068, n63069, n63070, n63071, n63072, n63073, n63074,
    n63075, n63076, n63077, n63078, n63079, n63080, n63081, n63082, n63083,
    n63084, n63085, n63086, n63087, n63088, n63089, n63090, n63091, n63092,
    n63093, n63094, n63095, n63096, n63097, n63098, n63099, n63100, n63101,
    n63102, n63103, n63104, n63105, n63106, n63107, n63108, n63109, n63110,
    n63111, n63112, n63113, n63114, n63115, n63116, n63117, n63119, n63120,
    n63121, n63122, n63123, n63124, n63125, n63126, n63127, n63128, n63129,
    n63130, n63131, n63132, n63133, n63134, n63135, n63136, n63137, n63138,
    n63139, n63140, n63141, n63142, n63143, n63144, n63145, n63146, n63147,
    n63148, n63149, n63150, n63151, n63152, n63153, n63154, n63155, n63156,
    n63157, n63158, n63159, n63160, n63161, n63162, n63163, n63164, n63165,
    n63166, n63167, n63168, n63169, n63170, n63171, n63172, n63173, n63174,
    n63175, n63176, n63177, n63178, n63179, n63180, n63181, n63182, n63183,
    n63184, n63185, n63186, n63187, n63188, n63189, n63190, n63191, n63192,
    n63193, n63194, n63196, n63197, n63198, n63199, n63200, n63201, n63202,
    n63203, n63204, n63205, n63206, n63207, n63208, n63209, n63210, n63211,
    n63212, n63213, n63214, n63215, n63216, n63217, n63218, n63219, n63220,
    n63221, n63222, n63223, n63224, n63225, n63226, n63227, n63228, n63229,
    n63230, n63231, n63232, n63233, n63234, n63235, n63236, n63237, n63238,
    n63239, n63240, n63241, n63242, n63243, n63244, n63245, n63246, n63247,
    n63248, n63249, n63250, n63251, n63252, n63253, n63254, n63255, n63256,
    n63257, n63258, n63259, n63260, n63261, n63262, n63263, n63264, n63265,
    n63266, n63267, n63268, n63270, n63271, n63272, n63273, n63274, n63275,
    n63276, n63277, n63278, n63279, n63280, n63281, n63282, n63283, n63284,
    n63285, n63286, n63287, n63288, n63289, n63290, n63291, n63292, n63293,
    n63294, n63295, n63296, n63297, n63298, n63299, n63300, n63301, n63302,
    n63303, n63304, n63305, n63306, n63307, n63308, n63309, n63310, n63311,
    n63312, n63313, n63314, n63315, n63316, n63317, n63318, n63319, n63320,
    n63321, n63322, n63323, n63324, n63325, n63326, n63327, n63328, n63329,
    n63330, n63331, n63332, n63333, n63334, n63335, n63336, n63337, n63338,
    n63339, n63340, n63341, n63342, n63343, n63344, n63345, n63346, n63348,
    n63349, n63350, n63351, n63352, n63353, n63354, n63355, n63356, n63357,
    n63358, n63359, n63360, n63361, n63362, n63363, n63364, n63365, n63366,
    n63367, n63368, n63369, n63370, n63371, n63372, n63373, n63374, n63375,
    n63376, n63377, n63378, n63379, n63380, n63381, n63382, n63383, n63384,
    n63385, n63386, n63387, n63388, n63389, n63390, n63391, n63392, n63393,
    n63394, n63395, n63396, n63397, n63398, n63399, n63400, n63401, n63402,
    n63403, n63404, n63405, n63406, n63407, n63408, n63409, n63410, n63411,
    n63412, n63413, n63414, n63415, n63416, n63417, n63418, n63419, n63420,
    n63421, n63423, n63424, n63425, n63426, n63427, n63428, n63429, n63430,
    n63431, n63432, n63433, n63434, n63435, n63436, n63437, n63438, n63439,
    n63440, n63441, n63442, n63443, n63444, n63445, n63446, n63447, n63448,
    n63449, n63450, n63451, n63452, n63453, n63454, n63455, n63456, n63457,
    n63458, n63459, n63460, n63461, n63462, n63463, n63464, n63465, n63466,
    n63467, n63468, n63469, n63470, n63471, n63472, n63473, n63474, n63475,
    n63476, n63477, n63478, n63479, n63480, n63481, n63482, n63483, n63484,
    n63485, n63486, n63487, n63488, n63489, n63490, n63491, n63492, n63494,
    n63495, n63496, n63497, n63498, n63499, n63500, n63501, n63502, n63503,
    n63504, n63505, n63506, n63507, n63508, n63509, n63510, n63511, n63512,
    n63513, n63514, n63515, n63516, n63517, n63518, n63519, n63520, n63521,
    n63522, n63523, n63524, n63525, n63526, n63527, n63528, n63529, n63530,
    n63531, n63532, n63533, n63534, n63535, n63536, n63537, n63538, n63539,
    n63540, n63541, n63542, n63543, n63544, n63545, n63546, n63547, n63548,
    n63549, n63550, n63551, n63552, n63553, n63554, n63555, n63556, n63557,
    n63558, n63559, n63560, n63561, n63562, n63563, n63564, n63565, n63566,
    n63567, n63568, n63569, n63570, n63571, n63572, n63574, n63575, n63576,
    n63577, n63578, n63579, n63580, n63581, n63582, n63583, n63584, n63585,
    n63586, n63587, n63588, n63589, n63590, n63591, n63592, n63593, n63594,
    n63595, n63596, n63597, n63598, n63599, n63600, n63601, n63602, n63603,
    n63604, n63605, n63606, n63607, n63608, n63609, n63610, n63611, n63612,
    n63613, n63614, n63615, n63616, n63617, n63618, n63619, n63620, n63621,
    n63622, n63623, n63624, n63625, n63626, n63627, n63628, n63629, n63630,
    n63631, n63632, n63633, n63634, n63635, n63636, n63637, n63638, n63639,
    n63640, n63641, n63642, n63643, n63645, n63646, n63647, n63648, n63649,
    n63650, n63651, n63652, n63653, n63654, n63655, n63656, n63657, n63658,
    n63659, n63660, n63661, n63662, n63663, n63664, n63665, n63666, n63667,
    n63668, n63669, n63670, n63671, n63672, n63673, n63674, n63675, n63676,
    n63677, n63678, n63679, n63680, n63681, n63682, n63683, n63684, n63685,
    n63686, n63687, n63688, n63689, n63690, n63691, n63692, n63693, n63694,
    n63695, n63696, n63697, n63698, n63699, n63700, n63701, n63702, n63703,
    n63704, n63705, n63706, n63707, n63708, n63709, n63710, n63711, n63712,
    n63713, n63714, n63715, n63717, n63718, n63719, n63720, n63721, n63722,
    n63723, n63724, n63725, n63726, n63727, n63728, n63729, n63730, n63731,
    n63732, n63733, n63734, n63735, n63736, n63737, n63738, n63739, n63740,
    n63741, n63742, n63743, n63744, n63745, n63746, n63747, n63748, n63749,
    n63750, n63751, n63752, n63753, n63754, n63755, n63756, n63757, n63758,
    n63759, n63760, n63761, n63762, n63763, n63764, n63765, n63766, n63767,
    n63768, n63769, n63770, n63771, n63772, n63773, n63774, n63775, n63776,
    n63777, n63778, n63779, n63780, n63781, n63782, n63783, n63784, n63785,
    n63786, n63787, n63788, n63789, n63790, n63791, n63792, n63793, n63794,
    n63795, n63796, n63797, n63799, n63800, n63801, n63802, n63803, n63804,
    n63805, n63806, n63807, n63808, n63809, n63810, n63811, n63812, n63813,
    n63814, n63815, n63816, n63817, n63818, n63819, n63820, n63821, n63822,
    n63823, n63824, n63825, n63826, n63827, n63828, n63829, n63830, n63832,
    n63833, n63834, n63835, n63836, n63837, n63838, n63839, n63840, n63841,
    n63842, n63843, n63844, n63845, n63847, n63848, n63849, n63850, n63851,
    n63852, n63853, n63854, n63855, n63856, n63857, n63858, n63859, n63860,
    n63861, n63862, n63863, n63865, n63866, n63867, n63868, n63869, n63870,
    n63871, n63872, n63873, n63874, n63875, n63876, n63877, n63878, n63879,
    n63880, n63881, n63882, n63883, n63884, n63885, n63887, n63888, n63889,
    n63890, n63891, n63892, n63893, n63894, n63895, n63896, n63897, n63898,
    n63899, n63900, n63901, n63902, n63903, n63904, n63905, n63906, n63907,
    n63908, n63910, n63911, n63912, n63913, n63914, n63915, n63916, n63917,
    n63918, n63919, n63920, n63921, n63922, n63923, n63924, n63925, n63926,
    n63927, n63928, n63929, n63930, n63931, n63933, n63934, n63935, n63936,
    n63937, n63938, n63939, n63940, n63941, n63942, n63943, n63944, n63945,
    n63946, n63947, n63948, n63949, n63950, n63951, n63952, n63953, n63954,
    n63956, n63957, n63958, n63959, n63960, n63961, n63962, n63963, n63964,
    n63965, n63966, n63967, n63968, n63969, n63970, n63971, n63972, n63973,
    n63974, n63975, n63976, n63977, n63979, n63980, n63981, n63982, n63983,
    n63984, n63985, n63986, n63987, n63988, n63989, n63990, n63991, n63992,
    n63993, n63994, n63995, n63996, n63997, n63998, n63999, n64000, n64002,
    n64003, n64004, n64005, n64006, n64007, n64008, n64009, n64010, n64011,
    n64012, n64013, n64014, n64015, n64016, n64017, n64018, n64019, n64020,
    n64021, n64022, n64023, n64025, n64026, n64027, n64028, n64029, n64030,
    n64031, n64032, n64033, n64034, n64035, n64036, n64037, n64038, n64039,
    n64040, n64041, n64042, n64043, n64044, n64045, n64046, n64048, n64049,
    n64050, n64051, n64052, n64053, n64054, n64055, n64056, n64057, n64058,
    n64059, n64060, n64061, n64062, n64063, n64064, n64065, n64066, n64067,
    n64068, n64069, n64071, n64072, n64073, n64074, n64075, n64076, n64077,
    n64078, n64079, n64080, n64081, n64082, n64083, n64084, n64085, n64086,
    n64087, n64088, n64089, n64090, n64091, n64092, n64094, n64095, n64096,
    n64097, n64098, n64099, n64100, n64101, n64102, n64103, n64104, n64105,
    n64106, n64107, n64108, n64109, n64110, n64111, n64112, n64113, n64114,
    n64115, n64117, n64118, n64119, n64120, n64121, n64122, n64123, n64124,
    n64125, n64126, n64127, n64128, n64129, n64130, n64131, n64132, n64133,
    n64134, n64135, n64136, n64137, n64138, n64140, n64141, n64142, n64143,
    n64144, n64145, n64146, n64147, n64148, n64149, n64150, n64151, n64152,
    n64153, n64154, n64155, n64156, n64157, n64158, n64159, n64160, n64161,
    n64163, n64164, n64165, n64166, n64167, n64168, n64169, n64170, n64171,
    n64172, n64173, n64174, n64175, n64176, n64177, n64178, n64179, n64180,
    n64181, n64182, n64183, n64184, n64186, n64187, n64188, n64189, n64190,
    n64191, n64192, n64193, n64194, n64195, n64196, n64197, n64198, n64199,
    n64200, n64201, n64202, n64203, n64204, n64205, n64206, n64207, n64209,
    n64210, n64211, n64212, n64213, n64214, n64215, n64216, n64217, n64218,
    n64219, n64220, n64221, n64222, n64223, n64224, n64225, n64226, n64227,
    n64228, n64229, n64230, n64232, n64233, n64234, n64235, n64236, n64237,
    n64238, n64239, n64240, n64241, n64242, n64243, n64244, n64245, n64246,
    n64247, n64248, n64249, n64250, n64251, n64252, n64253, n64255, n64256,
    n64257, n64258, n64259, n64260, n64261, n64262, n64263, n64264, n64265,
    n64266, n64267, n64268, n64269, n64270, n64271, n64272, n64273, n64274,
    n64275, n64276, n64278, n64279, n64280, n64281, n64282, n64283, n64284,
    n64285, n64286, n64287, n64288, n64289, n64290, n64291, n64292, n64293,
    n64294, n64295, n64296, n64297, n64298, n64299, n64301, n64302, n64303,
    n64304, n64305, n64306, n64307, n64308, n64309, n64310, n64311, n64312,
    n64313, n64314, n64315, n64316, n64317, n64318, n64319, n64320, n64321,
    n64322, n64324, n64325, n64326, n64327, n64328, n64329, n64330, n64331,
    n64332, n64333, n64334, n64335, n64336, n64337, n64338, n64339, n64340,
    n64341, n64342, n64343, n64344, n64345, n64347, n64348, n64349, n64350,
    n64351, n64352, n64353, n64354, n64355, n64356, n64357, n64358, n64359,
    n64360, n64361, n64362, n64363, n64364, n64365, n64366, n64367, n64368,
    n64370, n64371, n64372, n64373, n64374, n64375, n64376, n64377, n64378,
    n64379, n64380, n64381, n64382, n64383, n64384, n64385, n64386, n64387,
    n64388, n64389, n64390, n64391, n64393, n64394, n64395, n64396, n64397,
    n64398, n64399, n64400, n64401, n64402, n64403, n64404, n64405, n64406,
    n64407, n64408, n64409, n64410, n64411, n64412, n64413, n64414, n64416,
    n64417, n64418, n64419, n64420, n64421, n64422, n64423, n64424, n64425,
    n64426, n64427, n64428, n64429, n64430, n64431, n64432, n64433, n64434,
    n64435, n64436, n64437, n64439, n64440, n64441, n64442, n64443, n64444,
    n64445, n64446, n64447, n64448, n64449, n64450, n64451, n64452, n64453,
    n64454, n64455, n64456, n64457, n64458, n64459, n64460, n64462, n64463,
    n64464, n64465, n64466, n64467, n64468, n64469, n64470, n64471, n64472,
    n64473, n64474, n64475, n64476, n64477, n64478, n64479, n64480, n64481,
    n64482, n64483, n64485, n64486, n64487, n64488, n64489, n64490, n64491,
    n64492, n64493, n64494, n64495, n64496, n64497, n64498, n64499, n64500,
    n64501, n64502, n64503, n64504, n64505, n64506, n64508, n64509, n64510,
    n64511, n64512, n64513, n64514, n64515, n64516, n64517, n64518, n64519,
    n64520, n64521, n64522, n64523, n64524, n64525, n64526, n64527, n64528,
    n64529, n64531, n64532, n64533, n64534, n64535, n64536, n64537, n64538,
    n64539, n64540, n64542, n64543, n64544, n64545, n64547, n64548, n64549,
    n64550, n64552, n64553, n64554, n64555, n64557, n64558, n64559, n64560,
    n64562, n64563, n64564, n64565, n64567, n64568, n64569, n64570, n64572,
    n64573, n64574, n64575, n64577, n64578, n64579, n64580, n64582, n64583,
    n64584, n64585, n64587, n64588, n64589, n64590, n64592, n64593, n64594,
    n64595, n64597, n64598, n64599, n64600, n64602, n64603, n64604, n64605,
    n64607, n64608, n64609, n64610, n64612, n64613, n64614, n64615, n64617,
    n64618, n64619, n64621, n64622, n64623, n64625, n64626, n64627, n64629,
    n64630, n64631, n64633, n64634, n64635, n64637, n64638, n64639, n64641,
    n64642, n64643, n64645, n64646, n64647, n64649, n64650, n64651, n64653,
    n64654, n64655, n64657, n64658, n64659, n64661, n64662, n64663, n64665,
    n64666, n64667, n64669, n64670, n64671, n64673, n64674, n64675, n64677,
    n64678, n64679, n64680, n64681, n64682, n64683, n64684, n64685, n64686,
    n64688, n64689, n64690, n64691, n64693, n64694, n64695, n64696, n64698,
    n64699, n64700, n64701, n64703, n64704, n64705, n64706, n64708, n64709,
    n64710, n64711, n64713, n64714, n64715, n64716, n64718, n64719, n64720,
    n64721, n64723, n64724, n64725, n64726, n64728, n64729, n64730, n64731,
    n64733, n64734, n64735, n64736, n64738, n64739, n64740, n64741, n64743,
    n64744, n64745, n64746, n64748, n64749, n64750, n64751, n64753, n64754,
    n64755, n64756, n64758, n64759, n64760, n64761, n64763, n64764, n64765,
    n64766, n64767, n64769, n64770, n64771, n64772, n64774, n64775, n64776,
    n64777, n64779, n64780, n64781, n64782, n64784, n64785, n64786, n64787,
    n64789, n64790, n64791, n64792, n64794, n64795, n64796, n64797, n64799,
    n64800, n64801, n64802, n64804, n64805, n64806, n64807, n64809, n64810,
    n64811, n64812, n64814, n64815, n64816, n64817, n64819, n64820, n64821,
    n64822, n64824, n64825, n64826, n64827, n64829, n64830, n64831, n64832,
    n64834, n64835, n64836, n64837, n64840, n64841, n64842, n64843, n64844,
    n64845, n64846, n64847, n64848, n64849, n64850, n64851, n64853, n64854,
    n64855, n64856, n64857, n64858, n64859, n64860, n64861, n64863, n64864,
    n64865, n64866, n64867, n64868, n64869, n64870, n64871, n64872, n64874,
    n64875, n64876, n64877, n64878, n64879, n64880, n64881, n64882, n64883,
    n64884, n64886, n64887, n64888, n64889, n64890, n64891, n64892, n64893,
    n64894, n64895, n64897, n64898, n64899, n64900, n64901, n64902, n64903,
    n64904, n64905, n64906, n64907, n64909, n64910, n64911, n64912, n64913,
    n64914, n64915, n64916, n64917, n64918, n64920, n64921, n64922, n64923,
    n64924, n64925, n64926, n64927, n64928, n64929, n64930, n64932, n64933,
    n64934, n64935, n64936, n64937, n64938, n64939, n64940, n64941, n64942,
    n64943, n64944, n64945, n64946, n64947, n64948, n64949, n64950, n64951,
    n64952, n64953, n64954, n64955, n64956, n64957, n64958, n64959, n64960,
    n64961, n64962, n64963, n64964, n64965, n64966, n64967, n64968, n64969,
    n64970, n64971, n64972, n64973, n64974, n64975, n64976, n64977, n64978,
    n64979, n64980, n64981, n64982, n64983, n64984, n64985, n64986, n64987,
    n64988, n64989, n64990, n64991, n64992, n64993, n64995, n64996, n64997,
    n64998, n64999, n65000, n65001, n65002, n65003, n65004, n65005, n65006,
    n65007, n65008, n65009, n65010, n65011, n65012, n65013, n65014, n65015,
    n65016, n65017, n65018, n65019, n65020, n65021, n65022, n65023, n65024,
    n65025, n65026, n65027, n65028, n65029, n65030, n65031, n65032, n65033,
    n65034, n65035, n65036, n65038, n65039, n65040, n65041, n65042, n65043,
    n65044, n65045, n65046, n65047, n65048, n65049, n65050, n65051, n65052,
    n65053, n65054, n65055, n65056, n65057, n65058, n65059, n65060, n65061,
    n65062, n65063, n65064, n65065, n65066, n65067, n65068, n65069, n65070,
    n65071, n65072, n65073, n65074, n65075, n65076, n65077, n65078, n65080,
    n65081, n65082, n65083, n65084, n65085, n65086, n65087, n65088, n65089,
    n65090, n65091, n65092, n65093, n65094, n65095, n65096, n65097, n65098,
    n65099, n65100, n65101, n65102, n65103, n65104, n65105, n65106, n65107,
    n65108, n65109, n65110, n65111, n65112, n65113, n65114, n65115, n65116,
    n65117, n65118, n65119, n65120, n65121, n65123, n65124, n65125, n65126,
    n65127, n65128, n65129, n65130, n65131, n65132, n65133, n65134, n65135,
    n65136, n65137, n65138, n65139, n65140, n65141, n65142, n65143, n65144,
    n65145, n65146, n65147, n65148, n65149, n65150, n65151, n65152, n65153,
    n65154, n65155, n65156, n65157, n65158, n65159, n65160, n65161, n65162,
    n65163, n65165, n65166, n65167, n65168, n65169, n65170, n65171, n65172,
    n65173, n65174, n65175, n65176, n65177, n65178, n65179, n65180, n65181,
    n65182, n65183, n65184, n65185, n65186, n65187, n65188, n65189, n65190,
    n65191, n65192, n65193, n65194, n65195, n65196, n65197, n65198, n65199,
    n65200, n65201, n65202, n65203, n65204, n65205, n65206, n65208, n65209,
    n65210, n65211, n65212, n65213, n65214, n65215, n65216, n65217, n65218,
    n65219, n65220, n65221, n65222, n65223, n65224, n65225, n65226, n65227,
    n65228, n65229, n65230, n65231, n65232, n65233, n65234, n65235, n65236,
    n65237, n65238, n65239, n65240, n65241, n65242, n65243, n65244, n65245,
    n65246, n65247, n65248, n65250, n65251, n65252, n65253, n65254, n65255,
    n65256, n65257, n65258, n65259, n65260, n65261, n65262, n65263, n65264,
    n65265, n65266, n65267, n65268, n65269, n65270, n65271, n65272, n65273,
    n65274, n65275, n65276, n65277, n65278, n65279, n65280, n65281, n65282,
    n65283, n65284, n65285, n65286, n65287, n65288, n65289, n65290, n65291,
    n65293, n65294, n65295, n65296, n65297, n65298, n65299, n65300, n65301,
    n65302, n65303, n65304, n65305, n65306, n65307, n65308, n65309, n65310,
    n65311, n65312, n65313, n65314, n65315, n65316, n65317, n65318, n65319,
    n65320, n65321, n65322, n65323, n65324, n65325, n65326, n65327, n65328,
    n65329, n65330, n65331, n65332, n65333, n65334, n65335, n65336, n65337,
    n65338, n65339, n65340, n65341, n65342, n65343, n65344, n65345, n65346,
    n65347, n65348, n65349, n65350, n65351, n65352, n65353, n65354, n65355,
    n65356, n65357, n65358, n65359, n65360, n65361, n65362, n65364, n65365,
    n65366, n65367, n65368, n65369, n65370, n65371, n65372, n65373, n65374,
    n65375, n65376, n65377, n65378, n65379, n65380, n65381, n65382, n65383,
    n65384, n65385, n65386, n65387, n65388, n65389, n65390, n65391, n65392,
    n65393, n65394, n65395, n65396, n65397, n65398, n65399, n65400, n65401,
    n65402, n65403, n65404, n65405, n65406, n65407, n65409, n65410, n65411,
    n65412, n65413, n65414, n65415, n65416, n65417, n65418, n65419, n65420,
    n65421, n65422, n65423, n65424, n65425, n65426, n65427, n65428, n65429,
    n65430, n65431, n65432, n65433, n65434, n65435, n65436, n65437, n65438,
    n65439, n65440, n65441, n65442, n65443, n65444, n65445, n65446, n65447,
    n65448, n65449, n65450, n65451, n65453, n65454, n65455, n65456, n65457,
    n65458, n65459, n65460, n65461, n65462, n65463, n65464, n65465, n65466,
    n65467, n65468, n65469, n65470, n65471, n65472, n65473, n65474, n65475,
    n65476, n65477, n65478, n65479, n65480, n65481, n65482, n65483, n65484,
    n65485, n65486, n65487, n65488, n65489, n65490, n65491, n65492, n65493,
    n65494, n65495, n65496, n65498, n65499, n65500, n65501, n65502, n65503,
    n65504, n65505, n65506, n65507, n65508, n65509, n65510, n65511, n65512,
    n65513, n65514, n65515, n65516, n65517, n65518, n65519, n65520, n65521,
    n65522, n65523, n65524, n65525, n65526, n65527, n65528, n65529, n65530,
    n65531, n65532, n65533, n65534, n65535, n65536, n65537, n65538, n65539,
    n65540, n65542, n65543, n65544, n65545, n65546, n65547, n65548, n65549,
    n65550, n65551, n65552, n65553, n65554, n65555, n65556, n65557, n65558,
    n65559, n65560, n65561, n65562, n65563, n65564, n65565, n65566, n65567,
    n65568, n65569, n65570, n65571, n65572, n65573, n65574, n65575, n65576,
    n65577, n65578, n65579, n65580, n65581, n65582, n65583, n65584, n65585,
    n65587, n65588, n65589, n65590, n65591, n65592, n65593, n65594, n65595,
    n65596, n65597, n65598, n65599, n65600, n65601, n65602, n65603, n65604,
    n65605, n65606, n65607, n65608, n65609, n65610, n65611, n65612, n65613,
    n65614, n65615, n65616, n65617, n65618, n65619, n65620, n65621, n65622,
    n65623, n65624, n65625, n65626, n65627, n65628, n65629, n65631, n65632,
    n65633, n65634, n65635, n65636, n65637, n65638, n65639, n65640, n65641,
    n65642, n65643, n65644, n65645, n65646, n65647, n65648, n65649, n65650,
    n65651, n65652, n65653, n65654, n65655, n65656, n65657, n65658, n65659,
    n65660, n65661, n65662, n65663, n65664, n65665, n65666, n65667, n65668,
    n65669, n65670, n65671, n65672, n65673, n65674, n65675, n65676, n65677,
    n65678, n65679, n65680, n65681, n65682, n65683, n65684, n65685, n65686,
    n65687, n65688, n65689, n65690, n65691, n65692, n65693, n65694, n65695,
    n65696, n65697, n65698, n65699, n65700, n65701, n65702, n65703, n65704,
    n65705, n65706, n65707, n65708, n65709, n65710, n65711, n65712, n65713,
    n65714, n65715, n65716, n65717, n65718, n65719, n65720, n65721, n65722,
    n65723, n65724, n65725, n65726, n65727, n65728, n65730, n65731, n65732,
    n65733, n65734, n65735, n65736, n65737, n65738, n65739, n65740, n65741,
    n65742, n65743, n65744, n65745, n65746, n65747, n65748, n65749, n65750,
    n65751, n65752, n65753, n65754, n65755, n65756, n65757, n65758, n65759,
    n65760, n65761, n65762, n65763, n65764, n65765, n65766, n65767, n65768,
    n65769, n65770, n65771, n65772, n65773, n65774, n65775, n65776, n65778,
    n65779, n65780, n65781, n65782, n65783, n65784, n65785, n65786, n65787,
    n65788, n65789, n65790, n65791, n65792, n65793, n65794, n65795, n65796,
    n65797, n65798, n65799, n65800, n65801, n65802, n65803, n65804, n65805,
    n65806, n65807, n65808, n65809, n65810, n65811, n65812, n65813, n65814,
    n65815, n65816, n65817, n65818, n65819, n65820, n65821, n65822, n65823,
    n65824, n65825, n65827, n65828, n65829, n65830, n65831, n65832, n65833,
    n65834, n65835, n65836, n65837, n65838, n65839, n65840, n65841, n65842,
    n65843, n65844, n65845, n65846, n65847, n65848, n65849, n65850, n65851,
    n65852, n65853, n65854, n65855, n65856, n65857, n65858, n65859, n65860,
    n65861, n65862, n65863, n65864, n65865, n65866, n65867, n65868, n65869,
    n65870, n65871, n65872, n65873, n65875, n65876, n65877, n65878, n65879,
    n65880, n65881, n65882, n65883, n65884, n65885, n65886, n65887, n65888,
    n65889, n65890, n65891, n65892, n65893, n65894, n65895, n65896, n65897,
    n65898, n65899, n65900, n65901, n65902, n65903, n65904, n65905, n65906,
    n65907, n65908, n65909, n65910, n65911, n65912, n65913, n65914, n65915,
    n65916, n65917, n65918, n65919, n65920, n65921, n65922, n65924, n65925,
    n65926, n65927, n65928, n65929, n65930, n65931, n65932, n65933, n65934,
    n65935, n65936, n65937, n65938, n65939, n65940, n65941, n65942, n65943,
    n65944, n65945, n65946, n65947, n65948, n65949, n65950, n65951, n65952,
    n65953, n65954, n65955, n65956, n65957, n65958, n65959, n65960, n65961,
    n65962, n65963, n65964, n65965, n65966, n65967, n65968, n65969, n65970,
    n65972, n65973, n65974, n65975, n65976, n65977, n65978, n65979, n65980,
    n65981, n65982, n65983, n65984, n65985, n65986, n65987, n65988, n65989,
    n65990, n65991, n65992, n65993, n65994, n65995, n65996, n65997, n65998,
    n65999, n66000, n66001, n66002, n66003, n66004, n66005, n66006, n66007,
    n66008, n66009, n66010, n66011, n66012, n66013, n66014, n66015, n66016,
    n66017, n66018, n66019, n66021, n66022, n66023, n66024, n66025, n66026,
    n66027, n66028, n66029, n66030, n66031, n66032, n66033, n66034, n66035,
    n66036, n66037, n66038, n66039, n66040, n66041, n66042, n66043, n66044,
    n66045, n66046, n66047, n66048, n66049, n66050, n66051, n66052, n66053,
    n66054, n66055, n66056, n66057, n66058, n66059, n66060, n66061, n66062,
    n66063, n66064, n66065, n66066, n66067, n66069, n66070, n66071, n66072,
    n66073, n66074, n66075, n66076, n66078, n66079, n66080, n66081, n66082,
    n66083, n66084, n66085, n66087, n66088, n66089, n66090, n66091, n66092,
    n66093, n66095, n66096, n66097, n66098, n66099, n66100, n66101, n66102,
    n66104, n66105, n66106, n66107, n66108, n66109, n66110, n66111, n66112,
    n66114, n66115, n66116, n66117, n66118, n66119, n66120, n66121, n66123,
    n66124, n66125, n66126, n66127, n66128, n66129, n66130, n66131, n66133,
    n66134, n66135, n66136, n66137, n66138, n66139, n66140, n66142, n66143,
    n66144, n66145, n66146, n66147, n66148, n66149, n66150, n66152, n66153,
    n66154, n66155, n66156, n66157, n66158, n66159, n66161, n66162, n66163,
    n66164, n66165, n66166, n66167, n66168, n66169, n66171, n66172, n66173,
    n66174, n66175, n66176, n66177, n66178, n66180, n66181, n66182, n66183,
    n66184, n66185, n66186, n66187, n66188, n66190, n66191, n66192, n66193,
    n66194, n66195, n66196, n66197, n66199, n66200, n66201, n66202, n66203,
    n66204, n66205, n66206, n66207, n66209, n66210, n66211, n66212, n66213,
    n66214, n66215, n66216, n66218, n66219, n66220, n66221, n66222, n66223,
    n66224, n66225, n66226, n66228, n66229, n66230, n66231, n66232, n66233,
    n66234, n66235, n66237, n66238, n66239, n66240, n66241, n66242, n66243,
    n66244, n66245, n66247, n66248, n66249, n66250, n66251, n66252, n66253,
    n66254, n66256, n66257, n66258, n66259, n66260, n66261, n66262, n66263,
    n66264, n66266, n66267, n66268, n66269, n66270, n66271, n66272, n66273,
    n66275, n66276, n66277, n66278, n66279, n66280, n66281, n66282, n66283,
    n66285, n66286, n66287, n66288, n66289, n66290, n66291, n66292, n66294,
    n66295, n66296, n66297, n66298, n66299, n66300, n66301, n66302, n66304,
    n66305, n66306, n66307, n66308, n66309, n66310, n66311, n66313, n66314,
    n66315, n66316, n66317, n66318, n66319, n66320, n66321, n66323, n66324,
    n66325, n66326, n66327, n66328, n66329, n66330, n66332, n66333, n66334,
    n66335, n66336, n66337, n66338, n66339, n66340, n66342, n66343, n66344,
    n66345, n66346, n66347, n66348, n66349, n66351, n66352, n66353, n66354,
    n66355, n66356, n66357, n66358, n66359, n66361, n66362, n66363, n66364,
    n66365, n66366, n66367, n66368, n66370, n66371, n66372, n66373, n66374,
    n66375, n66377, n66378, n66379, n66380, n66381, n66382, n66383, n66384,
    n66385, n66386, n66387, n66388, n66389, n66390, n66391, n66392, n66393,
    n66394, n66395, n66396, n66397, n66398, n66399, n66400, n66401, n66402,
    n66403, n66404, n66405, n66406, n66407, n66408, n66409, n66410, n66411,
    n66412, n66413, n66414, n66415, n66416, n66417, n66418, n66420, n66421,
    n66422, n66423, n66424, n66425, n66426, n66427, n66428, n66429, n66430,
    n66431, n66432, n66433, n66434, n66435, n66436, n66437, n66438, n66439,
    n66440, n66441, n66443, n66444, n66445, n66446, n66447, n66448, n66449,
    n66450, n66451, n66452, n66453, n66454, n66455, n66456, n66457, n66458,
    n66459, n66460, n66461, n66462, n66463, n66464, n66465, n66466, n66467,
    n66468, n66469, n66470, n66471, n66473, n66474, n66475, n66476, n66477,
    n66478, n66479, n66480, n66481, n66482, n66483, n66484, n66485, n66486,
    n66487, n66488, n66489, n66490, n66491, n66492, n66493, n66494, n66495,
    n66496, n66497, n66498, n66499, n66500, n66501, n66502, n66504, n66505,
    n66506, n66507, n66508, n66509, n66510, n66511, n66512, n66513, n66514,
    n66515, n66516, n66517, n66518, n66519, n66520, n66521, n66522, n66523,
    n66524, n66525, n66526, n66527, n66528, n66529, n66530, n66531, n66532,
    n66533, n66534, n66535, n66536, n66537, n66538, n66539, n66541, n66542,
    n66543, n66544, n66545, n66546, n66547, n66548, n66549, n66550, n66551,
    n66552, n66553, n66554, n66555, n66556, n66557, n66558, n66559, n66560,
    n66561, n66562, n66563, n66564, n66565, n66566, n66567, n66568, n66569,
    n66570, n66572, n66573, n66574, n66575, n66576, n66577, n66578, n66579,
    n66580, n66581, n66582, n66583, n66584, n66585, n66586, n66587, n66588,
    n66589, n66590, n66591, n66592, n66593, n66594, n66595, n66596, n66597,
    n66598, n66600, n66601, n66602, n66603, n66604, n66605, n66606, n66607,
    n66608, n66609, n66610, n66611, n66612, n66613, n66614, n66615, n66616,
    n66617, n66618, n66619, n66620, n66621, n66622, n66623, n66624, n66626,
    n66627, n66628, n66629, n66630, n66631, n66632, n66633, n66634, n66635,
    n66636, n66637, n66638, n66639, n66640, n66641, n66642, n66643, n66644,
    n66645, n66646, n66647, n66648, n66649, n66650, n66651, n66652, n66654,
    n66655, n66656, n66657, n66658, n66659, n66660, n66661, n66662, n66663,
    n66664, n66665, n66666, n66667, n66668, n66669, n66670, n66671, n66672,
    n66673, n66674, n66675, n66676, n66677, n66678, n66680, n66681, n66682,
    n66683, n66684, n66685, n66686, n66687, n66688, n66689, n66690, n66691,
    n66692, n66693, n66694, n66695, n66696, n66697, n66698, n66699, n66700,
    n66701, n66702, n66703, n66704, n66705, n66706, n66708, n66709, n66710,
    n66711, n66712, n66713, n66714, n66715, n66716, n66717, n66718, n66719,
    n66720, n66721, n66722, n66723, n66724, n66725, n66726, n66727, n66728,
    n66729, n66730, n66731, n66732, n66734, n66735, n66736, n66737, n66738,
    n66739, n66740, n66741, n66742, n66743, n66744, n66745, n66746, n66747,
    n66748, n66749, n66750, n66751, n66752, n66753, n66754, n66755, n66756,
    n66757, n66758, n66759, n66760, n66762, n66763, n66764, n66765, n66766,
    n66767, n66768, n66769, n66770, n66771, n66772, n66773, n66774, n66775,
    n66776, n66777, n66778, n66779, n66780, n66781, n66782, n66783, n66784,
    n66785, n66786, n66788, n66789, n66790, n66791, n66792, n66793, n66794,
    n66795, n66796, n66797, n66798, n66799, n66800, n66801, n66802, n66803,
    n66804, n66805, n66806, n66807, n66808, n66809, n66810, n66811, n66812,
    n66813, n66814, n66816, n66817, n66818, n66819, n66820, n66821, n66822,
    n66823, n66824, n66825, n66826, n66827, n66828, n66829, n66830, n66831,
    n66832, n66833, n66834, n66835, n66836, n66837, n66838, n66839, n66840,
    n66842, n66843, n66844, n66845, n66846, n66847, n66848, n66849, n66850,
    n66851, n66852, n66853, n66854, n66855, n66856, n66857, n66858, n66859,
    n66860, n66861, n66862, n66863, n66864, n66865, n66866, n66867, n66868,
    n66870, n66871, n66872, n66873, n66874, n66875, n66876, n66877, n66878,
    n66879, n66880, n66881, n66882, n66883, n66884, n66885, n66886, n66887,
    n66888, n66889, n66890, n66891, n66892, n66893, n66894, n66896, n66897,
    n66898, n66899, n66900, n66901, n66902, n66903, n66904, n66905, n66906,
    n66907, n66908, n66909, n66910, n66911, n66912, n66913, n66914, n66915,
    n66916, n66917, n66918, n66919, n66920, n66921, n66922, n66924, n66925,
    n66926, n66927, n66928, n66929, n66930, n66931, n66932, n66933, n66934,
    n66935, n66936, n66937, n66938, n66939, n66940, n66941, n66942, n66943,
    n66944, n66945, n66946, n66947, n66948, n66950, n66951, n66952, n66953,
    n66954, n66955, n66956, n66957, n66958, n66959, n66960, n66961, n66962,
    n66963, n66964, n66965, n66966, n66967, n66968, n66969, n66970, n66971,
    n66972, n66973, n66974, n66975, n66977, n66978, n66979, n66980, n66981,
    n66982, n66983, n66984, n66985, n66986, n66987, n66988, n66989, n66990,
    n66991, n66992, n66993, n66994, n66995, n66996, n66997, n66998, n66999,
    n67000, n67002, n67003, n67004, n67005, n67006, n67007, n67008, n67009,
    n67010, n67011, n67012, n67013, n67014, n67015, n67016, n67017, n67018,
    n67019, n67020, n67021, n67022, n67023, n67024, n67025, n67026, n67027,
    n67029, n67030, n67031, n67032, n67033, n67034, n67035, n67036, n67037,
    n67038, n67039, n67040, n67041, n67042, n67043, n67044, n67045, n67046,
    n67047, n67048, n67049, n67050, n67051, n67052, n67054, n67055, n67056,
    n67057, n67058, n67059, n67060, n67061, n67062, n67063, n67064, n67065,
    n67066, n67067, n67068, n67069, n67070, n67071, n67072, n67073, n67074,
    n67075, n67076, n67077, n67078, n67079, n67081, n67082, n67083, n67084,
    n67085, n67086, n67087, n67088, n67089, n67090, n67091, n67092, n67093,
    n67094, n67095, n67096, n67097, n67098, n67099, n67100, n67101, n67102,
    n67103, n67104, n67106, n67107, n67108, n67109, n67110, n67111, n67112,
    n67113, n67114, n67115, n67116, n67117, n67118, n67119, n67120, n67121,
    n67122, n67123, n67124, n67125, n67126, n67127, n67128, n67129, n67130,
    n67131, n67133, n67134, n67135, n67136, n67137, n67138, n67139, n67140,
    n67141, n67142, n67143, n67144, n67145, n67146, n67147, n67148, n67149,
    n67150, n67151, n67152, n67153, n67154, n67155, n67156, n67158, n67159,
    n67160, n67161, n67162, n67163, n67164, n67165, n67166, n67167, n67168,
    n67169, n67170, n67171, n67172, n67173, n67174, n67175, n67176, n67177,
    n67178, n67179, n67180, n67181, n67182, n67183, n67185, n67186, n67187,
    n67188, n67189, n67190, n67191, n67192, n67193, n67194, n67195, n67196,
    n67197, n67198, n67199, n67200, n67201, n67202, n67203, n67204, n67205,
    n67206, n67207, n67208, n67210, n67211, n67212, n67213, n67214, n67215,
    n67216, n67217, n67218, n67219, n67220, n67221, n67222, n67223, n67224,
    n67225, n67226, n67227, n67228, n67229, n67230, n67231, n67232, n67233,
    n67235, n67236, n67237, n67238, n67239, n67240, n67241, n67242, n67243,
    n67244, n67245, n67246, n67247, n67248, n67249, n67250, n67251, n67252,
    n67253, n67254, n67255, n67256, n67257, n67258, n67259, n67260, n67262,
    n67263, n67264, n67265, n67266, n67267, n67268, n67269, n67270, n67271,
    n67272, n67273, n67274, n67275, n67276, n67277, n67278, n67279, n67280,
    n67281, n67282, n67283, n67284, n67285, n67286, n67287, n67288, n67289,
    n67290, n67291, n67292, n67293, n67294, n67295, n67296, n67297, n67298,
    n67299, n67301, n67302, n67303, n67304, n67305, n67306, n67307, n67308,
    n67310, n67311, n67312, n67314, n67315, n67316, n67318, n67319, n67321,
    n67322, n67323, n67325, n67326, n67328, n67329, n67330, n67331, n67333,
    n67334, n67335, n67336, n67337, n67338, n67339, n67340, n67341, n67342,
    n67343, n67344, n67345, n67346, n67347, n67349, n67350, n67351, n67353,
    n67354, n67356, n67357, n67358, n67360, n67362, n67363, n67364, n67365,
    n67366, n67368, n67369, n67370, n67372, n67373, n67374, n67376, n67377,
    n67379, n67380, n67382, n67383, n67385, n67386, n67387, n67388, n67389,
    n67390, n67392, n67393, n67394, n67395, n67397, n67398, n67399, n67400,
    n67402, n67403, n67404, n67405, n67407, n67408, n67409, n67410, n67412,
    n67413, n67414, n67415, n67417, n67418, n67419, n67420, n67422, n67423,
    n67424, n67425, n67427, n67428, n67429, n67430, n67432, n67433, n67434,
    n67435, n67437, n67438, n67439, n67440, n67442, n67443, n67444, n67445,
    n67447, n67448, n67449, n67450, n67452, n67453, n67454, n67455, n67457,
    n67458, n67459, n67460, n67462, n67463, n67464, n67465, n67467, n67468,
    n67469, n67470, n67472, n67473, n67474, n67475, n67477, n67478, n67479,
    n67480, n67482, n67483, n67484, n67485, n67487, n67488, n67489, n67490,
    n67492, n67493, n67494, n67495, n67497, n67498, n67499, n67500, n67502,
    n67503, n67504, n67505, n67507, n67508, n67509, n67510, n67512, n67513,
    n67514, n67515, n67517, n67518, n67519, n67520, n67522, n67523, n67524,
    n67525, n67527, n67528, n67529, n67530, n67532, n67533, n67534, n67535,
    n67537, n67538, n67539, n67540, n67541, n67542, n67543, n67544, n67545,
    n67546, n67547, n67548, n67549, n67550, n67551, n67552, n67553, n67554,
    n67555, n67556, n67557, n67558, n67559, n67560, n67562, n67563, n67564,
    n67565, n67566, n67567, n67568, n67569, n67570, n67571, n67572, n67573,
    n67574, n67576, n67577, n67578, n67579, n67580, n67581, n67582, n67583,
    n67584, n67586, n67587, n67588, n67589, n67590, n67591, n67593, n67594,
    n67626, n67627, n67628, n67629, n67630, n67631, n67632, n67633, n67634,
    n67635, n67636, n67637, n67638, n67639, n67640, n67641, n67642, n67643,
    n67644, n67645, n67646, n67647, n67648, n67649, n67650, n67651, n67652,
    n67653, n67654, n67655, n67656, n67657, n67658, n67659, n67660, n67661,
    n67662, n67663, n67664, n67665, n67666, n67667, n67668, n67669, n67670,
    n67671, n67672, n67673, n67674, n67675, n67676, n67677, n67678, n67679,
    n67680, n67681, n67682, n67683, n67684, n67685, n67686, n67687, n67688,
    n67689, n67690, n67691, n67692, n67693, n67694, n67695, n67696, n67697,
    n67698, n67699, n67700, n67701, n67702, n67703, n67704, n67705, n67706,
    n67707, n67708, n67709, n67710, n67711, n67712, n67713, n67714, n67715,
    n67716, n67717, n67718, n67719, n67720, n67721, n67722, n67723, n67724,
    n67725, n67726, n67727, n67728, n67729, n67730, n67731, n67732, n67733,
    n67734, n67735, n67736, n67737, n67738, n67739, n67740, n67741, n67742,
    n67743, n67744, n67745, n67746, n67747, n67748, n67749, n67750, n67751,
    n67752, n67753, n67754, n67755, n67756, n67757, n67758, n67759, n67760,
    n67761, n67762, n67763, n67764, n67765, n67766, n67767, n67768, n67769,
    n67770, n67771, n67772, n67773, n67774, n67775, n67776, n67777, n67778,
    n67779, n67780, n67781, n67782, n67783, n67784, n67785, n67786, n67787,
    n67788, n67789, n67790, n67791, n67792, n67793, n67794, n67795, n67796,
    n67797, n67798, n67799, n67800, n67801, n67802, n67803, n67804, n67805,
    n67806, n67807, n67808, n67809, n67810, n67811, n67812, n67813, n67814,
    n67815, n67816, n67817, n67818, n67819, n67820, n67821, n67822, n67823,
    n67824, n67825, n67826, n67827, n67828, n67829, n67830, n67831, n67832,
    n67833, n67834, n67835, n67836, n67837, n67838, n67839, n67840, n67841,
    n67842, n67843, n67844, n67845, n67846, n67847, n67848, n67849, n67850,
    n67851, n67852, n67853, n67854, n67855, n67856, n67857, n67858, n67859,
    n67860, n67861, n67862, n67863, n67864, n67865, n67866, n67867, n67868,
    n67869, n67870, n67871, n67872, n67873, n67874, n67875, n67876, n67877,
    n67878, n67879, n67880, n67881, n67882, n67883, n67884, n67885, n67886,
    n67887, n67888, n67889, n67890, n67891, n67892, n67893, n67894, n67895,
    n67896, n67897, n67898, n67899, n67900, n67901, n67902, n67903, n67904,
    n67905, n67906, n67907, n67908, n67909, n67910, n67911, n67912, n67913,
    n67914, n67915, n67916, n67917, n67918, n67919, n67920, n67921, n67922,
    n67923, n67924, n67925, n67926, n67927, n67928, n67929, n67930, n67931,
    n67932, n67933, n67934, n67935, n67936, n67937, n67938, n67939, n67940,
    n67941, n67942, n67943, n67944, n67945, n67946, n67947, n67948, n67949,
    n67950, n67951, n67952, n67953, n67954, n67955, n67956, n67957, n67958,
    n67959, n67960, n67961, n67962, n67963, n67964, n67965, n67966, n67967,
    n67968, n67969, n67970, n67971, n67972, n67973, n67974, n67975, n67976,
    n67977, n67978, n67979, n67980, n67981, n67982, n67983, n67984, n67985,
    n67986, n67987, n67988, n67989, n67990, n67991, n67992, n67993, n67994,
    n67995, n67996, n67997, n67998, n67999, n68000, n68001, n68002, n68003,
    n68004, n68005, n68006, n68007, n68008, n68009, n68010, n68011, n68012,
    n68013, n68014, n68015, n68016, n68017, n68018, n68019, n68020, n68021,
    n68022, n68023, n68024, n68025, n68026, n68027, n68028, n68029, n68030,
    n68031, n68032, n68033, n68034, n68035, n68036, n68037, n68038, n68039,
    n68040, n68041, n68042, n68043, n68044, n68045, n68046, n68047, n68048,
    n68049, n68050, n68051, n68052, n68053, n68054, n68055, n68056, n68057,
    n68058, n68059, n68060, n68061, n68062, n68063, n68064, n68065, n68066,
    n68067, n68068, n68069, n68070, n68071, n68072, n68073, n68074, n68075,
    n68076, n68077, n68078, n68079, n68080, n68081, n68082, n68083, n68084,
    n68085, n68086, n68087, n68088, n68089, n68090, n68091, n68092, n68093,
    n68094, n68095, n68096, n68097, n68098, n68099, n68100, n68101, n68102,
    n68103, n68104, n68105, n68106, n68107, n68108, n68109, n68110, n68111,
    n68112, n68113, n68114, n68115, n68116, n68117, n68118, n68119, n68120,
    n68121, n68122, n68123, n68124, n68125, n68126, n68127, n68128, n68129,
    n68130, n68131, n68132, n68133, n68134, n68135, n68136, n68137, n68138,
    n68139, n68140, n68141, n68142, n68143, n68144, n68145, n68146, n68147,
    n68148, n68149, n68150, n68151, n68152, n68153, n68154, n68155, n68156,
    n68157, n68158, n68159, n68160, n68161, n68162, n68163, n68164, n68165,
    n68166, n68167, n68168, n68169, n68170, n68171, n68172, n68173, n68174,
    n68175, n68176, n68177, n68178, n68179, n68180, n68181, n68182, n68183,
    n68184, n68185, n68186, n68187, n68188, n68189, n68190, n68191, n68192,
    n68193, n68194, n68195, n68196, n68197, n68198, n68199, n68200, n68201,
    n68202, n68203, n68204, n68205, n68206, n68207, n68208, n68209, n68210,
    n68211, n68212, n68213, n68214, n68215, n68216, n68217, n68218, n68219,
    n68220, n68221, n68222, n68223, n68224, n68225, n68226, n68227, n68228,
    n68229, n68230, n68231, n68232, n68233, n68234, n68235, n68236, n68237,
    n68238, n68239, n68240, n68241, n68242, n68243, n68244, n68245, n68246,
    n68247, n68248, n68249, n68250, n68251, n68252, n68253, n68254, n68255,
    n68256, n68257, n68259, n68260, n68261, n68262, n68263, n68264, n68265,
    n68266, n68268, n68269, n68270, n68271, n68272, n68273, n68274, n68275,
    n68276, n68277, n68278, n68279, n68280, n68281, n68283, n68284, n68285,
    n68286, n68287, n68288, n68289, n68290, n68291, n68292, n68293, n68294,
    n68295, n68296, n68297, n68298, n68299, n68300, n68301, n68302, n68303,
    n68304, n68305, n68306, n68307, n68308, n68309, n68310, n68311, n68312,
    n68313, n68314, n68315, n68316, n68317, n68318, n68319, n68320, n68321,
    n68322, n68324, n68325, n68326, n68327, n68328, n68329, n68330, n68331,
    n68332, n68333, n68334, n68335, n68336, n68337, n68338, n68339, n68340,
    n68341, n68342, n68343, n68344, n68345, n68346, n68347, n68348, n68349,
    n68350, n68351, n68352, n68353, n68354, n68355, n68356, n68357, n68358,
    n68359, n68360, n68361, n68362, n68363, n68364, n68365, n68366, n68367,
    n68368, n68369, n68370, n68371, n68372, n68373, n68374, n68375, n68376,
    n68377, n68378, n68379, n68380, n68381, n68382, n68383, n68384, n68385,
    n68386, n68387, n68388, n68389, n68390, n68391, n68392, n68393, n68394,
    n68395, n68396, n68397, n68398, n68399, n68400, n68401, n68402, n68403,
    n68404, n68405, n68406, n68407, n68408, n68410, n68411, n68412, n68413,
    n68414, n68415, n68416, n68417, n68418, n68419, n68420, n68421, n68422,
    n68423, n68424, n68425, n68426, n68427, n68428, n68429, n68430, n68432,
    n68433, n68434, n68435, n68436, n68437, n68438, n68439, n68440, n68441,
    n68442, n68443, n68444, n68445, n68446, n68447, n68448, n68449, n68450,
    n68451, n68452, n68454, n68455, n68456, n68457, n68458, n68459, n68460,
    n68461, n68462, n68463, n68464, n68465, n68466, n68467, n68468, n68469,
    n68470, n68471, n68472, n68473, n68474, n68476, n68477, n68478, n68479,
    n68480, n68481, n68482, n68483, n68484, n68485, n68486, n68487, n68488,
    n68489, n68490, n68491, n68492, n68493, n68494, n68495, n68496, n68498,
    n68499, n68500, n68501, n68502, n68503, n68504, n68505, n68506, n68507,
    n68508, n68509, n68510, n68511, n68512, n68513, n68514, n68515, n68516,
    n68517, n68518, n68520, n68521, n68522, n68523, n68524, n68525, n68526,
    n68527, n68528, n68529, n68530, n68531, n68532, n68533, n68534, n68535,
    n68536, n68537, n68538, n68539, n68540, n68542, n68543, n68544, n68545,
    n68546, n68547, n68548, n68549, n68550, n68551, n68552, n68553, n68554,
    n68555, n68556, n68557, n68558, n68559, n68560, n68561, n68562, n68564,
    n68565, n68566, n68567, n68568, n68569, n68570, n68571, n68572, n68573,
    n68574, n68575, n68576, n68577, n68578, n68579, n68580, n68581, n68582,
    n68583, n68584, n68585, n68586, n68587, n68588, n68590, n68591, n68592,
    n68593, n68594, n68595, n68596, n68597, n68599, n68600, n68601, n68602,
    n68603, n68604, n68605, n68606, n68608, n68609, n68610, n68611, n68612,
    n68613, n68614, n68615, n68617, n68618, n68619, n68620, n68621, n68622,
    n68623, n68624, n68626, n68627, n68628, n68629, n68630, n68631, n68632,
    n68633, n68635, n68636, n68637, n68638, n68639, n68640, n68641, n68642,
    n68644, n68645, n68646, n68647, n68648, n68649, n68650, n68651, n68653,
    n68654, n68655, n68656, n68657, n68658, n68659, n68660, n68661, n68662,
    n68663, n68664, n68665, n68666, n68667, n68668, n68669, n68670, n68671,
    n68672, n68673, n68674, n68675, n68676, n68678, n68679, n68680, n68681,
    n68682, n68683, n68684, n68685, n68687, n68688, n68689, n68690, n68691,
    n68692, n68693, n68694, n68696, n68697, n68698, n68699, n68700, n68701,
    n68702, n68703, n68705, n68706, n68707, n68708, n68709, n68710, n68711,
    n68712, n68714, n68715, n68716, n68717, n68718, n68719, n68720, n68721,
    n68723, n68724, n68725, n68726, n68727, n68728, n68729, n68730, n68732,
    n68733, n68734, n68735, n68736, n68737, n68738, n68739, n68741, n68742,
    n68743, n68744, n68745, n68746, n68747, n68748, n68749, n68750, n68751,
    n68752, n68753, n68754, n68755, n68756, n68757, n68758, n68759, n68760,
    n68761, n68762, n68763, n68764, n68766, n68767, n68768, n68769, n68770,
    n68771, n68772, n68773, n68775, n68776, n68777, n68778, n68779, n68780,
    n68781, n68782, n68784, n68785, n68786, n68787, n68788, n68789, n68790,
    n68791, n68793, n68794, n68795, n68796, n68797, n68798, n68799, n68800,
    n68802, n68803, n68804, n68805, n68806, n68807, n68808, n68809, n68811,
    n68812, n68813, n68814, n68815, n68816, n68817, n68818, n68820, n68821,
    n68822, n68823, n68824, n68825, n68826, n68827, n68829, n68830, n68831,
    n68832, n68833, n68834, n68835, n68836, n68837, n68838, n68839, n68840,
    n68841, n68842, n68843, n68844, n68845, n68846, n68847, n68848, n68849,
    n68850, n68851, n68852, n68853, n68855, n68856, n68857, n68858, n68859,
    n68860, n68861, n68862, n68864, n68865, n68866, n68867, n68868, n68869,
    n68870, n68871, n68873, n68874, n68875, n68876, n68877, n68878, n68879,
    n68880, n68882, n68883, n68884, n68885, n68886, n68887, n68888, n68889,
    n68891, n68892, n68893, n68894, n68895, n68896, n68897, n68898, n68900,
    n68901, n68902, n68903, n68904, n68905, n68906, n68907, n68909, n68910,
    n68911, n68912, n68913, n68914, n68915, n68916, n68918, n68919, n68920,
    n68921, n68922, n68923, n68924, n68925, n68926, n68927, n68928, n68929,
    n68930, n68931, n68932, n68933, n68934, n68935, n68936, n68937, n68938,
    n68939, n68940, n68942, n68943, n68944, n68945, n68946, n68947, n68948,
    n68949, n68951, n68952, n68953, n68954, n68955, n68956, n68957, n68958,
    n68960, n68961, n68962, n68963, n68964, n68965, n68966, n68967, n68969,
    n68970, n68971, n68972, n68973, n68974, n68975, n68976, n68978, n68979,
    n68980, n68981, n68982, n68983, n68984, n68985, n68987, n68988, n68989,
    n68990, n68991, n68992, n68993, n68994, n68996, n68997, n68998, n68999,
    n69000, n69001, n69002, n69003, n69005, n69006, n69007, n69008, n69009,
    n69010, n69011, n69012, n69013, n69014, n69015, n69016, n69017, n69018,
    n69019, n69020, n69021, n69022, n69023, n69024, n69025, n69026, n69028,
    n69029, n69030, n69031, n69032, n69033, n69034, n69035, n69037, n69038,
    n69039, n69040, n69041, n69042, n69043, n69044, n69046, n69047, n69048,
    n69049, n69050, n69051, n69052, n69053, n69055, n69056, n69057, n69058,
    n69059, n69060, n69061, n69062, n69064, n69065, n69066, n69067, n69068,
    n69069, n69070, n69071, n69073, n69074, n69075, n69076, n69077, n69078,
    n69079, n69080, n69082, n69083, n69084, n69085, n69086, n69087, n69088,
    n69089, n69091, n69092, n69093, n69094, n69095, n69096, n69097, n69098,
    n69099, n69100, n69101, n69102, n69103, n69104, n69105, n69106, n69107,
    n69108, n69109, n69110, n69111, n69113, n69114, n69115, n69116, n69117,
    n69118, n69119, n69120, n69122, n69123, n69124, n69125, n69126, n69127,
    n69128, n69129, n69131, n69132, n69133, n69134, n69135, n69136, n69137,
    n69138, n69140, n69141, n69142, n69143, n69144, n69145, n69146, n69147,
    n69149, n69150, n69151, n69152, n69153, n69154, n69155, n69156, n69158,
    n69159, n69160, n69161, n69162, n69163, n69164, n69165, n69167, n69168,
    n69169, n69170, n69171, n69172, n69173, n69174, n69176, n69177, n69178,
    n69179, n69180, n69181, n69182, n69183, n69184, n69185, n69186, n69187,
    n69188, n69189, n69190, n69191, n69192, n69193, n69194, n69195, n69197,
    n69198, n69199, n69200, n69201, n69202, n69203, n69204, n69206, n69207,
    n69208, n69209, n69210, n69211, n69212, n69213, n69215, n69216, n69217,
    n69218, n69219, n69220, n69221, n69222, n69224, n69225, n69226, n69227,
    n69228, n69229, n69230, n69231, n69233, n69234, n69235, n69236, n69237,
    n69238, n69239, n69240, n69242, n69243, n69244, n69245, n69246, n69247,
    n69248, n69249, n69251, n69252, n69253, n69254, n69255, n69256, n69257,
    n69258, n69260, n69261, n69262, n69263, n69264, n69265, n69266, n69267,
    n69268, n69269, n69270, n69271, n69272, n69273, n69274, n69275, n69276,
    n69277, n69278, n69279, n69280, n69281, n69282, n69284, n69285, n69286,
    n69287, n69288, n69289, n69290, n69291, n69293, n69294, n69295, n69296,
    n69297, n69298, n69299, n69300, n69302, n69303, n69304, n69305, n69306,
    n69307, n69308, n69309, n69311, n69312, n69313, n69314, n69315, n69316,
    n69317, n69318, n69320, n69321, n69322, n69323, n69324, n69325, n69326,
    n69327, n69329, n69330, n69331, n69332, n69333, n69334, n69335, n69336,
    n69338, n69339, n69340, n69341, n69342, n69343, n69344, n69345, n69347,
    n69348, n69349, n69350, n69351, n69352, n69353, n69354, n69355, n69356,
    n69357, n69358, n69359, n69360, n69361, n69362, n69363, n69364, n69365,
    n69366, n69367, n69368, n69369, n69371, n69372, n69373, n69374, n69375,
    n69376, n69377, n69378, n69380, n69381, n69382, n69383, n69384, n69385,
    n69386, n69387, n69389, n69390, n69391, n69392, n69393, n69394, n69395,
    n69396, n69398, n69399, n69400, n69401, n69402, n69403, n69404, n69405,
    n69407, n69408, n69409, n69410, n69411, n69412, n69413, n69414, n69416,
    n69417, n69418, n69419, n69420, n69421, n69422, n69423, n69425, n69426,
    n69427, n69428, n69429, n69430, n69431, n69432, n69434, n69435, n69436,
    n69437, n69438, n69439, n69440, n69441, n69442, n69443, n69444, n69445,
    n69446, n69447, n69448, n69449, n69450, n69451, n69452, n69453, n69454,
    n69456, n69457, n69458, n69459, n69460, n69461, n69462, n69463, n69465,
    n69466, n69467, n69468, n69469, n69470, n69471, n69472, n69474, n69475,
    n69476, n69477, n69478, n69479, n69480, n69481, n69483, n69484, n69485,
    n69486, n69487, n69488, n69489, n69490, n69492, n69493, n69494, n69495,
    n69496, n69497, n69498, n69499, n69501, n69502, n69503, n69504, n69505,
    n69506, n69507, n69508, n69510, n69511, n69512, n69513, n69514, n69515,
    n69516, n69517, n69519, n69520, n69521, n69522, n69523, n69524, n69525,
    n69526, n69527, n69528, n69529, n69530, n69531, n69532, n69533, n69534,
    n69535, n69536, n69537, n69538, n69539, n69540, n69541, n69542, n69544,
    n69545, n69546, n69547, n69548, n69549, n69550, n69551, n69553, n69554,
    n69555, n69556, n69557, n69558, n69559, n69560, n69562, n69563, n69564,
    n69565, n69566, n69567, n69568, n69569, n69571, n69572, n69573, n69574,
    n69575, n69576, n69577, n69578, n69580, n69581, n69582, n69583, n69584,
    n69585, n69586, n69587, n69589, n69590, n69591, n69592, n69593, n69594,
    n69595, n69596, n69598, n69599, n69600, n69601, n69602, n69603, n69604,
    n69605, n69607, n69608, n69609, n69610, n69611, n69612, n69613, n69614,
    n69615, n69616, n69617, n69618, n69619, n69620, n69621, n69622, n69623,
    n69624, n69625, n69626, n69628, n69629, n69630, n69631, n69632, n69633,
    n69634, n69635, n69637, n69638, n69639, n69640, n69641, n69642, n69643,
    n69644, n69646, n69647, n69648, n69649, n69650, n69651, n69652, n69653,
    n69655, n69656, n69657, n69658, n69659, n69660, n69661, n69662, n69664,
    n69665, n69666, n69667, n69668, n69669, n69670, n69671, n69673, n69674,
    n69675, n69676, n69677, n69678, n69679, n69680, n69682, n69683, n69684,
    n69685, n69686, n69687, n69688, n69689, n69691, n69692, n69693, n69694,
    n69695, n69696, n69697, n69698, n69699, n69700, n69701, n69702, n69703,
    n69704, n69705, n69706, n69707, n69708, n69709, n69710, n69712, n69713,
    n69714, n69715, n69716, n69717, n69718, n69719, n69721, n69722, n69723,
    n69724, n69725, n69726, n69727, n69728, n69730, n69731, n69732, n69733,
    n69734, n69735, n69736, n69737, n69739, n69740, n69741, n69742, n69743,
    n69744, n69745, n69746, n69748, n69749, n69750, n69751, n69752, n69753,
    n69754, n69755, n69757, n69758, n69759, n69760, n69761, n69762, n69763,
    n69764, n69766, n69767, n69768, n69769, n69770, n69771, n69772, n69773,
    n69775, n69776, n69777, n69778, n69779, n69780, n69781, n69782, n69783,
    n69784, n69785, n69786, n69787, n69788, n69789, n69790, n69791, n69792,
    n69793, n69795, n69796, n69797, n69798, n69799, n69800, n69801, n69802,
    n69804, n69805, n69806, n69807, n69808, n69809, n69810, n69811, n69813,
    n69814, n69815, n69816, n69817, n69818, n69819, n69820, n69822, n69823,
    n69824, n69825, n69826, n69827, n69828, n69829, n69831, n69832, n69833,
    n69834, n69835, n69836, n69837, n69838, n69840, n69841, n69842, n69843,
    n69844, n69845, n69846, n69847, n69849, n69850, n69851, n69852, n69853,
    n69854, n69855, n69856, n69858, n69859, n69860, n69861, n69862, n69863,
    n69864, n69865, n69866, n69867, n69869, n69870, n69871, n69872, n69873,
    n69874, n69876, n69877, n69878, n69879, n69880, n69881, n69882, n69883,
    n69885, n69886, n69887, n69888, n69889, n69890, n69891, n69893, n69894,
    n69895, n69896, n69897, n69898, n69899, n69901, n69902, n69903, n69904,
    n69906, n69907, n69908, n69909, n69910, n69911, n69912, n69913, n69914,
    n69915, n69916, n69917, n69918, n69920, n69921, n69922, n69923, n69924,
    n69925, n69926, n69927, n69928, n69929, n69930, n69931, n69932, n69934,
    n69935, n69936, n69937, n69938, n69939, n69940, n69941, n69942, n69943,
    n69944, n69945, n69947, n69948, n69949, n69950, n69951, n69953, n69954,
    n69955, n69956, n69957, n69958, n69959, n69960, n69961, n69962, n69963,
    n69964, n69965, n69966, n69967, n69968, n69969, n69970, n69971, n69972,
    n69973, n69974, n69975, n69976, n69977, n69978, n69979, n69980, n69981,
    n69982, n69983, n69984, n69985, n69986, n69987, n69988, n69989, n69990,
    n69991, n69992, n69993, n69994, n69995, n69996, n69997, n69998, n69999,
    n70000, n70001, n70002, n70003, n70004, n70005, n70006, n70007, n70008,
    n70009, n70010, n70011, n70012, n70013, n70014, n70015, n70016, n70017,
    n70018, n70019, n70020, n70021, n70022, n70023, n70024, n70025, n70026,
    n70027, n70028, n70029, n70030, n70031, n70032, n70033, n70034, n70035,
    n70036, n70037, n70038, n70039, n70040, n70041, n70042, n70043, n70044,
    n70045, n70046, n70047, n70048, n70049, n70050, n70051, n70052, n70053,
    n70054, n70055, n70056, n70057, n70058, n70059, n70060, n70061, n70062,
    n70063, n70064, n70065, n70066, n70067, n70068, n70069, n70070, n70071,
    n70072, n70073, n70074, n70075, n70076, n70077, n70078, n70079, n70080,
    n70081, n70082, n70083, n70084, n70085, n70086, n70087, n70088, n70089,
    n70090, n70091, n70092, n70093, n70094, n70095, n70096, n70097, n70098,
    n70099, n70100, n70101, n70102, n70103, n70104, n70105, n70106, n70107,
    n70108, n70109, n70110, n70111, n70112, n70113, n70114, n70115, n70116,
    n70117, n70118, n70119, n70120, n70121, n70122, n70123, n70124, n70125,
    n70126, n70127, n70129, n70130, n70131, n70132, n70133, n70134, n70135,
    n70136, n70137, n70138, n70139, n70140, n70141, n70142, n70143, n70144,
    n70145, n70146, n70147, n70148, n70149, n70150, n70151, n70152, n70153,
    n70154, n70155, n70156, n70157, n70158, n70159, n70160, n70161, n70162,
    n70163, n70164, n70165, n70166, n70167, n70168, n70169, n70170, n70171,
    n70172, n70173, n70174, n70175, n70176, n70177, n70178, n70179, n70180,
    n70181, n70182, n70183, n70184, n70185, n70186, n70187, n70188, n70189,
    n70190, n70191, n70192, n70193, n70194, n70195, n70196, n70197, n70198,
    n70199, n70200, n70201, n70202, n70203, n70204, n70205, n70206, n70207,
    n70208, n70209, n70210, n70211, n70212, n70213, n70214, n70215, n70216,
    n70217, n70218, n70219, n70220, n70221, n70222, n70223, n70224, n70225,
    n70226, n70227, n70228, n70229, n70230, n70231, n70232, n70233, n70234,
    n70235, n70237, n70238, n70239, n70240, n70241, n70242, n70243, n70244,
    n70245, n70246, n70247, n70248, n70249, n70250, n70251, n70252, n70253,
    n70254, n70255, n70256, n70257, n70258, n70259, n70260, n70261, n70262,
    n70263, n70264, n70265, n70266, n70267, n70268, n70269, n70270, n70271,
    n70272, n70273, n70274, n70275, n70276, n70277, n70278, n70279, n70280,
    n70281, n70282, n70283, n70284, n70285, n70286, n70287, n70288, n70289,
    n70290, n70291, n70292, n70293, n70294, n70295, n70296, n70297, n70298,
    n70299, n70300, n70301, n70302, n70303, n70304, n70305, n70306, n70307,
    n70308, n70309, n70310, n70311, n70312, n70313, n70314, n70315, n70316,
    n70317, n70318, n70319, n70320, n70321, n70322, n70323, n70324, n70325,
    n70326, n70327, n70328, n70329, n70330, n70331, n70332, n70333, n70334,
    n70335, n70336, n70337, n70338, n70339, n70340, n70341, n70342, n70343,
    n70344, n70345, n70346, n70347, n70348, n70349, n70350, n70351, n70352,
    n70353, n70354, n70355, n70356, n70358, n70359, n70360, n70361, n70362,
    n70363, n70364, n70365, n70366, n70367, n70368, n70369, n70370, n70371,
    n70372, n70373, n70374, n70375, n70376, n70377, n70378, n70379, n70380,
    n70381, n70382, n70383, n70384, n70385, n70386, n70387, n70388, n70389,
    n70390, n70391, n70392, n70393, n70394, n70395, n70396, n70397, n70398,
    n70399, n70400, n70401, n70402, n70403, n70404, n70405, n70406, n70407,
    n70408, n70409, n70410, n70411, n70412, n70413, n70414, n70415, n70416,
    n70417, n70418, n70419, n70420, n70421, n70422, n70423, n70424, n70425,
    n70426, n70427, n70428, n70429, n70430, n70431, n70432, n70433, n70434,
    n70435, n70436, n70437, n70438, n70439, n70440, n70441, n70442, n70443,
    n70444, n70445, n70446, n70447, n70448, n70449, n70450, n70451, n70452,
    n70453, n70454, n70455, n70456, n70457, n70458, n70459, n70460, n70461,
    n70462, n70463, n70464, n70465, n70466, n70467, n70468, n70469, n70470,
    n70471, n70472, n70473, n70474, n70475, n70476, n70477, n70478, n70479,
    n70480, n70481, n70482, n70483, n70484, n70485, n70486, n70487, n70489,
    n70490, n70491, n70492, n70493, n70494, n70495, n70496, n70497, n70498,
    n70499, n70500, n70501, n70502, n70503, n70504, n70505, n70506, n70507,
    n70508, n70509, n70510, n70511, n70512, n70513, n70514, n70515, n70516,
    n70517, n70518, n70519, n70520, n70521, n70522, n70523, n70524, n70525,
    n70526, n70527, n70528, n70529, n70530, n70531, n70532, n70533, n70534,
    n70535, n70536, n70537, n70538, n70539, n70540, n70541, n70542, n70543,
    n70544, n70545, n70546, n70547, n70548, n70549, n70550, n70551, n70552,
    n70553, n70554, n70555, n70556, n70557, n70558, n70559, n70560, n70561,
    n70562, n70563, n70564, n70565, n70566, n70567, n70568, n70569, n70570,
    n70571, n70572, n70573, n70574, n70575, n70576, n70577, n70578, n70579,
    n70580, n70581, n70582, n70583, n70584, n70585, n70586, n70587, n70588,
    n70589, n70590, n70591, n70592, n70593, n70594, n70595, n70596, n70597,
    n70598, n70599, n70600, n70601, n70602, n70603, n70604, n70605, n70606,
    n70607, n70608, n70609, n70610, n70611, n70612, n70613, n70614, n70615,
    n70616, n70617, n70618, n70619, n70620, n70621, n70622, n70623, n70625,
    n70626, n70627, n70628, n70629, n70630, n70631, n70632, n70633, n70634,
    n70635, n70636, n70637, n70638, n70639, n70640, n70641, n70642, n70643,
    n70644, n70645, n70646, n70647, n70648, n70649, n70650, n70651, n70652,
    n70653, n70654, n70655, n70656, n70657, n70658, n70659, n70660, n70661,
    n70662, n70663, n70664, n70665, n70666, n70667, n70668, n70669, n70670,
    n70671, n70672, n70673, n70674, n70675, n70676, n70677, n70678, n70679,
    n70680, n70681, n70682, n70683, n70684, n70685, n70686, n70687, n70688,
    n70689, n70690, n70691, n70692, n70693, n70694, n70695, n70696, n70697,
    n70698, n70699, n70700, n70701, n70702, n70703, n70704, n70705, n70706,
    n70707, n70708, n70709, n70710, n70711, n70712, n70713, n70714, n70715,
    n70716, n70717, n70718, n70719, n70720, n70721, n70722, n70723, n70724,
    n70725, n70726, n70727, n70728, n70729, n70730, n70731, n70732, n70733,
    n70734, n70735, n70736, n70737, n70738, n70739, n70740, n70741, n70742,
    n70743, n70744, n70745, n70746, n70747, n70748, n70749, n70750, n70751,
    n70752, n70753, n70754, n70755, n70756, n70758, n70759, n70760, n70761,
    n70762, n70763, n70764, n70765, n70766, n70767, n70768, n70769, n70770,
    n70771, n70772, n70773, n70774, n70775, n70776, n70777, n70778, n70779,
    n70780, n70781, n70782, n70783, n70784, n70785, n70786, n70787, n70788,
    n70789, n70790, n70791, n70792, n70793, n70794, n70795, n70796, n70797,
    n70798, n70799, n70800, n70801, n70802, n70803, n70804, n70805, n70806,
    n70807, n70808, n70809, n70810, n70811, n70812, n70813, n70814, n70815,
    n70816, n70817, n70818, n70819, n70820, n70821, n70822, n70823, n70824,
    n70825, n70826, n70827, n70828, n70829, n70830, n70831, n70832, n70833,
    n70834, n70835, n70836, n70837, n70838, n70839, n70840, n70841, n70842,
    n70843, n70844, n70845, n70846, n70847, n70848, n70849, n70850, n70851,
    n70852, n70853, n70854, n70855, n70856, n70857, n70858, n70859, n70860,
    n70861, n70862, n70863, n70864, n70865, n70866, n70867, n70868, n70869,
    n70870, n70871, n70872, n70873, n70874, n70875, n70876, n70877, n70878,
    n70879, n70880, n70881, n70882, n70883, n70884, n70885, n70886, n70887,
    n70889, n70890, n70891, n70892, n70893, n70894, n70895, n70896, n70897,
    n70898, n70899, n70900, n70901, n70902, n70903, n70904, n70905, n70906,
    n70907, n70908, n70909, n70910, n70911, n70912, n70913, n70914, n70915,
    n70916, n70917, n70918, n70919, n70920, n70921, n70922, n70923, n70924,
    n70925, n70926, n70927, n70928, n70929, n70930, n70931, n70932, n70933,
    n70934, n70935, n70936, n70937, n70938, n70939, n70940, n70941, n70942,
    n70943, n70944, n70945, n70946, n70947, n70948, n70949, n70950, n70951,
    n70952, n70953, n70954, n70955, n70956, n70957, n70958, n70959, n70960,
    n70961, n70962, n70963, n70964, n70965, n70966, n70967, n70968, n70969,
    n70970, n70971, n70972, n70973, n70974, n70975, n70976, n70977, n70978,
    n70979, n70980, n70981, n70982, n70983, n70984, n70985, n70987, n70988,
    n70989, n70990, n70991, n70992, n70993, n70994, n70995, n70996, n70997,
    n70998, n70999, n71000, n71001, n71002, n71003, n71004, n71005, n71006,
    n71007, n71008, n71009, n71010, n71011, n71012, n71013, n71014, n71015,
    n71016, n71017, n71018, n71019, n71020, n71021, n71022, n71023, n71024,
    n71025, n71026, n71027, n71028, n71029, n71030, n71031, n71032, n71033,
    n71034, n71035, n71036, n71037, n71038, n71039, n71040, n71041, n71042,
    n71043, n71044, n71045, n71046, n71047, n71048, n71049, n71050, n71051,
    n71052, n71053, n71054, n71055, n71056, n71057, n71058, n71059, n71060,
    n71061, n71062, n71063, n71064, n71065, n71066, n71067, n71068, n71069,
    n71070, n71071, n71072, n71073, n71074, n71075, n71077, n71078, n71079,
    n71080, n71081, n71082, n71083, n71084, n71085, n71086, n71087, n71088,
    n71089, n71090, n71091, n71092, n71093, n71094, n71095, n71096, n71097,
    n71098, n71099, n71100, n71101, n71102, n71103, n71104, n71105, n71106,
    n71107, n71108, n71109, n71110, n71111, n71112, n71113, n71114, n71115,
    n71116, n71117, n71118, n71119, n71120, n71121, n71122, n71123, n71124,
    n71125, n71126, n71127, n71128, n71129, n71130, n71131, n71132, n71133,
    n71134, n71135, n71136, n71137, n71138, n71139, n71140, n71141, n71142,
    n71143, n71144, n71145, n71146, n71147, n71148, n71149, n71150, n71151,
    n71152, n71153, n71154, n71155, n71156, n71157, n71158, n71160, n71161,
    n71162, n71163, n71164, n71165, n71166, n71167, n71168, n71169, n71170,
    n71171, n71172, n71173, n71174, n71175, n71176, n71177, n71178, n71179,
    n71180, n71181, n71182, n71183, n71184, n71185, n71186, n71187, n71188,
    n71189, n71190, n71191, n71192, n71193, n71194, n71195, n71196, n71197,
    n71198, n71199, n71200, n71201, n71202, n71203, n71204, n71205, n71206,
    n71207, n71208, n71209, n71210, n71211, n71212, n71213, n71214, n71215,
    n71216, n71217, n71218, n71219, n71220, n71221, n71222, n71223, n71224,
    n71225, n71226, n71227, n71228, n71229, n71230, n71231, n71232, n71233,
    n71234, n71236, n71237, n71238, n71239, n71240, n71241, n71242, n71243,
    n71244, n71245, n71246, n71247, n71248, n71249, n71250, n71251, n71252,
    n71253, n71254, n71255, n71256, n71257, n71258, n71259, n71260, n71261,
    n71262, n71263, n71264, n71265, n71266, n71267, n71268, n71269, n71270,
    n71271, n71272, n71273, n71274, n71275, n71276, n71277, n71278, n71279,
    n71280, n71281, n71282, n71283, n71284, n71285, n71286, n71287, n71288,
    n71289, n71290, n71291, n71292, n71293, n71294, n71295, n71296, n71297,
    n71298, n71299, n71300, n71301, n71302, n71303, n71304, n71305, n71306,
    n71308, n71309, n71310, n71311, n71312, n71313, n71314, n71315, n71316,
    n71317, n71318, n71319, n71320, n71321, n71322, n71323, n71324, n71325,
    n71326, n71327, n71328, n71329, n71330, n71331, n71332, n71333, n71334,
    n71335, n71336, n71337, n71338, n71339, n71340, n71341, n71342, n71343,
    n71344, n71345, n71346, n71347, n71348, n71349, n71350, n71351, n71352,
    n71353, n71354, n71355, n71356, n71357, n71358, n71359, n71360, n71361,
    n71362, n71363, n71364, n71365, n71366, n71367, n71368, n71369, n71370,
    n71371, n71372, n71373, n71374, n71375, n71376, n71377, n71378, n71379,
    n71380, n71381, n71382, n71383, n71384, n71386, n71387, n71388, n71389,
    n71390, n71391, n71392, n71393, n71394, n71395, n71396, n71397, n71398,
    n71399, n71400, n71401, n71402, n71403, n71404, n71405, n71406, n71407,
    n71408, n71409, n71410, n71411, n71412, n71413, n71414, n71415, n71416,
    n71417, n71418, n71419, n71420, n71421, n71422, n71423, n71424, n71425,
    n71426, n71427, n71428, n71429, n71430, n71431, n71432, n71433, n71434,
    n71435, n71436, n71437, n71438, n71439, n71440, n71441, n71442, n71443,
    n71444, n71445, n71446, n71447, n71448, n71449, n71450, n71451, n71452,
    n71453, n71454, n71455, n71456, n71457, n71458, n71459, n71461, n71462,
    n71463, n71464, n71465, n71466, n71467, n71468, n71469, n71470, n71471,
    n71472, n71473, n71474, n71475, n71476, n71477, n71478, n71479, n71480,
    n71481, n71482, n71483, n71484, n71485, n71486, n71487, n71488, n71489,
    n71490, n71491, n71492, n71493, n71494, n71495, n71496, n71497, n71498,
    n71499, n71500, n71501, n71502, n71503, n71504, n71505, n71506, n71507,
    n71508, n71509, n71510, n71511, n71512, n71513, n71514, n71515, n71516,
    n71517, n71518, n71519, n71520, n71521, n71522, n71523, n71524, n71525,
    n71526, n71527, n71528, n71529, n71530, n71531, n71532, n71534, n71535,
    n71536, n71537, n71538, n71539, n71540, n71541, n71542, n71543, n71544,
    n71545, n71546, n71547, n71548, n71549, n71550, n71551, n71552, n71553,
    n71554, n71555, n71556, n71557, n71558, n71559, n71560, n71561, n71562,
    n71563, n71564, n71565, n71566, n71567, n71568, n71569, n71570, n71571,
    n71572, n71573, n71574, n71575, n71576, n71577, n71578, n71579, n71580,
    n71581, n71582, n71583, n71584, n71585, n71586, n71587, n71588, n71589,
    n71590, n71591, n71592, n71593, n71594, n71595, n71596, n71597, n71598,
    n71599, n71600, n71601, n71602, n71603, n71604, n71605, n71606, n71607,
    n71608, n71609, n71610, n71612, n71613, n71614, n71615, n71616, n71617,
    n71618, n71619, n71620, n71621, n71622, n71623, n71624, n71625, n71626,
    n71627, n71628, n71629, n71630, n71631, n71632, n71633, n71634, n71635,
    n71636, n71637, n71638, n71639, n71640, n71641, n71642, n71643, n71644,
    n71645, n71646, n71647, n71648, n71649, n71650, n71651, n71652, n71653,
    n71654, n71655, n71656, n71657, n71658, n71659, n71660, n71661, n71662,
    n71663, n71664, n71665, n71666, n71667, n71668, n71669, n71670, n71671,
    n71672, n71673, n71674, n71675, n71676, n71677, n71678, n71679, n71680,
    n71681, n71682, n71684, n71685, n71686, n71687, n71688, n71689, n71690,
    n71691, n71692, n71693, n71694, n71695, n71696, n71697, n71698, n71699,
    n71700, n71701, n71702, n71703, n71704, n71705, n71706, n71707, n71708,
    n71709, n71710, n71711, n71712, n71713, n71714, n71715, n71716, n71717,
    n71718, n71719, n71720, n71721, n71722, n71723, n71724, n71725, n71726,
    n71727, n71728, n71729, n71730, n71731, n71732, n71733, n71734, n71735,
    n71736, n71737, n71738, n71739, n71740, n71741, n71742, n71743, n71744,
    n71745, n71746, n71747, n71748, n71749, n71750, n71751, n71752, n71753,
    n71754, n71755, n71756, n71757, n71758, n71759, n71760, n71761, n71763,
    n71764, n71765, n71766, n71767, n71768, n71769, n71770, n71771, n71772,
    n71773, n71774, n71775, n71776, n71777, n71778, n71779, n71780, n71781,
    n71782, n71783, n71784, n71785, n71786, n71787, n71788, n71789, n71790,
    n71791, n71792, n71793, n71794, n71795, n71796, n71797, n71798, n71799,
    n71800, n71801, n71802, n71803, n71804, n71805, n71806, n71807, n71808,
    n71809, n71810, n71811, n71812, n71813, n71814, n71815, n71816, n71817,
    n71818, n71819, n71820, n71821, n71822, n71823, n71824, n71825, n71826,
    n71827, n71828, n71829, n71830, n71831, n71832, n71834, n71835, n71836,
    n71837, n71838, n71839, n71840, n71841, n71842, n71843, n71844, n71845,
    n71846, n71847, n71848, n71849, n71850, n71851, n71852, n71853, n71854,
    n71855, n71856, n71857, n71858, n71859, n71860, n71861, n71862, n71863,
    n71864, n71865, n71866, n71867, n71868, n71869, n71870, n71871, n71872,
    n71873, n71874, n71875, n71876, n71877, n71878, n71879, n71880, n71881,
    n71882, n71883, n71884, n71885, n71886, n71887, n71888, n71889, n71890,
    n71891, n71892, n71893, n71894, n71895, n71896, n71897, n71898, n71899,
    n71900, n71901, n71902, n71903, n71904, n71905, n71906, n71907, n71908,
    n71909, n71910, n71912, n71913, n71914, n71915, n71916, n71917, n71918,
    n71919, n71920, n71921, n71922, n71923, n71924, n71925, n71926, n71927,
    n71928, n71929, n71930, n71931, n71932, n71933, n71934, n71935, n71936,
    n71937, n71938, n71939, n71940, n71941, n71942, n71943, n71944, n71945,
    n71946, n71947, n71948, n71949, n71950, n71951, n71952, n71953, n71954,
    n71955, n71956, n71957, n71958, n71959, n71960, n71961, n71962, n71963,
    n71964, n71965, n71966, n71967, n71968, n71969, n71970, n71971, n71972,
    n71973, n71974, n71975, n71976, n71977, n71978, n71979, n71980, n71981,
    n71982, n71983, n71984, n71985, n71986, n71988, n71989, n71990, n71991,
    n71992, n71993, n71994, n71995, n71996, n71997, n71998, n71999, n72000,
    n72001, n72002, n72003, n72004, n72005, n72006, n72007, n72008, n72009,
    n72010, n72011, n72012, n72013, n72014, n72015, n72016, n72017, n72018,
    n72019, n72020, n72021, n72022, n72023, n72024, n72025, n72026, n72027,
    n72028, n72029, n72030, n72031, n72032, n72033, n72034, n72035, n72036,
    n72037, n72038, n72039, n72040, n72041, n72042, n72043, n72044, n72045,
    n72046, n72047, n72048, n72049, n72050, n72051, n72052, n72053, n72054,
    n72055, n72056, n72057, n72058, n72059, n72061, n72062, n72063, n72064,
    n72065, n72066, n72067, n72068, n72069, n72070, n72071, n72072, n72073,
    n72074, n72075, n72076, n72077, n72078, n72079, n72080, n72081, n72082,
    n72083, n72084, n72085, n72086, n72087, n72088, n72089, n72090, n72091,
    n72092, n72093, n72094, n72095, n72096, n72097, n72098, n72099, n72100,
    n72101, n72102, n72103, n72104, n72105, n72106, n72107, n72108, n72109,
    n72110, n72111, n72112, n72113, n72114, n72115, n72116, n72117, n72118,
    n72119, n72120, n72121, n72122, n72123, n72124, n72125, n72126, n72127,
    n72128, n72129, n72130, n72131, n72132, n72133, n72134, n72135, n72136,
    n72138, n72139, n72140, n72141, n72142, n72143, n72144, n72145, n72146,
    n72147, n72148, n72149, n72150, n72151, n72152, n72153, n72154, n72155,
    n72156, n72157, n72158, n72159, n72160, n72161, n72162, n72163, n72164,
    n72165, n72166, n72167, n72168, n72169, n72170, n72171, n72172, n72173,
    n72174, n72175, n72176, n72177, n72178, n72179, n72180, n72181, n72182,
    n72183, n72184, n72185, n72186, n72187, n72188, n72189, n72190, n72191,
    n72192, n72193, n72194, n72195, n72196, n72197, n72198, n72199, n72200,
    n72201, n72202, n72203, n72204, n72205, n72206, n72207, n72208, n72209,
    n72210, n72211, n72212, n72213, n72215, n72216, n72217, n72218, n72219,
    n72220, n72221, n72222, n72223, n72224, n72225, n72226, n72227, n72228,
    n72229, n72230, n72231, n72232, n72233, n72234, n72235, n72236, n72237,
    n72238, n72239, n72240, n72241, n72242, n72243, n72244, n72245, n72246,
    n72247, n72248, n72249, n72250, n72251, n72252, n72253, n72254, n72255,
    n72256, n72257, n72258, n72259, n72260, n72261, n72262, n72263, n72264,
    n72265, n72266, n72267, n72268, n72269, n72270, n72271, n72272, n72273,
    n72274, n72275, n72276, n72277, n72278, n72279, n72280, n72281, n72282,
    n72283, n72284, n72285, n72286, n72287, n72289, n72290, n72291, n72292,
    n72293, n72294, n72295, n72296, n72297, n72298, n72299, n72300, n72301,
    n72302, n72303, n72304, n72305, n72306, n72307, n72308, n72309, n72310,
    n72311, n72312, n72313, n72314, n72315, n72316, n72317, n72318, n72319,
    n72320, n72321, n72322, n72323, n72324, n72325, n72326, n72327, n72328,
    n72329, n72330, n72331, n72332, n72333, n72334, n72335, n72336, n72337,
    n72338, n72339, n72340, n72341, n72342, n72343, n72344, n72345, n72346,
    n72347, n72348, n72349, n72350, n72351, n72352, n72353, n72354, n72355,
    n72356, n72357, n72358, n72359, n72360, n72361, n72362, n72363, n72364,
    n72365, n72367, n72368, n72369, n72370, n72371, n72372, n72373, n72374,
    n72375, n72376, n72377, n72378, n72379, n72380, n72381, n72382, n72383,
    n72384, n72385, n72386, n72387, n72388, n72389, n72390, n72391, n72392,
    n72393, n72394, n72395, n72396, n72397, n72398, n72399, n72400, n72401,
    n72402, n72403, n72404, n72405, n72406, n72407, n72408, n72409, n72410,
    n72411, n72412, n72413, n72414, n72415, n72416, n72417, n72418, n72419,
    n72420, n72421, n72422, n72423, n72424, n72425, n72426, n72427, n72428,
    n72429, n72430, n72431, n72432, n72433, n72434, n72435, n72436, n72437,
    n72438, n72439, n72440, n72442, n72443, n72444, n72445, n72446, n72447,
    n72448, n72449, n72450, n72451, n72452, n72453, n72454, n72455, n72456,
    n72457, n72458, n72459, n72460, n72461, n72462, n72463, n72464, n72465,
    n72466, n72467, n72468, n72469, n72470, n72471, n72472, n72473, n72474,
    n72475, n72476, n72477, n72478, n72479, n72480, n72481, n72482, n72483,
    n72484, n72485, n72486, n72487, n72488, n72489, n72490, n72491, n72492,
    n72493, n72494, n72495, n72496, n72497, n72498, n72499, n72500, n72501,
    n72502, n72503, n72504, n72505, n72506, n72507, n72508, n72509, n72510,
    n72511, n72513, n72514, n72515, n72516, n72517, n72518, n72519, n72520,
    n72521, n72522, n72523, n72524, n72525, n72526, n72527, n72528, n72529,
    n72530, n72531, n72532, n72533, n72534, n72535, n72536, n72537, n72538,
    n72539, n72540, n72541, n72542, n72543, n72544, n72545, n72546, n72547,
    n72548, n72549, n72550, n72551, n72552, n72553, n72554, n72555, n72556,
    n72557, n72558, n72559, n72560, n72561, n72562, n72563, n72564, n72565,
    n72566, n72567, n72568, n72569, n72570, n72571, n72572, n72573, n72574,
    n72575, n72576, n72577, n72578, n72579, n72580, n72581, n72582, n72583,
    n72584, n72585, n72586, n72587, n72588, n72589, n72590, n72591, n72593,
    n72594, n72595, n72596, n72597, n72598, n72599, n72600, n72601, n72602,
    n72603, n72604, n72605, n72606, n72607, n72608, n72609, n72610, n72611,
    n72612, n72613, n72614, n72615, n72616, n72617, n72618, n72619, n72620,
    n72621, n72622, n72623, n72624, n72625, n72626, n72627, n72628, n72629,
    n72630, n72631, n72632, n72633, n72634, n72635, n72636, n72637, n72638,
    n72639, n72640, n72641, n72642, n72643, n72644, n72645, n72646, n72647,
    n72648, n72649, n72650, n72651, n72652, n72653, n72654, n72655, n72656,
    n72657, n72658, n72659, n72660, n72661, n72662, n72664, n72665, n72666,
    n72667, n72668, n72669, n72670, n72671, n72672, n72673, n72674, n72675,
    n72676, n72677, n72678, n72679, n72680, n72681, n72682, n72683, n72684,
    n72685, n72686, n72687, n72688, n72689, n72690, n72691, n72692, n72693,
    n72694, n72695, n72696, n72697, n72698, n72699, n72700, n72701, n72702,
    n72703, n72704, n72705, n72706, n72707, n72708, n72709, n72710, n72711,
    n72712, n72713, n72714, n72715, n72716, n72717, n72718, n72719, n72720,
    n72721, n72722, n72723, n72724, n72725, n72726, n72727, n72728, n72729,
    n72730, n72731, n72732, n72733, n72734, n72736, n72737, n72738, n72739,
    n72740, n72741, n72742, n72743, n72744, n72745, n72746, n72747, n72748,
    n72749, n72750, n72751, n72752, n72753, n72754, n72755, n72756, n72757,
    n72758, n72759, n72760, n72761, n72762, n72763, n72764, n72765, n72766,
    n72767, n72768, n72769, n72770, n72771, n72772, n72773, n72774, n72775,
    n72776, n72777, n72778, n72779, n72780, n72781, n72782, n72783, n72784,
    n72785, n72786, n72787, n72788, n72789, n72790, n72791, n72792, n72793,
    n72794, n72795, n72796, n72797, n72798, n72799, n72800, n72801, n72802,
    n72803, n72804, n72805, n72806, n72807, n72808, n72809, n72810, n72811,
    n72812, n72813, n72814, n72815, n72816, n72818, n72819, n72820, n72821,
    n72822, n72823, n72824, n72825, n72826, n72827, n72828, n72829, n72830,
    n72831, n72832, n72833, n72834, n72835, n72836, n72837, n72838, n72839,
    n72840, n72841, n72842, n72843, n72844, n72845, n72846, n72847, n72848,
    n72849, n72851, n72852, n72853, n72854, n72855, n72856, n72857, n72858,
    n72859, n72860, n72861, n72862, n72863, n72864, n72866, n72867, n72868,
    n72869, n72870, n72871, n72872, n72873, n72874, n72875, n72876, n72877,
    n72878, n72879, n72880, n72881, n72882, n72884, n72885, n72886, n72887,
    n72888, n72889, n72890, n72891, n72892, n72893, n72894, n72895, n72896,
    n72897, n72898, n72899, n72900, n72901, n72902, n72903, n72904, n72906,
    n72907, n72908, n72909, n72910, n72911, n72912, n72913, n72914, n72915,
    n72916, n72917, n72918, n72919, n72920, n72921, n72922, n72923, n72924,
    n72925, n72926, n72927, n72929, n72930, n72931, n72932, n72933, n72934,
    n72935, n72936, n72937, n72938, n72939, n72940, n72941, n72942, n72943,
    n72944, n72945, n72946, n72947, n72948, n72949, n72950, n72952, n72953,
    n72954, n72955, n72956, n72957, n72958, n72959, n72960, n72961, n72962,
    n72963, n72964, n72965, n72966, n72967, n72968, n72969, n72970, n72971,
    n72972, n72973, n72975, n72976, n72977, n72978, n72979, n72980, n72981,
    n72982, n72983, n72984, n72985, n72986, n72987, n72988, n72989, n72990,
    n72991, n72992, n72993, n72994, n72995, n72996, n72998, n72999, n73000,
    n73001, n73002, n73003, n73004, n73005, n73006, n73007, n73008, n73009,
    n73010, n73011, n73012, n73013, n73014, n73015, n73016, n73017, n73018,
    n73019, n73021, n73022, n73023, n73024, n73025, n73026, n73027, n73028,
    n73029, n73030, n73031, n73032, n73033, n73034, n73035, n73036, n73037,
    n73038, n73039, n73040, n73041, n73042, n73044, n73045, n73046, n73047,
    n73048, n73049, n73050, n73051, n73052, n73053, n73054, n73055, n73056,
    n73057, n73058, n73059, n73060, n73061, n73062, n73063, n73064, n73065,
    n73067, n73068, n73069, n73070, n73071, n73072, n73073, n73074, n73075,
    n73076, n73077, n73078, n73079, n73080, n73081, n73082, n73083, n73084,
    n73085, n73086, n73087, n73088, n73090, n73091, n73092, n73093, n73094,
    n73095, n73096, n73097, n73098, n73099, n73100, n73101, n73102, n73103,
    n73104, n73105, n73106, n73107, n73108, n73109, n73110, n73111, n73113,
    n73114, n73115, n73116, n73117, n73118, n73119, n73120, n73121, n73122,
    n73123, n73124, n73125, n73126, n73127, n73128, n73129, n73130, n73131,
    n73132, n73133, n73134, n73136, n73137, n73138, n73139, n73140, n73141,
    n73142, n73143, n73144, n73145, n73146, n73147, n73148, n73149, n73150,
    n73151, n73152, n73153, n73154, n73155, n73156, n73157, n73159, n73160,
    n73161, n73162, n73163, n73164, n73165, n73166, n73167, n73168, n73169,
    n73170, n73171, n73172, n73173, n73174, n73175, n73176, n73177, n73178,
    n73179, n73180, n73182, n73183, n73184, n73185, n73186, n73187, n73188,
    n73189, n73190, n73191, n73192, n73193, n73194, n73195, n73196, n73197,
    n73198, n73199, n73200, n73201, n73202, n73203, n73205, n73206, n73207,
    n73208, n73209, n73210, n73211, n73212, n73213, n73214, n73215, n73216,
    n73217, n73218, n73219, n73220, n73221, n73222, n73223, n73224, n73225,
    n73226, n73228, n73229, n73230, n73231, n73232, n73233, n73234, n73235,
    n73236, n73237, n73238, n73239, n73240, n73241, n73242, n73243, n73244,
    n73245, n73246, n73247, n73248, n73249, n73251, n73252, n73253, n73254,
    n73255, n73256, n73257, n73258, n73259, n73260, n73261, n73262, n73263,
    n73264, n73265, n73266, n73267, n73268, n73269, n73270, n73271, n73272,
    n73274, n73275, n73276, n73277, n73278, n73279, n73280, n73281, n73282,
    n73283, n73284, n73285, n73286, n73287, n73288, n73289, n73290, n73291,
    n73292, n73293, n73294, n73295, n73297, n73298, n73299, n73300, n73301,
    n73302, n73303, n73304, n73305, n73306, n73307, n73308, n73309, n73310,
    n73311, n73312, n73313, n73314, n73315, n73316, n73317, n73318, n73320,
    n73321, n73322, n73323, n73324, n73325, n73326, n73327, n73328, n73329,
    n73330, n73331, n73332, n73333, n73334, n73335, n73336, n73337, n73338,
    n73339, n73340, n73341, n73343, n73344, n73345, n73346, n73347, n73348,
    n73349, n73350, n73351, n73352, n73353, n73354, n73355, n73356, n73357,
    n73358, n73359, n73360, n73361, n73362, n73363, n73364, n73366, n73367,
    n73368, n73369, n73370, n73371, n73372, n73373, n73374, n73375, n73376,
    n73377, n73378, n73379, n73380, n73381, n73382, n73383, n73384, n73385,
    n73386, n73387, n73389, n73390, n73391, n73392, n73393, n73394, n73395,
    n73396, n73397, n73398, n73399, n73400, n73401, n73402, n73403, n73404,
    n73405, n73406, n73407, n73408, n73409, n73410, n73412, n73413, n73414,
    n73415, n73416, n73417, n73418, n73419, n73420, n73421, n73422, n73423,
    n73424, n73425, n73426, n73427, n73428, n73429, n73430, n73431, n73432,
    n73433, n73435, n73436, n73437, n73438, n73439, n73440, n73441, n73442,
    n73443, n73444, n73445, n73446, n73447, n73448, n73449, n73450, n73451,
    n73452, n73453, n73454, n73455, n73456, n73458, n73459, n73460, n73461,
    n73462, n73463, n73464, n73465, n73466, n73467, n73468, n73469, n73470,
    n73471, n73472, n73473, n73474, n73475, n73476, n73477, n73478, n73479,
    n73481, n73482, n73483, n73484, n73485, n73486, n73487, n73488, n73489,
    n73490, n73491, n73492, n73493, n73494, n73495, n73496, n73497, n73498,
    n73499, n73500, n73501, n73502, n73504, n73505, n73506, n73507, n73508,
    n73509, n73510, n73511, n73512, n73513, n73514, n73515, n73516, n73517,
    n73518, n73519, n73520, n73521, n73522, n73523, n73524, n73525, n73527,
    n73528, n73529, n73530, n73531, n73532, n73533, n73534, n73535, n73536,
    n73537, n73538, n73539, n73540, n73541, n73542, n73543, n73544, n73545,
    n73546, n73547, n73548, n73550, n73551, n73552, n73553, n73554, n73555,
    n73556, n73557, n73558, n73559, n73560, n73561, n73562, n73564, n73565,
    n73566, n73567, n73568, n73569, n73570, n73572, n73573, n73574, n73575,
    n73576, n73577, n73578, n73580, n73581, n73582, n73583, n73584, n73585,
    n73586, n73588, n73589, n73590, n73591, n73592, n73593, n73594, n73596,
    n73597, n73598, n73599, n73600, n73601, n73602, n73604, n73605, n73606,
    n73607, n73608, n73609, n73610, n73612, n73613, n73614, n73615, n73616,
    n73617, n73618, n73620, n73621, n73622, n73623, n73625, n73626, n73627,
    n73628, n73630, n73631, n73632, n73633, n73635, n73636, n73637, n73638,
    n73640, n73641, n73642, n73643, n73645, n73646, n73647, n73648, n73650,
    n73651, n73652, n73653, n73655, n73656, n73657, n73658, n73660, n73661,
    n73662, n73664, n73665, n73666, n73668, n73669, n73670, n73672, n73673,
    n73674, n73676, n73677, n73678, n73680, n73681, n73682, n73684, n73685,
    n73686, n73688, n73689, n73690, n73692, n73693, n73694, n73696, n73697,
    n73698, n73700, n73701, n73702, n73704, n73705, n73706, n73708, n73709,
    n73710, n73712, n73713, n73714, n73716, n73717, n73718, n73720, n73721,
    n73722, n73723, n73724, n73725, n73726, n73727, n73728, n73729, n73731,
    n73732, n73733, n73734, n73736, n73737, n73738, n73739, n73741, n73742,
    n73743, n73744, n73746, n73747, n73748, n73749, n73751, n73752, n73753,
    n73754, n73756, n73757, n73758, n73759, n73761, n73762, n73763, n73764,
    n73766, n73767, n73768, n73769, n73771, n73772, n73773, n73774, n73776,
    n73777, n73778, n73779, n73781, n73782, n73783, n73784, n73786, n73787,
    n73788, n73789, n73791, n73792, n73793, n73794, n73796, n73797, n73798,
    n73799, n73801, n73802, n73803, n73804, n73806, n73807, n73808, n73809,
    n73810, n73812, n73813, n73814, n73815, n73817, n73818, n73819, n73820,
    n73822, n73823, n73824, n73825, n73827, n73828, n73829, n73830, n73832,
    n73833, n73834, n73835, n73837, n73838, n73839, n73840, n73842, n73843,
    n73844, n73845, n73847, n73848, n73849, n73850, n73852, n73853, n73854,
    n73855, n73857, n73858, n73859, n73860, n73862, n73863, n73864, n73865,
    n73867, n73868, n73869, n73870, n73872, n73873, n73874, n73875, n73877,
    n73878, n73879, n73880, n73883, n73884, n73885, n73886, n73887, n73888,
    n73889, n73890, n73891, n73892, n73893, n73894, n73896, n73897, n73898,
    n73899, n73900, n73901, n73902, n73903, n73904, n73906, n73907, n73908,
    n73909, n73910, n73911, n73912, n73913, n73914, n73915, n73917, n73918,
    n73919, n73920, n73921, n73922, n73923, n73924, n73925, n73926, n73927,
    n73929, n73930, n73931, n73932, n73933, n73934, n73935, n73936, n73937,
    n73938, n73940, n73941, n73942, n73943, n73944, n73945, n73946, n73947,
    n73948, n73949, n73950, n73952, n73953, n73954, n73955, n73956, n73957,
    n73958, n73959, n73960, n73961, n73963, n73964, n73965, n73966, n73967,
    n73968, n73969, n73970, n73971, n73972, n73973, n73975, n73976, n73977,
    n73978, n73979, n73980, n73981, n73982, n73983, n73984, n73985, n73986,
    n73987, n73988, n73989, n73990, n73991, n73992, n73993, n73994, n73995,
    n73996, n73997, n73998, n73999, n74000, n74001, n74002, n74003, n74004,
    n74005, n74006, n74007, n74008, n74009, n74010, n74011, n74012, n74013,
    n74014, n74015, n74016, n74017, n74018, n74019, n74020, n74021, n74022,
    n74023, n74024, n74025, n74026, n74027, n74028, n74029, n74030, n74031,
    n74032, n74033, n74034, n74035, n74036, n74038, n74039, n74040, n74041,
    n74042, n74043, n74044, n74045, n74046, n74047, n74048, n74049, n74050,
    n74051, n74052, n74053, n74054, n74055, n74056, n74057, n74058, n74059,
    n74060, n74061, n74062, n74063, n74064, n74065, n74066, n74067, n74068,
    n74069, n74070, n74071, n74072, n74073, n74074, n74075, n74076, n74077,
    n74078, n74079, n74081, n74082, n74083, n74084, n74085, n74086, n74087,
    n74088, n74089, n74090, n74091, n74092, n74093, n74094, n74095, n74096,
    n74097, n74098, n74099, n74100, n74101, n74102, n74103, n74104, n74105,
    n74106, n74107, n74108, n74109, n74110, n74111, n74112, n74113, n74114,
    n74115, n74116, n74117, n74118, n74119, n74120, n74121, n74123, n74124,
    n74125, n74126, n74127, n74128, n74129, n74130, n74131, n74132, n74133,
    n74134, n74135, n74136, n74137, n74138, n74139, n74140, n74141, n74142,
    n74143, n74144, n74145, n74146, n74147, n74148, n74149, n74150, n74151,
    n74152, n74153, n74154, n74155, n74156, n74157, n74158, n74159, n74160,
    n74161, n74162, n74163, n74164, n74166, n74167, n74168, n74169, n74170,
    n74171, n74172, n74173, n74174, n74175, n74176, n74177, n74178, n74179,
    n74180, n74181, n74182, n74183, n74184, n74185, n74186, n74187, n74188,
    n74189, n74190, n74191, n74192, n74193, n74194, n74195, n74196, n74197,
    n74198, n74199, n74200, n74201, n74202, n74203, n74204, n74205, n74206,
    n74208, n74209, n74210, n74211, n74212, n74213, n74214, n74215, n74216,
    n74217, n74218, n74219, n74220, n74221, n74222, n74223, n74224, n74225,
    n74226, n74227, n74228, n74229, n74230, n74231, n74232, n74233, n74234,
    n74235, n74236, n74237, n74238, n74239, n74240, n74241, n74242, n74243,
    n74244, n74245, n74246, n74247, n74248, n74249, n74251, n74252, n74253,
    n74254, n74255, n74256, n74257, n74258, n74259, n74260, n74261, n74262,
    n74263, n74264, n74265, n74266, n74267, n74268, n74269, n74270, n74271,
    n74272, n74273, n74274, n74275, n74276, n74277, n74278, n74279, n74280,
    n74281, n74282, n74283, n74284, n74285, n74286, n74287, n74288, n74289,
    n74290, n74291, n74293, n74294, n74295, n74296, n74297, n74298, n74299,
    n74300, n74301, n74302, n74303, n74304, n74305, n74306, n74307, n74308,
    n74309, n74310, n74311, n74312, n74313, n74314, n74315, n74316, n74317,
    n74318, n74319, n74320, n74321, n74322, n74323, n74324, n74325, n74326,
    n74327, n74328, n74329, n74330, n74331, n74332, n74333, n74334, n74336,
    n74337, n74338, n74339, n74340, n74341, n74342, n74343, n74344, n74345,
    n74346, n74347, n74348, n74349, n74350, n74351, n74352, n74353, n74354,
    n74355, n74356, n74357, n74358, n74359, n74360, n74361, n74362, n74363,
    n74364, n74365, n74366, n74367, n74368, n74369, n74370, n74371, n74372,
    n74373, n74374, n74375, n74376, n74377, n74378, n74379, n74380, n74381,
    n74382, n74383, n74384, n74385, n74386, n74387, n74388, n74389, n74390,
    n74391, n74392, n74393, n74394, n74395, n74396, n74397, n74398, n74399,
    n74400, n74401, n74402, n74403, n74404, n74405, n74407, n74408, n74409,
    n74410, n74411, n74412, n74413, n74414, n74415, n74416, n74417, n74418,
    n74419, n74420, n74421, n74422, n74423, n74424, n74425, n74426, n74427,
    n74428, n74429, n74430, n74431, n74432, n74433, n74434, n74435, n74436,
    n74437, n74438, n74439, n74440, n74441, n74442, n74443, n74444, n74445,
    n74446, n74447, n74448, n74449, n74450, n74452, n74453, n74454, n74455,
    n74456, n74457, n74458, n74459, n74460, n74461, n74462, n74463, n74464,
    n74465, n74466, n74467, n74468, n74469, n74470, n74471, n74472, n74473,
    n74474, n74475, n74476, n74477, n74478, n74479, n74480, n74481, n74482,
    n74483, n74484, n74485, n74486, n74487, n74488, n74489, n74490, n74491,
    n74492, n74493, n74494, n74496, n74497, n74498, n74499, n74500, n74501,
    n74502, n74503, n74504, n74505, n74506, n74507, n74508, n74509, n74510,
    n74511, n74512, n74513, n74514, n74515, n74516, n74517, n74518, n74519,
    n74520, n74521, n74522, n74523, n74524, n74525, n74526, n74527, n74528,
    n74529, n74530, n74531, n74532, n74533, n74534, n74535, n74536, n74537,
    n74538, n74539, n74541, n74542, n74543, n74544, n74545, n74546, n74547,
    n74548, n74549, n74550, n74551, n74552, n74553, n74554, n74555, n74556,
    n74557, n74558, n74559, n74560, n74561, n74562, n74563, n74564, n74565,
    n74566, n74567, n74568, n74569, n74570, n74571, n74572, n74573, n74574,
    n74575, n74576, n74577, n74578, n74579, n74580, n74581, n74582, n74583,
    n74585, n74586, n74587, n74588, n74589, n74590, n74591, n74592, n74593,
    n74594, n74595, n74596, n74597, n74598, n74599, n74600, n74601, n74602,
    n74603, n74604, n74605, n74606, n74607, n74608, n74609, n74610, n74611,
    n74612, n74613, n74614, n74615, n74616, n74617, n74618, n74619, n74620,
    n74621, n74622, n74623, n74624, n74625, n74626, n74627, n74628, n74630,
    n74631, n74632, n74633, n74634, n74635, n74636, n74637, n74638, n74639,
    n74640, n74641, n74642, n74643, n74644, n74645, n74646, n74647, n74648,
    n74649, n74650, n74651, n74652, n74653, n74654, n74655, n74656, n74657,
    n74658, n74659, n74660, n74661, n74662, n74663, n74664, n74665, n74666,
    n74667, n74668, n74669, n74670, n74671, n74672, n74674, n74675, n74676,
    n74677, n74678, n74679, n74680, n74681, n74682, n74683, n74684, n74685,
    n74686, n74687, n74688, n74689, n74690, n74691, n74692, n74693, n74694,
    n74695, n74696, n74697, n74698, n74699, n74700, n74701, n74702, n74703,
    n74704, n74705, n74706, n74707, n74708, n74709, n74710, n74711, n74712,
    n74713, n74714, n74715, n74716, n74717, n74718, n74719, n74720, n74721,
    n74722, n74723, n74724, n74725, n74726, n74727, n74728, n74729, n74730,
    n74731, n74732, n74733, n74734, n74735, n74736, n74737, n74738, n74739,
    n74740, n74741, n74742, n74743, n74744, n74745, n74746, n74747, n74748,
    n74749, n74750, n74751, n74752, n74753, n74754, n74755, n74756, n74757,
    n74758, n74759, n74760, n74761, n74762, n74763, n74764, n74765, n74766,
    n74767, n74768, n74769, n74770, n74771, n74773, n74774, n74775, n74776,
    n74777, n74778, n74779, n74780, n74781, n74782, n74783, n74784, n74785,
    n74786, n74787, n74788, n74789, n74790, n74791, n74792, n74793, n74794,
    n74795, n74796, n74797, n74798, n74799, n74800, n74801, n74802, n74803,
    n74804, n74805, n74806, n74807, n74808, n74809, n74810, n74811, n74812,
    n74813, n74814, n74815, n74816, n74817, n74818, n74819, n74821, n74822,
    n74823, n74824, n74825, n74826, n74827, n74828, n74829, n74830, n74831,
    n74832, n74833, n74834, n74835, n74836, n74837, n74838, n74839, n74840,
    n74841, n74842, n74843, n74844, n74845, n74846, n74847, n74848, n74849,
    n74850, n74851, n74852, n74853, n74854, n74855, n74856, n74857, n74858,
    n74859, n74860, n74861, n74862, n74863, n74864, n74865, n74866, n74867,
    n74868, n74870, n74871, n74872, n74873, n74874, n74875, n74876, n74877,
    n74878, n74879, n74880, n74881, n74882, n74883, n74884, n74885, n74886,
    n74887, n74888, n74889, n74890, n74891, n74892, n74893, n74894, n74895,
    n74896, n74897, n74898, n74899, n74900, n74901, n74902, n74903, n74904,
    n74905, n74906, n74907, n74908, n74909, n74910, n74911, n74912, n74913,
    n74914, n74915, n74916, n74918, n74919, n74920, n74921, n74922, n74923,
    n74924, n74925, n74926, n74927, n74928, n74929, n74930, n74931, n74932,
    n74933, n74934, n74935, n74936, n74937, n74938, n74939, n74940, n74941,
    n74942, n74943, n74944, n74945, n74946, n74947, n74948, n74949, n74950,
    n74951, n74952, n74953, n74954, n74955, n74956, n74957, n74958, n74959,
    n74960, n74961, n74962, n74963, n74964, n74965, n74967, n74968, n74969,
    n74970, n74971, n74972, n74973, n74974, n74975, n74976, n74977, n74978,
    n74979, n74980, n74981, n74982, n74983, n74984, n74985, n74986, n74987,
    n74988, n74989, n74990, n74991, n74992, n74993, n74994, n74995, n74996,
    n74997, n74998, n74999, n75000, n75001, n75002, n75003, n75004, n75005,
    n75006, n75007, n75008, n75009, n75010, n75011, n75012, n75013, n75015,
    n75016, n75017, n75018, n75019, n75020, n75021, n75022, n75023, n75024,
    n75025, n75026, n75027, n75028, n75029, n75030, n75031, n75032, n75033,
    n75034, n75035, n75036, n75037, n75038, n75039, n75040, n75041, n75042,
    n75043, n75044, n75045, n75046, n75047, n75048, n75049, n75050, n75051,
    n75052, n75053, n75054, n75055, n75056, n75057, n75058, n75059, n75060,
    n75061, n75062, n75064, n75065, n75066, n75067, n75068, n75069, n75070,
    n75071, n75072, n75073, n75074, n75075, n75076, n75077, n75078, n75079,
    n75080, n75081, n75082, n75083, n75084, n75085, n75086, n75087, n75088,
    n75089, n75090, n75091, n75092, n75093, n75094, n75095, n75096, n75097,
    n75098, n75099, n75100, n75101, n75102, n75103, n75104, n75105, n75106,
    n75107, n75108, n75109, n75110, n75112, n75113, n75114, n75115, n75116,
    n75117, n75118, n75119, n75121, n75122, n75123, n75124, n75125, n75126,
    n75127, n75128, n75130, n75131, n75132, n75133, n75134, n75135, n75136,
    n75138, n75139, n75140, n75141, n75142, n75143, n75144, n75145, n75147,
    n75148, n75149, n75150, n75151, n75152, n75153, n75154, n75155, n75157,
    n75158, n75159, n75160, n75161, n75162, n75163, n75164, n75166, n75167,
    n75168, n75169, n75170, n75171, n75172, n75173, n75174, n75176, n75177,
    n75178, n75179, n75180, n75181, n75182, n75183, n75185, n75186, n75187,
    n75188, n75189, n75190, n75191, n75192, n75193, n75195, n75196, n75197,
    n75198, n75199, n75200, n75201, n75202, n75204, n75205, n75206, n75207,
    n75208, n75209, n75210, n75211, n75212, n75214, n75215, n75216, n75217,
    n75218, n75219, n75220, n75221, n75223, n75224, n75225, n75226, n75227,
    n75228, n75229, n75230, n75231, n75233, n75234, n75235, n75236, n75237,
    n75238, n75239, n75240, n75242, n75243, n75244, n75245, n75246, n75247,
    n75248, n75249, n75250, n75252, n75253, n75254, n75255, n75256, n75257,
    n75258, n75259, n75261, n75262, n75263, n75264, n75265, n75266, n75267,
    n75268, n75269, n75271, n75272, n75273, n75274, n75275, n75276, n75277,
    n75278, n75280, n75281, n75282, n75283, n75284, n75285, n75286, n75287,
    n75288, n75290, n75291, n75292, n75293, n75294, n75295, n75296, n75297,
    n75299, n75300, n75301, n75302, n75303, n75304, n75305, n75306, n75307,
    n75309, n75310, n75311, n75312, n75313, n75314, n75315, n75316, n75318,
    n75319, n75320, n75321, n75322, n75323, n75324, n75325, n75326, n75328,
    n75329, n75330, n75331, n75332, n75333, n75334, n75335, n75337, n75338,
    n75339, n75340, n75341, n75342, n75343, n75344, n75345, n75347, n75348,
    n75349, n75350, n75351, n75352, n75353, n75354, n75356, n75357, n75358,
    n75359, n75360, n75361, n75362, n75363, n75364, n75366, n75367, n75368,
    n75369, n75370, n75371, n75372, n75373, n75375, n75376, n75377, n75378,
    n75379, n75380, n75381, n75382, n75383, n75385, n75386, n75387, n75388,
    n75389, n75390, n75391, n75392, n75394, n75395, n75396, n75397, n75398,
    n75399, n75400, n75401, n75402, n75404, n75405, n75406, n75407, n75408,
    n75409, n75410, n75411, n75413, n75414, n75415, n75416, n75417, n75418,
    n75420, n75421, n75422, n75423, n75424, n75425, n75426, n75427, n75428,
    n75429, n75430, n75431, n75432, n75433, n75434, n75435, n75436, n75437,
    n75438, n75439, n75440, n75441, n75442, n75443, n75444, n75445, n75446,
    n75447, n75448, n75449, n75450, n75451, n75452, n75453, n75454, n75455,
    n75456, n75457, n75458, n75459, n75460, n75461, n75463, n75464, n75465,
    n75466, n75467, n75468, n75469, n75470, n75471, n75472, n75473, n75474,
    n75475, n75476, n75477, n75478, n75479, n75480, n75481, n75482, n75483,
    n75484, n75486, n75487, n75488, n75489, n75490, n75491, n75492, n75493,
    n75494, n75495, n75496, n75497, n75498, n75499, n75500, n75501, n75502,
    n75503, n75504, n75505, n75506, n75507, n75508, n75509, n75510, n75511,
    n75512, n75513, n75514, n75516, n75517, n75518, n75519, n75520, n75521,
    n75522, n75523, n75524, n75525, n75526, n75527, n75528, n75529, n75530,
    n75531, n75532, n75533, n75534, n75535, n75536, n75537, n75538, n75539,
    n75540, n75541, n75542, n75543, n75544, n75545, n75547, n75548, n75549,
    n75550, n75551, n75552, n75553, n75554, n75555, n75556, n75557, n75558,
    n75559, n75560, n75561, n75562, n75563, n75564, n75565, n75566, n75567,
    n75568, n75569, n75570, n75571, n75572, n75573, n75574, n75575, n75576,
    n75577, n75578, n75579, n75580, n75581, n75582, n75584, n75585, n75586,
    n75587, n75588, n75589, n75590, n75591, n75592, n75593, n75594, n75595,
    n75596, n75597, n75598, n75599, n75600, n75601, n75602, n75603, n75604,
    n75605, n75606, n75607, n75608, n75609, n75610, n75611, n75612, n75613,
    n75615, n75616, n75617, n75618, n75619, n75620, n75621, n75622, n75623,
    n75624, n75625, n75626, n75627, n75628, n75629, n75630, n75631, n75632,
    n75633, n75634, n75635, n75636, n75637, n75638, n75639, n75640, n75641,
    n75643, n75644, n75645, n75646, n75647, n75648, n75649, n75650, n75651,
    n75652, n75653, n75654, n75655, n75656, n75657, n75658, n75659, n75660,
    n75661, n75662, n75663, n75664, n75665, n75666, n75667, n75669, n75670,
    n75671, n75672, n75673, n75674, n75675, n75676, n75677, n75678, n75679,
    n75680, n75681, n75682, n75683, n75684, n75685, n75686, n75687, n75688,
    n75689, n75690, n75691, n75692, n75693, n75694, n75695, n75697, n75698,
    n75699, n75700, n75701, n75702, n75703, n75704, n75705, n75706, n75707,
    n75708, n75709, n75710, n75711, n75712, n75713, n75714, n75715, n75716,
    n75717, n75718, n75719, n75720, n75721, n75723, n75724, n75725, n75726,
    n75727, n75728, n75729, n75730, n75731, n75732, n75733, n75734, n75735,
    n75736, n75737, n75738, n75739, n75740, n75741, n75742, n75743, n75744,
    n75745, n75746, n75747, n75748, n75749, n75751, n75752, n75753, n75754,
    n75755, n75756, n75757, n75758, n75759, n75760, n75761, n75762, n75763,
    n75764, n75765, n75766, n75767, n75768, n75769, n75770, n75771, n75772,
    n75773, n75774, n75775, n75777, n75778, n75779, n75780, n75781, n75782,
    n75783, n75784, n75785, n75786, n75787, n75788, n75789, n75790, n75791,
    n75792, n75793, n75794, n75795, n75796, n75797, n75798, n75799, n75800,
    n75801, n75802, n75803, n75805, n75806, n75807, n75808, n75809, n75810,
    n75811, n75812, n75813, n75814, n75815, n75816, n75817, n75818, n75819,
    n75820, n75821, n75822, n75823, n75824, n75825, n75826, n75827, n75828,
    n75829, n75831, n75832, n75833, n75834, n75835, n75836, n75837, n75838,
    n75839, n75840, n75841, n75842, n75843, n75844, n75845, n75846, n75847,
    n75848, n75849, n75850, n75851, n75852, n75853, n75854, n75855, n75856,
    n75857, n75859, n75860, n75861, n75862, n75863, n75864, n75865, n75866,
    n75867, n75868, n75869, n75870, n75871, n75872, n75873, n75874, n75875,
    n75876, n75877, n75878, n75879, n75880, n75881, n75882, n75883, n75885,
    n75886, n75887, n75888, n75889, n75890, n75891, n75892, n75893, n75894,
    n75895, n75896, n75897, n75898, n75899, n75900, n75901, n75902, n75903,
    n75904, n75905, n75906, n75907, n75908, n75909, n75910, n75911, n75913,
    n75914, n75915, n75916, n75917, n75918, n75919, n75920, n75921, n75922,
    n75923, n75924, n75925, n75926, n75927, n75928, n75929, n75930, n75931,
    n75932, n75933, n75934, n75935, n75936, n75937, n75939, n75940, n75941,
    n75942, n75943, n75944, n75945, n75946, n75947, n75948, n75949, n75950,
    n75951, n75952, n75953, n75954, n75955, n75956, n75957, n75958, n75959,
    n75960, n75961, n75962, n75963, n75964, n75965, n75967, n75968, n75969,
    n75970, n75971, n75972, n75973, n75974, n75975, n75976, n75977, n75978,
    n75979, n75980, n75981, n75982, n75983, n75984, n75985, n75986, n75987,
    n75988, n75989, n75990, n75991, n75993, n75994, n75995, n75996, n75997,
    n75998, n75999, n76000, n76001, n76002, n76003, n76004, n76005, n76006,
    n76007, n76008, n76009, n76010, n76011, n76012, n76013, n76014, n76015,
    n76016, n76017, n76018, n76020, n76021, n76022, n76023, n76024, n76025,
    n76026, n76027, n76028, n76029, n76030, n76031, n76032, n76033, n76034,
    n76035, n76036, n76037, n76038, n76039, n76040, n76041, n76042, n76043,
    n76045, n76046, n76047, n76048, n76049, n76050, n76051, n76052, n76053,
    n76054, n76055, n76056, n76057, n76058, n76059, n76060, n76061, n76062,
    n76063, n76064, n76065, n76066, n76067, n76068, n76069, n76070, n76072,
    n76073, n76074, n76075, n76076, n76077, n76078, n76079, n76080, n76081,
    n76082, n76083, n76084, n76085, n76086, n76087, n76088, n76089, n76090,
    n76091, n76092, n76093, n76094, n76095, n76097, n76098, n76099, n76100,
    n76101, n76102, n76103, n76104, n76105, n76106, n76107, n76108, n76109,
    n76110, n76111, n76112, n76113, n76114, n76115, n76116, n76117, n76118,
    n76119, n76120, n76121, n76122, n76124, n76125, n76126, n76127, n76128,
    n76129, n76130, n76131, n76132, n76133, n76134, n76135, n76136, n76137,
    n76138, n76139, n76140, n76141, n76142, n76143, n76144, n76145, n76146,
    n76147, n76149, n76150, n76151, n76152, n76153, n76154, n76155, n76156,
    n76157, n76158, n76159, n76160, n76161, n76162, n76163, n76164, n76165,
    n76166, n76167, n76168, n76169, n76170, n76171, n76172, n76173, n76174,
    n76176, n76177, n76178, n76179, n76180, n76181, n76182, n76183, n76184,
    n76185, n76186, n76187, n76188, n76189, n76190, n76191, n76192, n76193,
    n76194, n76195, n76196, n76197, n76198, n76199, n76201, n76202, n76203,
    n76204, n76205, n76206, n76207, n76208, n76209, n76210, n76211, n76212,
    n76213, n76214, n76215, n76216, n76217, n76218, n76219, n76220, n76221,
    n76222, n76223, n76224, n76225, n76226, n76228, n76229, n76230, n76231,
    n76232, n76233, n76234, n76235, n76236, n76237, n76238, n76239, n76240,
    n76241, n76242, n76243, n76244, n76245, n76246, n76247, n76248, n76249,
    n76250, n76251, n76253, n76254, n76255, n76256, n76257, n76258, n76259,
    n76260, n76261, n76262, n76263, n76264, n76265, n76266, n76267, n76268,
    n76269, n76270, n76271, n76272, n76273, n76274, n76275, n76276, n76278,
    n76279, n76280, n76281, n76282, n76283, n76284, n76285, n76286, n76287,
    n76288, n76289, n76290, n76291, n76292, n76293, n76294, n76295, n76296,
    n76297, n76298, n76299, n76300, n76301, n76302, n76303, n76305, n76306,
    n76307, n76308, n76309, n76310, n76311, n76312, n76313, n76314, n76315,
    n76316, n76317, n76318, n76319, n76320, n76321, n76322, n76323, n76324,
    n76325, n76326, n76327, n76328, n76329, n76330, n76331, n76332, n76333,
    n76334, n76335, n76336, n76337, n76338, n76339, n76340, n76341, n76342,
    n76344, n76345, n76346, n76347, n76348, n76349, n76350, n76351, n76353,
    n76354, n76355, n76357, n76358, n76359, n76361, n76362, n76364, n76365,
    n76366, n76368, n76369, n76371, n76372, n76373, n76374, n76376, n76377,
    n76378, n76379, n76380, n76381, n76382, n76383, n76384, n76385, n76386,
    n76387, n76388, n76389, n76390, n76392, n76393, n76394, n76396, n76397,
    n76399, n76400, n76401, n76403, n76405, n76406, n76407, n76408, n76409,
    n76411, n76412, n76413, n76415, n76416, n76417, n76419, n76420, n76422,
    n76423, n76425, n76426, n76428, n76429, n76430, n76431, n76432, n76433,
    n76435, n76436, n76437, n76438, n76440, n76441, n76442, n76443, n76445,
    n76446, n76447, n76448, n76450, n76451, n76452, n76453, n76455, n76456,
    n76457, n76458, n76460, n76461, n76462, n76463, n76465, n76466, n76467,
    n76468, n76470, n76471, n76472, n76473, n76475, n76476, n76477, n76478,
    n76480, n76481, n76482, n76483, n76485, n76486, n76487, n76488, n76490,
    n76491, n76492, n76493, n76495, n76496, n76497, n76498, n76500, n76501,
    n76502, n76503, n76505, n76506, n76507, n76508, n76510, n76511, n76512,
    n76513, n76515, n76516, n76517, n76518, n76520, n76521, n76522, n76523,
    n76525, n76526, n76527, n76528, n76530, n76531, n76532, n76533, n76535,
    n76536, n76537, n76538, n76540, n76541, n76542, n76543, n76545, n76546,
    n76547, n76548, n76550, n76551, n76552, n76553, n76555, n76556, n76557,
    n76558, n76560, n76561, n76562, n76563, n76565, n76566, n76567, n76568,
    n76570, n76571, n76572, n76573, n76575, n76576, n76577, n76578, n76580,
    n76581, n76582, n76583, n76584, n76585, n76586, n76587, n76588, n76589,
    n76590, n76591, n76592, n76593, n76594, n76595, n76596, n76597, n76598,
    n76599, n76600, n76601, n76602, n76603, n76605, n76606, n76607, n76608,
    n76609, n76610, n76611, n76612, n76613, n76614, n76615, n76616, n76617,
    n76619, n76620, n76621, n76622, n76623, n76624, n76625, n76626, n76627,
    n76629, n76630, n76631, n76632, n76633, n76634, n76636, n76637, n76669,
    n76670, n76671, n76672, n76673, n76674, n76675, n76676, n76677, n76678,
    n76679, n76680, n76681, n76682, n76683, n76684, n76685, n76686, n76687,
    n76688, n76689, n76690, n76691, n76692, n76693, n76694, n76695, n76696,
    n76697, n76698, n76699, n76700, n76701, n76702, n76703, n76704, n76705,
    n76706, n76707, n76708, n76709, n76710, n76711, n76712, n76713, n76714,
    n76715, n76716, n76717, n76718, n76719, n76720, n76721, n76722, n76723,
    n76724, n76725, n76726, n76727, n76728, n76729, n76730, n76731, n76732,
    n76733, n76734, n76735, n76736, n76737, n76738, n76739, n76740, n76741,
    n76742, n76743, n76744, n76745, n76746, n76747, n76748, n76749, n76750,
    n76751, n76752, n76753, n76754, n76755, n76756, n76757, n76758, n76759,
    n76760, n76761, n76762, n76763, n76764, n76765, n76766, n76767, n76768,
    n76769, n76770, n76771, n76772, n76773, n76774, n76775, n76776, n76777,
    n76778, n76779, n76780, n76781, n76782, n76783, n76784, n76785, n76786,
    n76787, n76788, n76789, n76790, n76791, n76792, n76793, n76794, n76795,
    n76796, n76797, n76798, n76799, n76800, n76801, n76802, n76803, n76804,
    n76805, n76806, n76807, n76808, n76809, n76810, n76811, n76812, n76813,
    n76814, n76815, n76816, n76817, n76818, n76819, n76820, n76821, n76822,
    n76823, n76824, n76825, n76826, n76827, n76828, n76829, n76830, n76831,
    n76832, n76833, n76834, n76835, n76836, n76837, n76838, n76839, n76840,
    n76841, n76842, n76843, n76844, n76845, n76846, n76847, n76848, n76849,
    n76850, n76851, n76852, n76853, n76854, n76855, n76856, n76857, n76858,
    n76859, n76860, n76861, n76862, n76863, n76864, n76865, n76866, n76867,
    n76868, n76869, n76870, n76871, n76872, n76873, n76874, n76875, n76876,
    n76877, n76878, n76879, n76880, n76881, n76882, n76883, n76884, n76885,
    n76886, n76887, n76888, n76889, n76890, n76891, n76892, n76893, n76894,
    n76895, n76896, n76897, n76898, n76899, n76900, n76901, n76902, n76903,
    n76904, n76905, n76906, n76907, n76908, n76909, n76910, n76911, n76912,
    n76913, n76914, n76915, n76916, n76917, n76918, n76919, n76920, n76921,
    n76922, n76923, n76924, n76925, n76926, n76927, n76928, n76929, n76930,
    n76931, n76932, n76933, n76934, n76935, n76936, n76937, n76938, n76939,
    n76940, n76941, n76942, n76943, n76944, n76945, n76946, n76947, n76948,
    n76949, n76950, n76951, n76952, n76953, n76954, n76955, n76956, n76957,
    n76958, n76959, n76960, n76961, n76962, n76963, n76964, n76965, n76966,
    n76967, n76968, n76969, n76970, n76971, n76972, n76973, n76974, n76975,
    n76976, n76977, n76978, n76979, n76980, n76981, n76982, n76983, n76984,
    n76985, n76986, n76987, n76988, n76989, n76990, n76991, n76992, n76993,
    n76994, n76995, n76996, n76997, n76998, n76999, n77000, n77001, n77002,
    n77003, n77004, n77005, n77006, n77007, n77008, n77009, n77010, n77011,
    n77012, n77013, n77014, n77015, n77016, n77017, n77018, n77019, n77020,
    n77021, n77022, n77023, n77024, n77025, n77026, n77027, n77028, n77029,
    n77030, n77031, n77032, n77033, n77034, n77035, n77036, n77037, n77038,
    n77039, n77040, n77041, n77042, n77043, n77044, n77045, n77046, n77047,
    n77048, n77049, n77050, n77051, n77052, n77053, n77054, n77055, n77056,
    n77057, n77058, n77059, n77060, n77061, n77062, n77063, n77064, n77065,
    n77066, n77067, n77068, n77069, n77070, n77071, n77072, n77073, n77074,
    n77075, n77076, n77077, n77078, n77079, n77080, n77081, n77082, n77083,
    n77084, n77085, n77086, n77087, n77088, n77089, n77090, n77091, n77092,
    n77093, n77094, n77095, n77096, n77097, n77098, n77099, n77100, n77101,
    n77102, n77103, n77104, n77105, n77106, n77107, n77108, n77109, n77110,
    n77111, n77112, n77113, n77114, n77115, n77116, n77117, n77118, n77119,
    n77120, n77121, n77122, n77123, n77124, n77125, n77126, n77127, n77128,
    n77129, n77130, n77131, n77132, n77133, n77134, n77135, n77136, n77137,
    n77138, n77139, n77140, n77141, n77142, n77143, n77144, n77145, n77146,
    n77147, n77148, n77149, n77150, n77151, n77152, n77153, n77154, n77155,
    n77156, n77157, n77158, n77159, n77160, n77161, n77162, n77163, n77164,
    n77165, n77166, n77167, n77168, n77169, n77170, n77171, n77172, n77173,
    n77174, n77175, n77176, n77177, n77178, n77179, n77180, n77181, n77182,
    n77183, n77184, n77185, n77186, n77187, n77188, n77189, n77190, n77191,
    n77192, n77193, n77194, n77195, n77196, n77197, n77198, n77199, n77200,
    n77201, n77202, n77203, n77204, n77205, n77206, n77207, n77208, n77209,
    n77210, n77211, n77212, n77213, n77214, n77215, n77216, n77217, n77218,
    n77219, n77220, n77221, n77222, n77223, n77224, n77225, n77226, n77227,
    n77228, n77229, n77230, n77231, n77232, n77233, n77234, n77235, n77236,
    n77237, n77238, n77239, n77240, n77241, n77242, n77243, n77244, n77245,
    n77246, n77247, n77248, n77249, n77250, n77251, n77252, n77253, n77254,
    n77255, n77256, n77257, n77258, n77259, n77260, n77261, n77262, n77263,
    n77264, n77265, n77266, n77267, n77268, n77269, n77270, n77271, n77272,
    n77273, n77274, n77275, n77276, n77277, n77278, n77279, n77280, n77281,
    n77282, n77283, n77284, n77285, n77286, n77287, n77288, n77289, n77290,
    n77291, n77292, n77293, n77294, n77295, n77296, n77297, n77298, n77299,
    n77300, n77302, n77303, n77304, n77305, n77306, n77307, n77308, n77309,
    n77311, n77312, n77313, n77314, n77315, n77316, n77317, n77318, n77319,
    n77320, n77321, n77322, n77323, n77324, n77326, n77327, n77328, n77329,
    n77330, n77331, n77332, n77333, n77334, n77335, n77336, n77337, n77338,
    n77339, n77340, n77341, n77342, n77343, n77344, n77345, n77346, n77347,
    n77348, n77349, n77350, n77351, n77352, n77353, n77354, n77355, n77356,
    n77357, n77358, n77359, n77360, n77361, n77362, n77363, n77364, n77365,
    n77367, n77368, n77369, n77370, n77371, n77372, n77373, n77374, n77375,
    n77376, n77377, n77378, n77379, n77380, n77381, n77382, n77383, n77384,
    n77385, n77386, n77387, n77388, n77389, n77390, n77391, n77392, n77393,
    n77394, n77395, n77396, n77397, n77398, n77399, n77400, n77401, n77402,
    n77403, n77404, n77405, n77406, n77407, n77408, n77409, n77410, n77411,
    n77412, n77413, n77414, n77415, n77416, n77417, n77418, n77419, n77420,
    n77421, n77422, n77423, n77424, n77425, n77426, n77427, n77428, n77429,
    n77430, n77431, n77432, n77433, n77434, n77435, n77436, n77437, n77438,
    n77439, n77440, n77441, n77442, n77443, n77444, n77445, n77446, n77447,
    n77448, n77449, n77450, n77451, n77452, n77453, n77454, n77455, n77456,
    n77457, n77458, n77459, n77460, n77461, n77462, n77463, n77464, n77465,
    n77466, n77467, n77468, n77469, n77470, n77471, n77472, n77473, n77474,
    n77475, n77476, n77477, n77478, n77479, n77480, n77481, n77482, n77483,
    n77484, n77485, n77486, n77487, n77488, n77489, n77490, n77491, n77492,
    n77493, n77494, n77495, n77496, n77497, n77498, n77499, n77500, n77501,
    n77502, n77503, n77504, n77505, n77506, n77507, n77508, n77509, n77510,
    n77511, n77512, n77513, n77514, n77515, n77516, n77517, n77518, n77519,
    n77520, n77521, n77522, n77523, n77524, n77525, n77526, n77527, n77528,
    n77529, n77530, n77531, n77532, n77533, n77534, n77535, n77536, n77537,
    n77538, n77539, n77540, n77541, n77542, n77543, n77544, n77545, n77546,
    n77547, n77548, n77549, n77550, n77551, n77552, n77553, n77554, n77555,
    n77556, n77557, n77558, n77559, n77560, n77561, n77562, n77563, n77564,
    n77565, n77566, n77567, n77568, n77569, n77570, n77571, n77572, n77573,
    n77574, n77575, n77576, n77577, n77578, n77579, n77580, n77581, n77582,
    n77583, n77584, n77585, n77586, n77587, n77588, n77589, n77590, n77591,
    n77592, n77593, n77594, n77595, n77596, n77597, n77598, n77599, n77600,
    n77601, n77602, n77603, n77604, n77605, n77606, n77607, n77608, n77609,
    n77610, n77611, n77612, n77613, n77614, n77615, n77616, n77617, n77618,
    n77619, n77620, n77621, n77622, n77623, n77624, n77625, n77626, n77627,
    n77628, n77629, n77630, n77631, n77632, n77633, n77634, n77635, n77636,
    n77637, n77638, n77639, n77640, n77641, n77642, n77643, n77644, n77645,
    n77646, n77647, n77648, n77649, n77650, n77651, n77652, n77653, n77654,
    n77655, n77656, n77657, n77658, n77659, n77660, n77661, n77662, n77663,
    n77664, n77665, n77666, n77667, n77668, n77669, n77670, n77671, n77672,
    n77673, n77674, n77675, n77676, n77677, n77678, n77679, n77680, n77681,
    n77682, n77683, n77684, n77685, n77686, n77687, n77688, n77689, n77690,
    n77691, n77692, n77693, n77694, n77695, n77696, n77697, n77698, n77699,
    n77700, n77701, n77702, n77703, n77704, n77705, n77706, n77707, n77708,
    n77709, n77710, n77711, n77712, n77713, n77714, n77715, n77716, n77717,
    n77718, n77719, n77720, n77721, n77722, n77723, n77724, n77725, n77726,
    n77727, n77728, n77729, n77730, n77731, n77732, n77733, n77734, n77735,
    n77736, n77737, n77738, n77739, n77740, n77741, n77742, n77743, n77744,
    n77745, n77746, n77747, n77748, n77749, n77750, n77751, n77752, n77753,
    n77754, n77755, n77756, n77757, n77758, n77759, n77760, n77761, n77762,
    n77763, n77764, n77765, n77766, n77767, n77768, n77769, n77770, n77771,
    n77772, n77773, n77774, n77775, n77776, n77777, n77778, n77779, n77780,
    n77781, n77782, n77783, n77784, n77785, n77786, n77787, n77788, n77789,
    n77790, n77791, n77792, n77793, n77794, n77795, n77796, n77797, n77798,
    n77799, n77800, n77801, n77802, n77803, n77804, n77805, n77806, n77807,
    n77808, n77809, n77810, n77811, n77812, n77813, n77814, n77815, n77816,
    n77817, n77818, n77819, n77820, n77821, n77822, n77823, n77824, n77825,
    n77826, n77827, n77828, n77829, n77830, n77831, n77832, n77833, n77834,
    n77835, n77836, n77837, n77838, n77839, n77840, n77841, n77842, n77843,
    n77844, n77845, n77846, n77847, n77848, n77849, n77850, n77851, n77852,
    n77853, n77854, n77855, n77856, n77857, n77858, n77859, n77860, n77861,
    n77862, n77863, n77864, n77865, n77866, n77867, n77868, n77869, n77870,
    n77871, n77872, n77873, n77874, n77875, n77876, n77877, n77878, n77879,
    n77880, n77881, n77882, n77883, n77884, n77885, n77886, n77887, n77888,
    n77889, n77890, n77891, n77892, n77893, n77894, n77895, n77896, n77897,
    n77898, n77899, n77900, n77901, n77902, n77903, n77904, n77905, n77906,
    n77907, n77908, n77909, n77910, n77911, n77912, n77913, n77914, n77915,
    n77916, n77917, n77918, n77919, n77920, n77921, n77922, n77923, n77924,
    n77925, n77926, n77927, n77928, n77929, n77930, n77931, n77932, n77933,
    n77934, n77935, n77936, n77937, n77938, n77939, n77940, n77941, n77942,
    n77943, n77944, n77945, n77946, n77947, n77948, n77949, n77950, n77951,
    n77952, n77953, n77954, n77955, n77956, n77957, n77958, n77959, n77960,
    n77961, n77962, n77963, n77964, n77965, n77966, n77967, n77968, n77969,
    n77970, n77971, n77972, n77973, n77974, n77975, n77976, n77977, n77978,
    n77979, n77980, n77981, n77982, n77983, n77984, n77985, n77986, n77987,
    n77988, n77989, n77990, n77991, n77992, n77993, n77994, n77995, n77996,
    n77997, n77998, n77999, n78000, n78001, n78002, n78003, n78004, n78005,
    n78006, n78007, n78008, n78009, n78010, n78011, n78012, n78013, n78014,
    n78015, n78016, n78017, n78018, n78019, n78020, n78021, n78022, n78023,
    n78024, n78025, n78026, n78027, n78028, n78029, n78030, n78031, n78032,
    n78033, n78034, n78035, n78036, n78037, n78038, n78039, n78040, n78041,
    n78042, n78043, n78044, n78045, n78046, n78047, n78048, n78049, n78050,
    n78051, n78052, n78053, n78054, n78055, n78056, n78057, n78058, n78059,
    n78060, n78061, n78062, n78063, n78064, n78065, n78066, n78067, n78068,
    n78069, n78070, n78071, n78072, n78073, n78074, n78075, n78076, n78077,
    n78078, n78079, n78080, n78081, n78082, n78083, n78084, n78085, n78086,
    n78087, n78088, n78089, n78090, n78091, n78092, n78093, n78094, n78095,
    n78096, n78097, n78098, n78099, n78100, n78101, n78102, n78103, n78104,
    n78105, n78106, n78107, n78108, n78109, n78110, n78111, n78112, n78113,
    n78114, n78115, n78116, n78117, n78118, n78119, n78120, n78121, n78122,
    n78123, n78124, n78125, n78126, n78127, n78128, n78129, n78130, n78131,
    n78132, n78133, n78134, n78135, n78136, n78137, n78138, n78139, n78140,
    n78141, n78142, n78143, n78144, n78145, n78146, n78147, n78148, n78149,
    n78150, n78151, n78152, n78153, n78154, n78155, n78156, n78157, n78158,
    n78159, n78160, n78161, n78162, n78163, n78164, n78165, n78166, n78167,
    n78168, n78169, n78170, n78171, n78172, n78173, n78174, n78175, n78176,
    n78177, n78178, n78179, n78180, n78181, n78182, n78183, n78184, n78185,
    n78186, n78187, n78188, n78189, n78190, n78191, n78192, n78193, n78194,
    n78195, n78196, n78197, n78198, n78199, n78200, n78201, n78202, n78203,
    n78204, n78205, n78206, n78207, n78208, n78209, n78210, n78211, n78212,
    n78213, n78214, n78215, n78216, n78217, n78218, n78219, n78220, n78221,
    n78222, n78223, n78224, n78225, n78226, n78227, n78228, n78229, n78230,
    n78231, n78232, n78233, n78234, n78235, n78236, n78237, n78238, n78239,
    n78240, n78241, n78242, n78243, n78244, n78245, n78246, n78247, n78248,
    n78249, n78250, n78251, n78252, n78253, n78254, n78255, n78256, n78257,
    n78258, n78259, n78260, n78261, n78262, n78263, n78264, n78265, n78266,
    n78267, n78268, n78269, n78270, n78271, n78272, n78273, n78274, n78275,
    n78276, n78277, n78278, n78279, n78280, n78281, n78282, n78283, n78284,
    n78285, n78286, n78287, n78288, n78289, n78290, n78291, n78292, n78293,
    n78294, n78295, n78296, n78297, n78298, n78299, n78300, n78301, n78302,
    n78303, n78304, n78305, n78306, n78307, n78308, n78309, n78310, n78311,
    n78312, n78313, n78314, n78315, n78316, n78317, n78318, n78319, n78320,
    n78321, n78322, n78323, n78324, n78325, n78326, n78327, n78328, n78329,
    n78330, n78331, n78332, n78333, n78334, n78335, n78336, n78337, n78338,
    n78339, n78340, n78341, n78342, n78343, n78344, n78345, n78346, n78347,
    n78348, n78349, n78350, n78351, n78352, n78353, n78354, n78355, n78356,
    n78357, n78358, n78359, n78360, n78361, n78362, n78363, n78364, n78365,
    n78366, n78367, n78368, n78369, n78370, n78371, n78372, n78373, n78374,
    n78375, n78376, n78377, n78378, n78379, n78380, n78381, n78382, n78383,
    n78384, n78385, n78386, n78387, n78388, n78389, n78390, n78391, n78392,
    n78393, n78394, n78395, n78396, n78397, n78398, n78399, n78400, n78401,
    n78402, n78403, n78404, n78405, n78406, n78407, n78408, n78409, n78410,
    n78411, n78412, n78413, n78414, n78415, n78416, n78417, n78418, n78419,
    n78420, n78421, n78422, n78423, n78424, n78425, n78426, n78427, n78428,
    n78429, n78430, n78431, n78432, n78433, n78434, n78435, n78436, n78437,
    n78438, n78439, n78440, n78441, n78442, n78443, n78444, n78445, n78446,
    n78447, n78448, n78449, n78450, n78451, n78452, n78453, n78454, n78455,
    n78456, n78457, n78458, n78459, n78460, n78461, n78462, n78463, n78464,
    n78465, n78466, n78467, n78468, n78469, n78470, n78471, n78472, n78473,
    n78474, n78475, n78476, n78477, n78478, n78479, n78480, n78481, n78482,
    n78483, n78484, n78485, n78486, n78487, n78488, n78489, n78490, n78491,
    n78492, n78493, n78494, n78495, n78496, n78497, n78498, n78499, n78500,
    n78501, n78502, n78503, n78504, n78505, n78506, n78507, n78508, n78509,
    n78510, n78511, n78512, n78513, n78514, n78515, n78516, n78517, n78518,
    n78519, n78520, n78521, n78522, n78523, n78524, n78525, n78526, n78527,
    n78528, n78529, n78530, n78531, n78532, n78533, n78534, n78535, n78536,
    n78537, n78538, n78539, n78540, n78541, n78542, n78543, n78544, n78545,
    n78546, n78547, n78548, n78549, n78550, n78551, n78552, n78553, n78554,
    n78555, n78556, n78557, n78558, n78559, n78560, n78561, n78562, n78563,
    n78564, n78565, n78566, n78567, n78568, n78569, n78570, n78571, n78572,
    n78573, n78574, n78575, n78576, n78577, n78578, n78579, n78580, n78581,
    n78582, n78583, n78584, n78585, n78586, n78587, n78588, n78589, n78590,
    n78591, n78592, n78593, n78594, n78595, n78596, n78597, n78598, n78599,
    n78600, n78601, n78602, n78603, n78604, n78605, n78606, n78607, n78608,
    n78609, n78610, n78611, n78612, n78613, n78614, n78615, n78616, n78617,
    n78618, n78619, n78620, n78621, n78622, n78623, n78624, n78625, n78626,
    n78627, n78628, n78629, n78630, n78631, n78632, n78633, n78634, n78635,
    n78636, n78637, n78638, n78639, n78640, n78641, n78642, n78643, n78644,
    n78645, n78646, n78647, n78648, n78649, n78650, n78651, n78652, n78653,
    n78654, n78655, n78656, n78657, n78658, n78659, n78660, n78661, n78662,
    n78663, n78664, n78665, n78666, n78667, n78668, n78669, n78670, n78671,
    n78672, n78673, n78674, n78675, n78676, n78677, n78678, n78679, n78680,
    n78681, n78682, n78683, n78684, n78685, n78686, n78687, n78688, n78689,
    n78690, n78691, n78692, n78693, n78694, n78695, n78696, n78697, n78698,
    n78699, n78700, n78701, n78702, n78703, n78704, n78705, n78706, n78707,
    n78708, n78709, n78710, n78711, n78712, n78713, n78714, n78715, n78716,
    n78717, n78718, n78719, n78720, n78721, n78722, n78723, n78724, n78725,
    n78726, n78727, n78728, n78729, n78730, n78731, n78732, n78733, n78734,
    n78735, n78736, n78737, n78738, n78739, n78740, n78741, n78742, n78743,
    n78744, n78745, n78746, n78747, n78748, n78749, n78750, n78751, n78752,
    n78753, n78754, n78755, n78756, n78757, n78758, n78759, n78760, n78761,
    n78762, n78763, n78764, n78765, n78766, n78767, n78768, n78769, n78770,
    n78771, n78772, n78773, n78774, n78775, n78776, n78777, n78778, n78779,
    n78780, n78781, n78782, n78783, n78784, n78785, n78786, n78787, n78788,
    n78789, n78790, n78791, n78792, n78793, n78794, n78795, n78796, n78797,
    n78798, n78799, n78800, n78801, n78802, n78803, n78804, n78805, n78806,
    n78807, n78808, n78809, n78810, n78811, n78812, n78813, n78814, n78815,
    n78816, n78817, n78818, n78819, n78820, n78821, n78822, n78823, n78824,
    n78825, n78826, n78827, n78828, n78829, n78830, n78831, n78832, n78833,
    n78834, n78835, n78836, n78837, n78838, n78839, n78840, n78841, n78842,
    n78843, n78844, n78845, n78846, n78847, n78848, n78849, n78850, n78851,
    n78852, n78853, n78854, n78855, n78856, n78857, n78858, n78859, n78860,
    n78861, n78862, n78863, n78864, n78865, n78866, n78867, n78868, n78869,
    n78870, n78871, n78872, n78873, n78874, n78875, n78876, n78877, n78878,
    n78879, n78880, n78881, n78882, n78883, n78884, n78885, n78886, n78887,
    n78888, n78889, n78890, n78891, n78892, n78893, n78894, n78895, n78896,
    n78897, n78898, n78899, n78900, n78901, n78902, n78903, n78904, n78905,
    n78906, n78907, n78908, n78909, n78910, n78911, n78912, n78913, n78914,
    n78915, n78916, n78917, n78918, n78919, n78920, n78921, n78922, n78923,
    n78924, n78925, n78926, n78927, n78928, n78929, n78930, n78931, n78932,
    n78933, n78934, n78935, n78936, n78937, n78938, n78939, n78940, n78941,
    n78942, n78943, n78944, n78945, n78946, n78947, n78948, n78949, n78950,
    n78951, n78952, n78953, n78954, n78955, n78956, n78957, n78958, n78959,
    n78960, n78961, n78962, n78963, n78964, n78965, n78966, n78967, n78968,
    n78969, n78970, n78971, n78972, n78973, n78974, n78975, n78976, n78977,
    n78978, n78979, n78980, n78981, n78982, n78983, n78984, n78985, n78986,
    n78987, n78988, n78989, n78990, n78991, n78992, n78993, n78994, n78995,
    n78996, n78997, n78998, n78999, n79000, n79001, n79002, n79003, n79004,
    n79005, n79006, n79007, n79008, n79009, n79010, n79011, n79012, n79013,
    n79014, n79015, n79016, n79017, n79018, n79019, n79020, n79021, n79022,
    n79023, n79024, n79025, n79026, n79027, n79028, n79029, n79030, n79031,
    n79032, n79033, n79034, n79035, n79036, n79037, n79038, n79039, n79040,
    n79041, n79042, n79043, n79044, n79045, n79046, n79047, n79048, n79049,
    n79050, n79051, n79052, n79053, n79054, n79055, n79056, n79057, n79058,
    n79059, n79060, n79061, n79062, n79063, n79064, n79065, n79066, n79067,
    n79068, n79069, n79070, n79071, n79072, n79073, n79074, n79075, n79076,
    n79077, n79078, n79079, n79080, n79081, n79082, n79083, n79084, n79085,
    n79086, n79087, n79088, n79089, n79090, n79091, n79092, n79093, n79094,
    n79095, n79096, n79097, n79098, n79099, n79100, n79101, n79102, n79103,
    n79104, n79105, n79106, n79107, n79108, n79109, n79110, n79111, n79112,
    n79113, n79114, n79115, n79116, n79117, n79118, n79119, n79120, n79121,
    n79122, n79123, n79124, n79125, n79126, n79127, n79128, n79129, n79130,
    n79131, n79132, n79133, n79134, n79135, n79136, n79137, n79138, n79139,
    n79140, n79141, n79142, n79143, n79144, n79145, n79146, n79147, n79148,
    n79149, n79150, n79151, n79152, n79153, n79154, n79155, n79156, n79157,
    n79158, n79159, n79160, n79161, n79162, n79163, n79164, n79165, n79166,
    n79167, n79168, n79169, n79170, n79171, n79172, n79173, n79174, n79175,
    n79176, n79177, n79178, n79179, n79180, n79181, n79182, n79183, n79184,
    n79185, n79186, n79187, n79188, n79189, n79190, n79191, n79192, n79193,
    n79194, n79195, n79196, n79197, n79198, n79199, n79200, n79201, n79202,
    n79203, n79204, n79205, n79206, n79207, n79208, n79209, n79210, n79211,
    n79212, n79213, n79214, n79215, n79216, n79217, n79218, n79219, n79220,
    n79221, n79222, n79223, n79224, n79225, n79226, n79227, n79228, n79229,
    n79230, n79231, n79232, n79233, n79234, n79235, n79236, n79237, n79238,
    n79239, n79240, n79241, n79242, n79243, n79244, n79245, n79246, n79247,
    n79248, n79249, n79250, n79251, n79252, n79253, n79254, n79255, n79256,
    n79257, n79258, n79259, n79260, n79261, n79262, n79263, n79264, n79265,
    n79266, n79267, n79268, n79269, n79270, n79271, n79272, n79273, n79274,
    n79275, n79276, n79277, n79278, n79279, n79280, n79281, n79282, n79283,
    n79284, n79285, n79286, n79287, n79288, n79289, n79290, n79291, n79292,
    n79293, n79294, n79295, n79296, n79297, n79298, n79299, n79300, n79301,
    n79302, n79303, n79304, n79305, n79306, n79307, n79308, n79309, n79310,
    n79311, n79312, n79313, n79314, n79315, n79316, n79317, n79318, n79319,
    n79320, n79321, n79322, n79323, n79324, n79325, n79326, n79327, n79328,
    n79329, n79330, n79331, n79332, n79333, n79334, n79335, n79336, n79337,
    n79338, n79339, n79340, n79341, n79342, n79343, n79344, n79345, n79346,
    n79347, n79348, n79349, n79350, n79351, n79352, n79353, n79354, n79355,
    n79356, n79357, n79358, n79359, n79360, n79361, n79362, n79363, n79364,
    n79365, n79366, n79367, n79368, n79369, n79370, n79371, n79372, n79373,
    n79374, n79375, n79376, n79377, n79378, n79379, n79380, n79381, n79382,
    n79383, n79384, n79385, n79386, n79387, n79388, n79389, n79390, n79391,
    n79392, n79393, n79394, n79395, n79396, n79397, n79398, n79399, n79400,
    n79401, n79402, n79403, n79404, n79405, n79406, n79407, n79408, n79409,
    n79410, n79411, n79412, n79413, n79414, n79415, n79416, n79417, n79418,
    n79419, n79420, n79421, n79422, n79423, n79424, n79425, n79426, n79427,
    n79428, n79429, n79430, n79431, n79432, n79433, n79434, n79435, n79436,
    n79437, n79438, n79439, n79440, n79441, n79442, n79443, n79444, n79445,
    n79446, n79447, n79448, n79449, n79450, n79451, n79452, n79453, n79454,
    n79455, n79456, n79457, n79458, n79459, n79460, n79461, n79462, n79463,
    n79464, n79465, n79466, n79467, n79468, n79469, n79470, n79471, n79472,
    n79473, n79474, n79475, n79476, n79477, n79478, n79479, n79480, n79481,
    n79482, n79483, n79484, n79485, n79486, n79487, n79488, n79489, n79490,
    n79491, n79492, n79493, n79494, n79495, n79496, n79497, n79498, n79499,
    n79500, n79501, n79502, n79503, n79504, n79505, n79506, n79507, n79508,
    n79509, n79510, n79511, n79512, n79513, n79514, n79515, n79516, n79517,
    n79518, n79519, n79520, n79521, n79522, n79523, n79524, n79525, n79526,
    n79527, n79528, n79529, n79530, n79531, n79532, n79533, n79534, n79535,
    n79536, n79537, n79538, n79539, n79540, n79541, n79542, n79543, n79544,
    n79545, n79546, n79547, n79548, n79549, n79550, n79551, n79552, n79553,
    n79554, n79555, n79556, n79557, n79558, n79559, n79560, n79561, n79562,
    n79563, n79564, n79565, n79566, n79567, n79568, n79569, n79570, n79571,
    n79572, n79573, n79574, n79575, n79576, n79577, n79578, n79579, n79580,
    n79581, n79582, n79583, n79584, n79585, n79586, n79587, n79588, n79589,
    n79590, n79591, n79592, n79593, n79594, n79595, n79596, n79597, n79598,
    n79599, n79600, n79601, n79602, n79603, n79604, n79605, n79606, n79607,
    n79608, n79609, n79610, n79611, n79612, n79613, n79614, n79615, n79616,
    n79617, n79618, n79619, n79620, n79621, n79622, n79623, n79624, n79625,
    n79626, n79627, n79628, n79629, n79630, n79631, n79632, n79633, n79634,
    n79635, n79636, n79637, n79638, n79639, n79640, n79641, n79642, n79643,
    n79644, n79645, n79646, n79647, n79648, n79649, n79650, n79651, n79652,
    n79653, n79654, n79655, n79656, n79657, n79658, n79659, n79660, n79661,
    n79662, n79663, n79664, n79665, n79666, n79667, n79668, n79669, n79670,
    n79671, n79672, n79673, n79674, n79675, n79676, n79677, n79678, n79679,
    n79680, n79681, n79682, n79683, n79684, n79685, n79686, n79687, n79688,
    n79689, n79690, n79691, n79692, n79693, n79694, n79695, n79696, n79697,
    n79698, n79699, n79700, n79701, n79702, n79703, n79704, n79705, n79706,
    n79707, n79708, n79709, n79710, n79711, n79712, n79713, n79714, n79715,
    n79716, n79717, n79718, n79719, n79720, n79721, n79722, n79723, n79724,
    n79725, n79726, n79727, n79728, n79729, n79730, n79731, n79732, n79733,
    n79734, n79735, n79736, n79737, n79738, n79739, n79740, n79741, n79742,
    n79743, n79744, n79745, n79746, n79747, n79748, n79749, n79750, n79751,
    n79752, n79753, n79754, n79755, n79756, n79757, n79758, n79759, n79760,
    n79761, n79762, n79763, n79764, n79765, n79766, n79767, n79768, n79769,
    n79770, n79771, n79772, n79773, n79774, n79775, n79776, n79777, n79778,
    n79779, n79780, n79781, n79782, n79783, n79784, n79785, n79786, n79787,
    n79788, n79789, n79790, n79791, n79792, n79793, n79794, n79795, n79796,
    n79797, n79798, n79799, n79800, n79801, n79802, n79803, n79804, n79805,
    n79806, n79807, n79808, n79809, n79810, n79811, n79812, n79813, n79814,
    n79815, n79816, n79817, n79818, n79819, n79820, n79821, n79822, n79823,
    n79824, n79825, n79826, n79827, n79828, n79829, n79830, n79831, n79832,
    n79833, n79834, n79835, n79836, n79837, n79838, n79839, n79840, n79841,
    n79842, n79843, n79844, n79845, n79846, n79847, n79848, n79849, n79850,
    n79851, n79852, n79853, n79854, n79855, n79856, n79857, n79858, n79859,
    n79860, n79861, n79862, n79863, n79864, n79865, n79866, n79867, n79868,
    n79869, n79870, n79871, n79872, n79873, n79874, n79875, n79876, n79877,
    n79878, n79879, n79880, n79881, n79882, n79883, n79884, n79885, n79886,
    n79887, n79888, n79889, n79890, n79891, n79892, n79893, n79894, n79895,
    n79896, n79897, n79898, n79899, n79900, n79901, n79902, n79903, n79904,
    n79905, n79906, n79907, n79908, n79909, n79910, n79911, n79912, n79913,
    n79914, n79915, n79916, n79917, n79918, n79919, n79920, n79921, n79922,
    n79923, n79924, n79925, n79926, n79927, n79928, n79929, n79930, n79931,
    n79932, n79933, n79934, n79935, n79936, n79937, n79938, n79939, n79940,
    n79941, n79942, n79943, n79944, n79945, n79946, n79947, n79948, n79949,
    n79950, n79951, n79952, n79953, n79954, n79955, n79956, n79957, n79958,
    n79959, n79960, n79961, n79962, n79963, n79964, n79965, n79966, n79967,
    n79968, n79969, n79970, n79971, n79972, n79973, n79974, n79975, n79976,
    n79977, n79978, n79979, n79980, n79981, n79982, n79983, n79984, n79985,
    n79986, n79987, n79988, n79989, n79990, n79991, n79992, n79993, n79994,
    n79995, n79996, n79997, n79998, n79999, n80000, n80001, n80002, n80003,
    n80004, n80005, n80006, n80007, n80008, n80009, n80010, n80011, n80012,
    n80013, n80014, n80015, n80016, n80017, n80018, n80019, n80020, n80021,
    n80022, n80023, n80024, n80025, n80026, n80027, n80028, n80029, n80030,
    n80031, n80032, n80033, n80034, n80035, n80036, n80037, n80038, n80039,
    n80040, n80041, n80042, n80043, n80044, n80045, n80046, n80047, n80048,
    n80049, n80050, n80051, n80052, n80053, n80054, n80055, n80056, n80057,
    n80058, n80059, n80060, n80061, n80062, n80063, n80064, n80065, n80066,
    n80067, n80068, n80069, n80070, n80071, n80072, n80073, n80074, n80075,
    n80076, n80077, n80078, n80079, n80080, n80081, n80082, n80083, n80084,
    n80085, n80086, n80087, n80088, n80089, n80090, n80091, n80092, n80093,
    n80094, n80095, n80096, n80097, n80098, n80099, n80100, n80101, n80102,
    n80103, n80104, n80105, n80106, n80107, n80108, n80109, n80110, n80111,
    n80112, n80113, n80114, n80115, n80116, n80117, n80118, n80119, n80120,
    n80121, n80122, n80123, n80124, n80125, n80126, n80127, n80128, n80129,
    n80130, n80131, n80132, n80133, n80134, n80135, n80136, n80137, n80138,
    n80139, n80140, n80141, n80142, n80143, n80144, n80145, n80146, n80147,
    n80148, n80149, n80150, n80151, n80152, n80153, n80154, n80155, n80156,
    n80157, n80158, n80159, n80160, n80161, n80162, n80163, n80164, n80165,
    n80166, n80167, n80168, n80169, n80170, n80171, n80172, n80173, n80174,
    n80175, n80176, n80177, n80178, n80179, n80180, n80181, n80182, n80183,
    n80184, n80185, n80186, n80187, n80188, n80189, n80190, n80191, n80192,
    n80193, n80194, n80195, n80196, n80197, n80198, n80199, n80200, n80201,
    n80202, n80203, n80204, n80205, n80206, n80207, n80208, n80209, n80210,
    n80211, n80212, n80213, n80214, n80215, n80216, n80217, n80218, n80219,
    n80220, n80221, n80222, n80223, n80224, n80225, n80226, n80227, n80228,
    n80229, n80230, n80231, n80232, n80233, n80234, n80235, n80236, n80237,
    n80238, n80239, n80240, n80241, n80242, n80243, n80244, n80245, n80246,
    n80247, n80248, n80249, n80250, n80251, n80252, n80253, n80254, n80255,
    n80256, n80257, n80258, n80259, n80260, n80261, n80262, n80263, n80264,
    n80265, n80266, n80267, n80268, n80269, n80270, n80271, n80272, n80273,
    n80274, n80275, n80276, n80277, n80278, n80279, n80280, n80281, n80282,
    n80283, n80284, n80285, n80286, n80287, n80288, n80289, n80290, n80291,
    n80292, n80293, n80294, n80295, n80296, n80297, n80298, n80299, n80300,
    n80301, n80302, n80303, n80304, n80305, n80306, n80307, n80308, n80309,
    n80310, n80311, n80312, n80313, n80314, n80315, n80316, n80317, n80318,
    n80319, n80320, n80321, n80322, n80323, n80324, n80325, n80326, n80327,
    n80328, n80329, n80330, n80331, n80332, n80333, n80334, n80335, n80336,
    n80337, n80338, n80339, n80340, n80341, n80342, n80343, n80344, n80345,
    n80346, n80347, n80348, n80349, n80350, n80351, n80352, n80353, n80354,
    n80355, n80356, n80357, n80358, n80359, n80360, n80361, n80362, n80363,
    n80364, n80365, n80366, n80367, n80368, n80369, n80370, n80371, n80372,
    n80373, n80374, n80375, n80376, n80377, n80378, n80379, n80380, n80381,
    n80382, n80383, n80384, n80385, n80386, n80387, n80388, n80389, n80390,
    n80391, n80392, n80393, n80394, n80395, n80396, n80397, n80398, n80399,
    n80400, n80401, n80402, n80403, n80404, n80405, n80406, n80407, n80408,
    n80409, n80410, n80411, n80412, n80413, n80414, n80415, n80416, n80417,
    n80418, n80419, n80420, n80421, n80422, n80423, n80424, n80425, n80426,
    n80427, n80428, n80429, n80430, n80431, n80432, n80433, n80434, n80435,
    n80436, n80437, n80438, n80439, n80440, n80441, n80442, n80443, n80444,
    n80445, n80446, n80447, n80448, n80449, n80450, n80451, n80452, n80453,
    n80454, n80455, n80456, n80457, n80458, n80459, n80460, n80461, n80462,
    n80463, n80464, n80465, n80466, n80467, n80468, n80469, n80470, n80471,
    n80472, n80473, n80474, n80475, n80476, n80477, n80478, n80479, n80480,
    n80481, n80482, n80483, n80484, n80485, n80486, n80487, n80488, n80489,
    n80490, n80491, n80492, n80493, n80494, n80495, n80496, n80497, n80498,
    n80499, n80500, n80501, n80502, n80503, n80504, n80505, n80506, n80507,
    n80508, n80509, n80510, n80511, n80512, n80513, n80514, n80515, n80516,
    n80517, n80518, n80519, n80520, n80521, n80522, n80523, n80524, n80525,
    n80526, n80527, n80528, n80529, n80530, n80531, n80532, n80533, n80534,
    n80535, n80536, n80537, n80538, n80539, n80540, n80541, n80542, n80543,
    n80544, n80545, n80546, n80547, n80548, n80549, n80550, n80551, n80552,
    n80553, n80554, n80555, n80556, n80557, n80558, n80559, n80560, n80561,
    n80562, n80563, n80564, n80565, n80566, n80567, n80568, n80569, n80570,
    n80571, n80572, n80573, n80574, n80575, n80576, n80577, n80578, n80579,
    n80580, n80581, n80582, n80583, n80584, n80585, n80586, n80587, n80588,
    n80589, n80590, n80591, n80592, n80593, n80594, n80595, n80596, n80597,
    n80598, n80599, n80600, n80601, n80602, n80603, n80604, n80605, n80606,
    n80607, n80608, n80609, n80610, n80611, n80612, n80613, n80614, n80615,
    n80616, n80617, n80618, n80619, n80620, n80621, n80622, n80623, n80624,
    n80625, n80626, n80627, n80628, n80629, n80630, n80631, n80632, n80633,
    n80634, n80635, n80636, n80637, n80638, n80639, n80640, n80641, n80642,
    n80643, n80644, n80645, n80646, n80647, n80648, n80649, n80650, n80651,
    n80652, n80653, n80654, n80655, n80656, n80657, n80658, n80659, n80660,
    n80661, n80662, n80663, n80664, n80665, n80666, n80667, n80668, n80669,
    n80670, n80671, n80672, n80673, n80674, n80675, n80676, n80677, n80678,
    n80679, n80680, n80681, n80682, n80683, n80684, n80685, n80686, n80687,
    n80688, n80689, n80690, n80691, n80692, n80693, n80694, n80695, n80696,
    n80697, n80698, n80699, n80700, n80701, n80702, n80703, n80704, n80705,
    n80706, n80707, n80708, n80709, n80710, n80711, n80712, n80713, n80714,
    n80715, n80716, n80717, n80718, n80719, n80720, n80721, n80722, n80723,
    n80724, n80725, n80726, n80727, n80728, n80729, n80730, n80731, n80732,
    n80733, n80734, n80735, n80736, n80737, n80738, n80739, n80740, n80741,
    n80742, n80743, n80744, n80745, n80746, n80747, n80748, n80749, n80750,
    n80751, n80752, n80753, n80754, n80755, n80756, n80757, n80758, n80759,
    n80760, n80761, n80762, n80763, n80764, n80765, n80766, n80767, n80768,
    n80769, n80770, n80771, n80772, n80773, n80774, n80775, n80776, n80777,
    n80778, n80779, n80780, n80781, n80782, n80783, n80784, n80785, n80786,
    n80787, n80788, n80789, n80790, n80791, n80792, n80793, n80794, n80795,
    n80796, n80797, n80798, n80799, n80800, n80801, n80802, n80803, n80804,
    n80805, n80806, n80807, n80808, n80809, n80810, n80811, n80812, n80813,
    n80814, n80815, n80816, n80817, n80818, n80819, n80820, n80821, n80822,
    n80823, n80824, n80825, n80826, n80827, n80828, n80829, n80830, n80831,
    n80832, n80833, n80834, n80835, n80836, n80837, n80838, n80839, n80840,
    n80841, n80842, n80843, n80844, n80845, n80846, n80847, n80848, n80849,
    n80850, n80851, n80852, n80853, n80854, n80855, n80856, n80857, n80858,
    n80859, n80860, n80861, n80862, n80863, n80864, n80865, n80866, n80867,
    n80868, n80869, n80870, n80871, n80872, n80873, n80874, n80875, n80876,
    n80877, n80878, n80879, n80880, n80881, n80882, n80883, n80884, n80885,
    n80886, n80887, n80888, n80889, n80890, n80891, n80892, n80893, n80894,
    n80895, n80896, n80897, n80898, n80899, n80900, n80901, n80902, n80903,
    n80904, n80905, n80906, n80907, n80908, n80909, n80910, n80911, n80912,
    n80913, n80914, n80915, n80916, n80917, n80918, n80919, n80920, n80921,
    n80922, n80923, n80924, n80925, n80926, n80927, n80928, n80929, n80930,
    n80931, n80932, n80933, n80934, n80935, n80936, n80937, n80938, n80939,
    n80940, n80941, n80942, n80943, n80944, n80945, n80946, n80947, n80948,
    n80949, n80950, n80951, n80952, n80953, n80954, n80955, n80956, n80957,
    n80958, n80959, n80960, n80961, n80962, n80963, n80964, n80965, n80966,
    n80967, n80968, n80969, n80970, n80971, n80972, n80973, n80974, n80975,
    n80976, n80977, n80978, n80979, n80980, n80981, n80982, n80983, n80984,
    n80985, n80986, n80987, n80988, n80989, n80990, n80991, n80992, n80993,
    n80994, n80995, n80996, n80997, n80998, n80999, n81000, n81001, n81002,
    n81003, n81004, n81005, n81006, n81007, n81008, n81009, n81010, n81011,
    n81012, n81013, n81014, n81015, n81016, n81017, n81018, n81019, n81020,
    n81021, n81022, n81023, n81024, n81025, n81026, n81027, n81028, n81029,
    n81030, n81031, n81032, n81033, n81034, n81035, n81036, n81037, n81038,
    n81039, n81040, n81041, n81042, n81043, n81044, n81045, n81046, n81047,
    n81048, n81049, n81050, n81051, n81052, n81053, n81054, n81055, n81056,
    n81057, n81058, n81059, n81060, n81061, n81062, n81063, n81064, n81065,
    n81066, n81067, n81068, n81069, n81070, n81071, n81072, n81073, n81074,
    n81075, n81076, n81077, n81078, n81079, n81080, n81081, n81082, n81083,
    n81084, n81085, n81086, n81087, n81088, n81089, n81090, n81091, n81092,
    n81093, n81094, n81095, n81096, n81097, n81098, n81099, n81100, n81101,
    n81102, n81103, n81104, n81105, n81106, n81107, n81108, n81109, n81110,
    n81111, n81112, n81113, n81114, n81115, n81116, n81117, n81118, n81119,
    n81120, n81121, n81122, n81123, n81124, n81125, n81126, n81127, n81128,
    n81129, n81130, n81131, n81132, n81133, n81134, n81135, n81136, n81137,
    n81138, n81139, n81140, n81141, n81142, n81143, n81144, n81145, n81146,
    n81147, n81148, n81149, n81150, n81151, n81152, n81153, n81154, n81155,
    n81156, n81157, n81158, n81159, n81160, n81161, n81162, n81163, n81164,
    n81165, n81166, n81167, n81168, n81169, n81170, n81171, n81172, n81173,
    n81174, n81175, n81176, n81177, n81178, n81179, n81180, n81181, n81182,
    n81183, n81184, n81185, n81186, n81187, n81188, n81189, n81190, n81191,
    n81192, n81193, n81194, n81195, n81196, n81197, n81198, n81199, n81200,
    n81201, n81202, n81203, n81204, n81205, n81206, n81207, n81208, n81209,
    n81210, n81211, n81212, n81213, n81214, n81215, n81216, n81217, n81218,
    n81219, n81220, n81221, n81222, n81223, n81224, n81225, n81226, n81227,
    n81228, n81229, n81230, n81231, n81232, n81233, n81234, n81235, n81236,
    n81237, n81238, n81239, n81240, n81241, n81242, n81243, n81244, n81245,
    n81246, n81247, n81248, n81249, n81250, n81251, n81252, n81253, n81254,
    n81255, n81256, n81257, n81258, n81259, n81260, n81261, n81262, n81263,
    n81264, n81265, n81266, n81267, n81268, n81269, n81270, n81271, n81272,
    n81273, n81274, n81275, n81276, n81277, n81278, n81279, n81280, n81281,
    n81282, n81283, n81284, n81285, n81286, n81287, n81288, n81289, n81290,
    n81291, n81292, n81293, n81294, n81295, n81296, n81297, n81298, n81299,
    n81300, n81301, n81302, n81303, n81304, n81305, n81306, n81307, n81308,
    n81309, n81310, n81311, n81312, n81313, n81314, n81315, n81316, n81317,
    n81318, n81319, n81320, n81321, n81322, n81323, n81324, n81325, n81326,
    n81327, n81328, n81329, n81330, n81331, n81332, n81333, n81334, n81335,
    n81336, n81337, n81338, n81339, n81340, n81341, n81342, n81343, n81344,
    n81345, n81346, n81347, n81348, n81349, n81350, n81351, n81352, n81353,
    n81354, n81355, n81356, n81357, n81358, n81359, n81360, n81361, n81362,
    n81363, n81364, n81365, n81366, n81367, n81368, n81369, n81370, n81371,
    n81372, n81373, n81374, n81375, n81376, n81377, n81378, n81379, n81380,
    n81381, n81382, n81383, n81384, n81385, n81386, n81387, n81388, n81389,
    n81390, n81391, n81392, n81393, n81394, n81395, n81396, n81397, n81398,
    n81399, n81400, n81401, n81402, n81403, n81404, n81405, n81406, n81407,
    n81408, n81409, n81410, n81411, n81412, n81413, n81414, n81415, n81416,
    n81417, n81418, n81419, n81420, n81421, n81422, n81423, n81424, n81425,
    n81426, n81427, n81428, n81429, n81430, n81431, n81432, n81433, n81434,
    n81435, n81436, n81437, n81438, n81439, n81440, n81441, n81442, n81443,
    n81444, n81445, n81446, n81447, n81448, n81449, n81450, n81451, n81452,
    n81453, n81454, n81455, n81456, n81457, n81458, n81459, n81460, n81461,
    n81462, n81463, n81464, n81465, n81466, n81467, n81468, n81469, n81470,
    n81471, n81472, n81473, n81474, n81475, n81476, n81477, n81478, n81479,
    n81480, n81481, n81482, n81483, n81484, n81485, n81486, n81487, n81488,
    n81489, n81490, n81491, n81492, n81493, n81494, n81495, n81496, n81497,
    n81498, n81499, n81500, n81501, n81502, n81503, n81504, n81505, n81506,
    n81507, n81508, n81509, n81510, n81511, n81512, n81513, n81514, n81515,
    n81516, n81517, n81518, n81519, n81520, n81521, n81522, n81523, n81524,
    n81525, n81526, n81527, n81528, n81529, n81530, n81531, n81532, n81533,
    n81534, n81535, n81536, n81537, n81538, n81539, n81540, n81541, n81542,
    n81543, n81544, n81545, n81546, n81547, n81548, n81549, n81550, n81551,
    n81552, n81553, n81554, n81555, n81556, n81557, n81558, n81559, n81560,
    n81561, n81562, n81563, n81564, n81565, n81566, n81567, n81568, n81569,
    n81570, n81571, n81572, n81573, n81574, n81575, n81576, n81577, n81578,
    n81579, n81580, n81581, n81582, n81583, n81584, n81585, n81586, n81587,
    n81588, n81589, n81590, n81591, n81592, n81593, n81594, n81595, n81596,
    n81597, n81598, n81599, n81600, n81601, n81602, n81603, n81604, n81605,
    n81606, n81607, n81608, n81609, n81610, n81611, n81612, n81613, n81614,
    n81615, n81616, n81617, n81618, n81619, n81620, n81621, n81622, n81623,
    n81624, n81625, n81626, n81627, n81628, n81629, n81630, n81631, n81632,
    n81633, n81634, n81635, n81636, n81637, n81638, n81639, n81640, n81641,
    n81642, n81643, n81644, n81645, n81646, n81647, n81648, n81649, n81650,
    n81651, n81652, n81653, n81654, n81655, n81656, n81657, n81658, n81659,
    n81660, n81661, n81662, n81663, n81664, n81665, n81666, n81667, n81668,
    n81669, n81670, n81671, n81672, n81673, n81674, n81675, n81676, n81677,
    n81678, n81679, n81680, n81681, n81682, n81683, n81684, n81685, n81686,
    n81687, n81688, n81689, n81690, n81691, n81692, n81693, n81694, n81695,
    n81696, n81697, n81698, n81699, n81700, n81701, n81702, n81703, n81704,
    n81705, n81706, n81707, n81708, n81709, n81710, n81711, n81712, n81713,
    n81714, n81715, n81716, n81717, n81718, n81719, n81720, n81721, n81722,
    n81723, n81724, n81725, n81726, n81727, n81728, n81729, n81730, n81731,
    n81732, n81733, n81734, n81735, n81736, n81737, n81738, n81739, n81740,
    n81741, n81742, n81743, n81744, n81745, n81746, n81747, n81748, n81749,
    n81750, n81751, n81752, n81753, n81754, n81755, n81756, n81757, n81758,
    n81759, n81760, n81761, n81762, n81763, n81764, n81765, n81766, n81767,
    n81768, n81769, n81770, n81771, n81772, n81773, n81774, n81775, n81776,
    n81777, n81778, n81779, n81780, n81781, n81782, n81783, n81784, n81785,
    n81786, n81787, n81788, n81789, n81790, n81791, n81792, n81793, n81794,
    n81795, n81796, n81797, n81798, n81799, n81800, n81801, n81802, n81803,
    n81804, n81805, n81806, n81807, n81808, n81809, n81810, n81811, n81812,
    n81813, n81814, n81815, n81816, n81817, n81818, n81819, n81820, n81821,
    n81822, n81823, n81824, n81825, n81826, n81827, n81828, n81829, n81830,
    n81831, n81832, n81833, n81834, n81835, n81836, n81837, n81838, n81839,
    n81840, n81841, n81842, n81843, n81844, n81845, n81846, n81847, n81848,
    n81849, n81850, n81851, n81852, n81853, n81854, n81855, n81856, n81857,
    n81858, n81859, n81860, n81861, n81862, n81863, n81864, n81865, n81866,
    n81867, n81868, n81869, n81870, n81871, n81872, n81873, n81874, n81875,
    n81876, n81877, n81878, n81879, n81880, n81881, n81882, n81883, n81884,
    n81885, n81886, n81887, n81888, n81889, n81890, n81891, n81892, n81893,
    n81894, n81895, n81896, n81897, n81898, n81899, n81900, n81901, n81902,
    n81903, n81904, n81905, n81906, n81907, n81908, n81909, n81910, n81911,
    n81912, n81913, n81914, n81915, n81916, n81917, n81918, n81919, n81920,
    n81921, n81922, n81923, n81924, n81925, n81926, n81927, n81928, n81929,
    n81930, n81931, n81932, n81933, n81934, n81935, n81936, n81937, n81938,
    n81939, n81940, n81941, n81942, n81943, n81944, n81945, n81946, n81947,
    n81948, n81949, n81950, n81951, n81952, n81953, n81954, n81955, n81956,
    n81957, n81958, n81959, n81960, n81961, n81962, n81963, n81964, n81965,
    n81966, n81967, n81968, n81969, n81970, n81971, n81972, n81973, n81974,
    n81975, n81976, n81977, n81978, n81979, n81980, n81981, n81982, n81983,
    n81984, n81985, n81986, n81987, n81988, n81989, n81990, n81991, n81992,
    n81993, n81994, n81995, n81996, n81997, n81998, n81999, n82000, n82001,
    n82002, n82003, n82004, n82005, n82006, n82007, n82008, n82009, n82010,
    n82011, n82012, n82013, n82014, n82015, n82016, n82017, n82018, n82019,
    n82020, n82021, n82022, n82023, n82024, n82025, n82026, n82027, n82028,
    n82029, n82030, n82031, n82032, n82033, n82034, n82035, n82036, n82037,
    n82038, n82039, n82040, n82041, n82042, n82043, n82044, n82045, n82046,
    n82047, n82048, n82049, n82050, n82051, n82052, n82053, n82054, n82055,
    n82056, n82057, n82058, n82059, n82060, n82061, n82062, n82063, n82064,
    n82065, n82066, n82067, n82068, n82069, n82070, n82071, n82072, n82073,
    n82074, n82075, n82076, n82077, n82078, n82079, n82080, n82081, n82082,
    n82083, n82084, n82085, n82086, n82087, n82088, n82089, n82090, n82091,
    n82092, n82093, n82094, n82095, n82096, n82097, n82098, n82099, n82100,
    n82101, n82102, n82103, n82104, n82105, n82106, n82107, n82108, n82109,
    n82110, n82111, n82112, n82113, n82114, n82115, n82116, n82117, n82118,
    n82119, n82120, n82121, n82122, n82123, n82124, n82125, n82126, n82127,
    n82128, n82129, n82130, n82131, n82132, n82133, n82134, n82135, n82136,
    n82137, n82138, n82139, n82140, n82141, n82142, n82143, n82144, n82145,
    n82146, n82147, n82148, n82149, n82150, n82151, n82152, n82153, n82154,
    n82155, n82156, n82157, n82158, n82159, n82160, n82161, n82162, n82163,
    n82164, n82165, n82166, n82167, n82168, n82169, n82170, n82171, n82172,
    n82173, n82174, n82175, n82176, n82177, n82178, n82179, n82180, n82181,
    n82182, n82183, n82184, n82185, n82186, n82187, n82188, n82189, n82190,
    n82191, n82192, n82193, n82194, n82195, n82196, n82197, n82198, n82199,
    n82200, n82201, n82202, n82203, n82204, n82205, n82206, n82207, n82208,
    n82209, n82210, n82211, n82212, n82213, n82214, n82215, n82216, n82217,
    n82218, n82219, n82220, n82221, n82222, n82223, n82224, n82225, n82226,
    n82227, n82228, n82229, n82230, n82231, n82232, n82233, n82234, n82235,
    n82236, n82237, n82238, n82239, n82240, n82241, n82242, n82243, n82244,
    n82245, n82246, n82247, n82248, n82249, n82250, n82251, n82252, n82253,
    n82254, n82255, n82256, n82257, n82258, n82259, n82260, n82261, n82262,
    n82263, n82264, n82265, n82266, n82267, n82268, n82269, n82270, n82271,
    n82272, n82273, n82274, n82275, n82276, n82277, n82278, n82279, n82280,
    n82281, n82282, n82283, n82284, n82285, n82286, n82287, n82288, n82289,
    n82290, n82291, n82292, n82293, n82294, n82295, n82296, n82297, n82298,
    n82299, n82300, n82301, n82302, n82303, n82304, n82305, n82306, n82307,
    n82308, n82309, n82310, n82311, n82312, n82313, n82314, n82315, n82316,
    n82317, n82318, n82319, n82320, n82321, n82322, n82323, n82324, n82325,
    n82326, n82327, n82328, n82329, n82330, n82331, n82332, n82333, n82334,
    n82335, n82336, n82337, n82338, n82339, n82340, n82341, n82342, n82343,
    n82344, n82345, n82346, n82347, n82348, n82349, n82350, n82351, n82352,
    n82353, n82354, n82355, n82356, n82357, n82358, n82359, n82360, n82361,
    n82362, n82363, n82364, n82365, n82366, n82367, n82368, n82369, n82370,
    n82371, n82372, n82373, n82374, n82375, n82376, n82377, n82378, n82379,
    n82380, n82381, n82382, n82383, n82384, n82385, n82386, n82387, n82388,
    n82389, n82390, n82391, n82392, n82393, n82394, n82395, n82396, n82397,
    n82398, n82399, n82400, n82401, n82402, n82403, n82404, n82405, n82406,
    n82407, n82408, n82409, n82410, n82411, n82412, n82413, n82414, n82415,
    n82416, n82417, n82418, n82419, n82420, n82421, n82422, n82423, n82424,
    n82425, n82426, n82427, n82428, n82429, n82430, n82431, n82432, n82433,
    n82434, n82435, n82436, n82437, n82438, n82439, n82440, n82441, n82442,
    n82443, n82444, n82445, n82446, n82447, n82448, n82449, n82450, n82451,
    n82452, n82453, n82454, n82455, n82456, n82457, n82458, n82459, n82460,
    n82461, n82462, n82463, n82464, n82465, n82466, n82467, n82468, n82469,
    n82470, n82471, n82472, n82473, n82474, n82475, n82476, n82477, n82478,
    n82479, n82480, n82481, n82482, n82483, n82484, n82485, n82486, n82487,
    n82488, n82489, n82490, n82491, n82492, n82493, n82494, n82495, n82496,
    n82497, n82498, n82499, n82500, n82501, n82502, n82503, n82504, n82505,
    n82506, n82507, n82508, n82509, n82510, n82511, n82512, n82513, n82514,
    n82515, n82516, n82517, n82518, n82519, n82520, n82521, n82522, n82523,
    n82524, n82525, n82526, n82527, n82528, n82529, n82530, n82531, n82532,
    n82533, n82534, n82535, n82536, n82537, n82538, n82539, n82540, n82541,
    n82542, n82543, n82544, n82545, n82546, n82547, n82548, n82549, n82550,
    n82551, n82552, n82553, n82554, n82555, n82556, n82557, n82558, n82559,
    n82560, n82561, n82562, n82563, n82564, n82565, n82566, n82567, n82568,
    n82569, n82570, n82571, n82572, n82573, n82574, n82575, n82576, n82577,
    n82578, n82579, n82580, n82581, n82582, n82583, n82584, n82585, n82586,
    n82587, n82588, n82589, n82590, n82591, n82592, n82593, n82594, n82595,
    n82596, n82597, n82598, n82599, n82600, n82601, n82602, n82603, n82604,
    n82605, n82606, n82607, n82608, n82609, n82610, n82611, n82612, n82613,
    n82614, n82615, n82616, n82617, n82618, n82619, n82620, n82621, n82622,
    n82623, n82624, n82625, n82626, n82627, n82628, n82629, n82630, n82631,
    n82632, n82633, n82634, n82635, n82636, n82637, n82638, n82639, n82640,
    n82641, n82642, n82643, n82644, n82645, n82646, n82647, n82648, n82649,
    n82650, n82651, n82652, n82653, n82654, n82655, n82656, n82657, n82658,
    n82659, n82660, n82661, n82662, n82663, n82664, n82665, n82666, n82667,
    n82668, n82669, n82670, n82671, n82672, n82673, n82674, n82675, n82676,
    n82677, n82678, n82679, n82680, n82681, n82682, n82683, n82684, n82685,
    n82686, n82687, n82688, n82689, n82690, n82691, n82692, n82693, n82694,
    n82695, n82696, n82697, n82698, n82699, n82700, n82701, n82702, n82703,
    n82704, n82705, n82706, n82707, n82708, n82709, n82710, n82711, n82712,
    n82713, n82714, n82715, n82716, n82717, n82718, n82719, n82720, n82721,
    n82722, n82723, n82724, n82725, n82726, n82727, n82728, n82729, n82730,
    n82731, n82732, n82733, n82734, n82735, n82736, n82737, n82738, n82739,
    n82740, n82741, n82742, n82743, n82744, n82745, n82746, n82747, n82748,
    n82749, n82750, n82751, n82752, n82753, n82754, n82755, n82756, n82757,
    n82758, n82759, n82760, n82761, n82762, n82763, n82764, n82765, n82766,
    n82767, n82768, n82769, n82770, n82771, n82772, n82773, n82774, n82775,
    n82776, n82777, n82778, n82779, n82780, n82781, n82782, n82783, n82784,
    n82785, n82786, n82787, n82788, n82789, n82790, n82791, n82792, n82793,
    n82794, n82795, n82796, n82797, n82798, n82799, n82800, n82801, n82802,
    n82803, n82804, n82805, n82806, n82807, n82808, n82809, n82810, n82811,
    n82812, n82813, n82814, n82815, n82816, n82817, n82818, n82819, n82820,
    n82821, n82822, n82823, n82824, n82825, n82826, n82827, n82828, n82829,
    n82830, n82831, n82832, n82833, n82834, n82835, n82836, n82837, n82838,
    n82839, n82840, n82841, n82842, n82843, n82844, n82845, n82846, n82847,
    n82848, n82849, n82850, n82851, n82852, n82853, n82854, n82855, n82856,
    n82857, n82858, n82859, n82860, n82861, n82862, n82863, n82864, n82865,
    n82866, n82867, n82868, n82869, n82870, n82871, n82872, n82873, n82874,
    n82875, n82876, n82877, n82878, n82879, n82880, n82881, n82882, n82883,
    n82884, n82885, n82886, n82887, n82888, n82889, n82890, n82891, n82892,
    n82893, n82894, n82895, n82896, n82897, n82898, n82899, n82900, n82901,
    n82902, n82903, n82904, n82905, n82906, n82907, n82908, n82909, n82910,
    n82911, n82912, n82913, n82914, n82915, n82916, n82917, n82918, n82919,
    n82920, n82921, n82922, n82923, n82924, n82925, n82926, n82927, n82928,
    n82929, n82930, n82931, n82932, n82933, n82934, n82935, n82936, n82937,
    n82938, n82939, n82940, n82941, n82942, n82943, n82944, n82945, n82946,
    n82947, n82948, n82949, n82950, n82951, n82952, n82953, n82954, n82955,
    n82956, n82957, n82958, n82959, n82960, n82961, n82962, n82963, n82964,
    n82965, n82966, n82967, n82968, n82969, n82970, n82971, n82972, n82973,
    n82974, n82975, n82976, n82977, n82978, n82979, n82980, n82981, n82982,
    n82983, n82984, n82985, n82986, n82987, n82988, n82989, n82990, n82991,
    n82992, n82993, n82994, n82995, n82996, n82997, n82998, n82999, n83000,
    n83001, n83002, n83003, n83004, n83005, n83006, n83007, n83008, n83009,
    n83010, n83011, n83012, n83013, n83014, n83015, n83016, n83017, n83018,
    n83019, n83020, n83021, n83022, n83023, n83024, n83025, n83026, n83027,
    n83028, n83029, n83030, n83031, n83032, n83033, n83034, n83035, n83036,
    n83037, n83038, n83039, n83040, n83041, n83042, n83043, n83044, n83045,
    n83046, n83047, n83048, n83049, n83050, n83051, n83052, n83053, n83054,
    n83055, n83056, n83057, n83058, n83059, n83060, n83061, n83062, n83063,
    n83064, n83065, n83066, n83067, n83068, n83069, n83070, n83071, n83072,
    n83073, n83074, n83075, n83076, n83077, n83078, n83079, n83080, n83081,
    n83082, n83083, n83084, n83085, n83086, n83087, n83088, n83089, n83090,
    n83091, n83092, n83093, n83094, n83095, n83096, n83097, n83098, n83099,
    n83100, n83101, n83102, n83103, n83104, n83105, n83106, n83107, n83108,
    n83109, n83110, n83111, n83112, n83113, n83114, n83115, n83116, n83117,
    n83118, n83119, n83120, n83121, n83122, n83123, n83124, n83125, n83126,
    n83127, n83128, n83129, n83130, n83131, n83132, n83133, n83134, n83135,
    n83136, n83137, n83138, n83139, n83140, n83141, n83142, n83143, n83144,
    n83145, n83146, n83147, n83148, n83149, n83150, n83151, n83152, n83153,
    n83154, n83155, n83156, n83157, n83158, n83159, n83160, n83161, n83162,
    n83163, n83164, n83165, n83166, n83167, n83168, n83169, n83170, n83171,
    n83172, n83173, n83174, n83175, n83176, n83177, n83178, n83179, n83180,
    n83181, n83182, n83183, n83184, n83185, n83186, n83187, n83188, n83189,
    n83190, n83191, n83192, n83193, n83194, n83195, n83196, n83197, n83198,
    n83199, n83200, n83201, n83202, n83203, n83204, n83205, n83206, n83207,
    n83208, n83209, n83210, n83211, n83212, n83213, n83214, n83215, n83216,
    n83217, n83218, n83219, n83220, n83221, n83222, n83223, n83224, n83225,
    n83226, n83227, n83228, n83229, n83230, n83231, n83232, n83233, n83234,
    n83235, n83236, n83237, n83238, n83239, n83240, n83241, n83242, n83243,
    n83244, n83245, n83246, n83247, n83248, n83249, n83250, n83251, n83252,
    n83253, n83254, n83255, n83256, n83257, n83258, n83259, n83260, n83261,
    n83262, n83263, n83264, n83265, n83266, n83267, n83268, n83269, n83270,
    n83271, n83272, n83273, n83274, n83275, n83276, n83277, n83278, n83279,
    n83280, n83281, n83282, n83283, n83284, n83285, n83286, n83287, n83288,
    n83289, n83290, n83291, n83292, n83293, n83294, n83295, n83296, n83297,
    n83298, n83299, n83300, n83301, n83302, n83303, n83304, n83305, n83306,
    n83307, n83308, n83309, n83310, n83311, n83312, n83313, n83314, n83315,
    n83316, n83317, n83318, n83319, n83320, n83321, n83322, n83323, n83324,
    n83325, n83326, n83327, n83328, n83329, n83330, n83331, n83332, n83333,
    n83334, n83335, n83336, n83337, n83338, n83339, n83340, n83341, n83342,
    n83343, n83344, n83345, n83346, n83347, n83348, n83349, n83350, n83351,
    n83352, n83353, n83354, n83355, n83356, n83357, n83358, n83359, n83360,
    n83361, n83362, n83363, n83364, n83365, n83366, n83367, n83368, n83369,
    n83370, n83371, n83372, n83373, n83374, n83375, n83376, n83377, n83378,
    n83379, n83380, n83381, n83382, n83383, n83384, n83385, n83386, n83387,
    n83388, n83389, n83390, n83391, n83392, n83393, n83394, n83395, n83396,
    n83397, n83398, n83399, n83400, n83401, n83402, n83403, n83404, n83405,
    n83406, n83407, n83408, n83409, n83410, n83411, n83412, n83413, n83414,
    n83415, n83416, n83417, n83418, n83419, n83420, n83421, n83422, n83423,
    n83424, n83425, n83426, n83427, n83428, n83429, n83430, n83431, n83432,
    n83433, n83434, n83435, n83436, n83437, n83438, n83439, n83440, n83441,
    n83442, n83443, n83444, n83445, n83446, n83447, n83448, n83449, n83450,
    n83451, n83452, n83453, n83454, n83455, n83456, n83457, n83458, n83459,
    n83460, n83461, n83462, n83463, n83464, n83465, n83466, n83467, n83468,
    n83469, n83470, n83471, n83472, n83473, n83474, n83475, n83476, n83477,
    n83478, n83479, n83480, n83481, n83482, n83483, n83484, n83485, n83486,
    n83487, n83488, n83489, n83490, n83491, n83492, n83493, n83494, n83495,
    n83496, n83497, n83498, n83499, n83500, n83501, n83502, n83503, n83504,
    n83505, n83506, n83507, n83508, n83509, n83510, n83511, n83512, n83513,
    n83514, n83515, n83516, n83517, n83518, n83519, n83520, n83521, n83523,
    n83524, n83525, n83526, n83527, n83528, n83529, n83530, n83531, n83532,
    n83533, n83534, n83535, n83536, n83537, n83538, n83539, n83540, n83541,
    n83542, n83543, n83544, n83545, n83546, n83547, n83548, n83549, n83550,
    n83551, n83552, n83553, n83554, n83555, n83556, n83557, n83558, n83559,
    n83560, n83561, n83562, n83563, n83564, n83565, n83566, n83567, n83568,
    n83569, n83570, n83572, n83573, n83574, n83575, n83576, n83577, n83578,
    n83579, n83580, n83581, n83582, n83583, n83584, n83585, n83586, n83587,
    n83588, n83589, n83590, n83591, n83592, n83593, n83594, n83595, n83596,
    n83597, n83598, n83599, n83600, n83601, n83602, n83603, n83604, n83605,
    n83606, n83607, n83608, n83609, n83610, n83611, n83612, n83614, n83615,
    n83616, n83617, n83618, n83619, n83620, n83621, n83622, n83623, n83624,
    n83625, n83626, n83627, n83628, n83629, n83630, n83631, n83632, n83633,
    n83634, n83635, n83636, n83637, n83638, n83639, n83640, n83641, n83642,
    n83643, n83644, n83645, n83646, n83647, n83648, n83649, n83650, n83651,
    n83652, n83653, n83654, n83655, n83656, n83657, n83658, n83660, n83661,
    n83662, n83663, n83664, n83665, n83666, n83667, n83668, n83669, n83670,
    n83671, n83672, n83673, n83674, n83675, n83676, n83677, n83678, n83679,
    n83680, n83681, n83682, n83683, n83684, n83685, n83686, n83687, n83688,
    n83689, n83690, n83691, n83692, n83693, n83694, n83695, n83696, n83697,
    n83698, n83699, n83701, n83702, n83703, n83704, n83705, n83706, n83707,
    n83708, n83709, n83710, n83711, n83712, n83713, n83714, n83715, n83716,
    n83717, n83718, n83719, n83720, n83721, n83722, n83723, n83724, n83725,
    n83726, n83727, n83728, n83729, n83730, n83731, n83732, n83733, n83734,
    n83735, n83736, n83737, n83738, n83739, n83740, n83741, n83742, n83743,
    n83744, n83745, n83746, n83747, n83749, n83750, n83751, n83752, n83753,
    n83754, n83755, n83756, n83757, n83758, n83759, n83760, n83761, n83762,
    n83763, n83764, n83765, n83766, n83767, n83768, n83769, n83770, n83771,
    n83772, n83773, n83774, n83775, n83776, n83777, n83778, n83779, n83780,
    n83781, n83782, n83783, n83784, n83785, n83787, n83788, n83789, n83790,
    n83791, n83792, n83793, n83794, n83795, n83796, n83797, n83798, n83799,
    n83800, n83801, n83802, n83803, n83804, n83805, n83806, n83807, n83808,
    n83809, n83810, n83811, n83812, n83813, n83814, n83815, n83816, n83817,
    n83818, n83819, n83820, n83821, n83822, n83823, n83824, n83826, n83827,
    n83828, n83829, n83830, n83831, n83832, n83833, n83834, n83835, n83836,
    n83837, n83838, n83839, n83840, n83841, n83842, n83843, n83844, n83845,
    n83846, n83847, n83848, n83849, n83850, n83851, n83853, n83854, n83855,
    n83856, n83857, n83858, n83859, n83860, n83862, n83863, n83864, n83865,
    n83866, n83867, n83868, n83869, n83871, n83872, n83873, n83874, n83875,
    n83876, n83877, n83878, n83880, n83881, n83882, n83883, n83884, n83885,
    n83886, n83887, n83889, n83890, n83891, n83892, n83893, n83894, n83895,
    n83896, n83898, n83899, n83900, n83901, n83902, n83903, n83904, n83905,
    n83907, n83908, n83909, n83910, n83911, n83912, n83913, n83914, n83916,
    n83917, n83918, n83919, n83920, n83921, n83922, n83923, n83924, n83925,
    n83926, n83927, n83928, n83929, n83930, n83931, n83932, n83933, n83934,
    n83935, n83936, n83937, n83938, n83939, n83940, n83942, n83943, n83944,
    n83945, n83946, n83947, n83948, n83949, n83951, n83952, n83953, n83954,
    n83955, n83956, n83957, n83958, n83960, n83961, n83962, n83963, n83964,
    n83965, n83966, n83967, n83969, n83970, n83971, n83972, n83973, n83974,
    n83975, n83976, n83978, n83979, n83980, n83981, n83982, n83983, n83984,
    n83985, n83987, n83988, n83989, n83990, n83991, n83992, n83993, n83994,
    n83996, n83997, n83998, n83999, n84000, n84001, n84002, n84003, n84005,
    n84006, n84007, n84008, n84009, n84010, n84011, n84012, n84013, n84014,
    n84015, n84016, n84017, n84018, n84019, n84020, n84021, n84022, n84023,
    n84024, n84025, n84026, n84027, n84028, n84029, n84031, n84032, n84033,
    n84034, n84035, n84036, n84037, n84038, n84040, n84041, n84042, n84043,
    n84044, n84045, n84046, n84047, n84049, n84050, n84051, n84052, n84053,
    n84054, n84055, n84056, n84058, n84059, n84060, n84061, n84062, n84063,
    n84064, n84065, n84067, n84068, n84069, n84070, n84071, n84072, n84073,
    n84074, n84076, n84077, n84078, n84079, n84080, n84081, n84082, n84083,
    n84085, n84086, n84087, n84088, n84089, n84090, n84091, n84092, n84094,
    n84095, n84096, n84097, n84098, n84099, n84100, n84101, n84102, n84103,
    n84104, n84105, n84106, n84107, n84108, n84109, n84110, n84111, n84112,
    n84113, n84114, n84115, n84116, n84117, n84118, n84119, n84121, n84122,
    n84123, n84124, n84125, n84126, n84127, n84128, n84130, n84131, n84132,
    n84133, n84134, n84135, n84136, n84137, n84139, n84140, n84141, n84142,
    n84143, n84144, n84145, n84146, n84148, n84149, n84150, n84151, n84152,
    n84153, n84154, n84155, n84157, n84158, n84159, n84160, n84161, n84162,
    n84163, n84164, n84166, n84167, n84168, n84169, n84170, n84171, n84172,
    n84173, n84175, n84176, n84177, n84178, n84179, n84180, n84181, n84182,
    n84184, n84185, n84186, n84187, n84188, n84189, n84190, n84191, n84192,
    n84193, n84194, n84195, n84196, n84197, n84198, n84199, n84200, n84201,
    n84202, n84203, n84204, n84205, n84206, n84207, n84209, n84210, n84211,
    n84212, n84213, n84214, n84215, n84216, n84218, n84219, n84220, n84221,
    n84222, n84223, n84224, n84225, n84227, n84228, n84229, n84230, n84231,
    n84232, n84233, n84234, n84236, n84237, n84238, n84239, n84240, n84241,
    n84242, n84243, n84245, n84246, n84247, n84248, n84249, n84250, n84251,
    n84252, n84254, n84255, n84256, n84257, n84258, n84259, n84260, n84261,
    n84263, n84264, n84265, n84266, n84267, n84268, n84269, n84270, n84272,
    n84273, n84274, n84275, n84276, n84277, n84278, n84279, n84280, n84281,
    n84282, n84283, n84284, n84285, n84286, n84287, n84288, n84289, n84290,
    n84291, n84292, n84293, n84294, n84296, n84297, n84298, n84299, n84300,
    n84301, n84302, n84303, n84305, n84306, n84307, n84308, n84309, n84310,
    n84311, n84312, n84314, n84315, n84316, n84317, n84318, n84319, n84320,
    n84321, n84323, n84324, n84325, n84326, n84327, n84328, n84329, n84330,
    n84332, n84333, n84334, n84335, n84336, n84337, n84338, n84339, n84341,
    n84342, n84343, n84344, n84345, n84346, n84347, n84348, n84350, n84351,
    n84352, n84353, n84354, n84355, n84356, n84357, n84359, n84360, n84361,
    n84362, n84363, n84364, n84365, n84366, n84367, n84368, n84369, n84370,
    n84371, n84372, n84373, n84374, n84375, n84376, n84377, n84378, n84379,
    n84380, n84382, n84383, n84384, n84385, n84386, n84387, n84388, n84389,
    n84391, n84392, n84393, n84394, n84395, n84396, n84397, n84398, n84400,
    n84401, n84402, n84403, n84404, n84405, n84406, n84407, n84409, n84410,
    n84411, n84412, n84413, n84414, n84415, n84416, n84418, n84419, n84420,
    n84421, n84422, n84423, n84424, n84425, n84427, n84428, n84429, n84430,
    n84431, n84432, n84433, n84434, n84436, n84437, n84438, n84439, n84440,
    n84441, n84442, n84443, n84445, n84446, n84447, n84448, n84449, n84450,
    n84451, n84452, n84453, n84454, n84455, n84456, n84457, n84458, n84459,
    n84460, n84461, n84462, n84463, n84464, n84465, n84467, n84468, n84469,
    n84470, n84471, n84472, n84473, n84474, n84476, n84477, n84478, n84479,
    n84480, n84481, n84482, n84483, n84485, n84486, n84487, n84488, n84489,
    n84490, n84491, n84492, n84494, n84495, n84496, n84497, n84498, n84499,
    n84500, n84501, n84503, n84504, n84505, n84506, n84507, n84508, n84509,
    n84510, n84512, n84513, n84514, n84515, n84516, n84517, n84518, n84519,
    n84521, n84522, n84523, n84524, n84525, n84526, n84527, n84528, n84530,
    n84531, n84532, n84533, n84534, n84535, n84536, n84537, n84538, n84539,
    n84540, n84541, n84542, n84543, n84544, n84545, n84546, n84547, n84548,
    n84549, n84550, n84551, n84552, n84553, n84555, n84556, n84557, n84558,
    n84559, n84560, n84561, n84562, n84564, n84565, n84566, n84567, n84568,
    n84569, n84570, n84571, n84573, n84574, n84575, n84576, n84577, n84578,
    n84579, n84580, n84582, n84583, n84584, n84585, n84586, n84587, n84588,
    n84589, n84591, n84592, n84593, n84594, n84595, n84596, n84597, n84598,
    n84600, n84601, n84602, n84603, n84604, n84605, n84606, n84607, n84609,
    n84610, n84611, n84612, n84613, n84614, n84615, n84616, n84618, n84619,
    n84620, n84621, n84622, n84623, n84624, n84625, n84626, n84627, n84628,
    n84629, n84630, n84631, n84632, n84633, n84634, n84635, n84636, n84637,
    n84638, n84639, n84640, n84641, n84643, n84644, n84645, n84646, n84647,
    n84648, n84649, n84650, n84652, n84653, n84654, n84655, n84656, n84657,
    n84658, n84659, n84661, n84662, n84663, n84664, n84665, n84666, n84667,
    n84668, n84670, n84671, n84672, n84673, n84674, n84675, n84676, n84677,
    n84679, n84680, n84681, n84682, n84683, n84684, n84685, n84686, n84688,
    n84689, n84690, n84691, n84692, n84693, n84694, n84695, n84697, n84698,
    n84699, n84700, n84701, n84702, n84703, n84704, n84706, n84707, n84708,
    n84709, n84710, n84711, n84712, n84713, n84714, n84715, n84716, n84717,
    n84718, n84719, n84720, n84721, n84722, n84723, n84724, n84725, n84726,
    n84727, n84729, n84730, n84731, n84732, n84733, n84734, n84735, n84736,
    n84738, n84739, n84740, n84741, n84742, n84743, n84744, n84745, n84747,
    n84748, n84749, n84750, n84751, n84752, n84753, n84754, n84756, n84757,
    n84758, n84759, n84760, n84761, n84762, n84763, n84765, n84766, n84767,
    n84768, n84769, n84770, n84771, n84772, n84774, n84775, n84776, n84777,
    n84778, n84779, n84780, n84781, n84783, n84784, n84785, n84786, n84787,
    n84788, n84789, n84790, n84792, n84793, n84794, n84795, n84796, n84797,
    n84798, n84799, n84800, n84801, n84802, n84803, n84804, n84805, n84806,
    n84807, n84808, n84809, n84810, n84811, n84812, n84813, n84814, n84815,
    n84816, n84818, n84819, n84820, n84821, n84822, n84823, n84824, n84825,
    n84827, n84828, n84829, n84830, n84831, n84832, n84833, n84834, n84836,
    n84837, n84838, n84839, n84840, n84841, n84842, n84843, n84845, n84846,
    n84847, n84848, n84849, n84850, n84851, n84852, n84854, n84855, n84856,
    n84857, n84858, n84859, n84860, n84861, n84863, n84864, n84865, n84866,
    n84867, n84868, n84869, n84870, n84872, n84873, n84874, n84875, n84876,
    n84877, n84878, n84879, n84881, n84882, n84883, n84884, n84885, n84886,
    n84887, n84888, n84889, n84890, n84891, n84892, n84893, n84894, n84895,
    n84896, n84897, n84898, n84899, n84900, n84901, n84903, n84904, n84905,
    n84906, n84907, n84908, n84909, n84910, n84912, n84913, n84914, n84915,
    n84916, n84917, n84918, n84919, n84921, n84922, n84923, n84924, n84925,
    n84926, n84927, n84928, n84930, n84931, n84932, n84933, n84934, n84935,
    n84936, n84937, n84939, n84940, n84941, n84942, n84943, n84944, n84945,
    n84946, n84948, n84949, n84950, n84951, n84952, n84953, n84954, n84955,
    n84957, n84958, n84959, n84960, n84961, n84962, n84963, n84964, n84966,
    n84967, n84968, n84969, n84970, n84971, n84972, n84973, n84974, n84975,
    n84976, n84977, n84978, n84979, n84980, n84981, n84982, n84983, n84984,
    n84985, n84986, n84988, n84989, n84990, n84991, n84992, n84993, n84994,
    n84995, n84997, n84998, n84999, n85000, n85001, n85002, n85003, n85004,
    n85006, n85007, n85008, n85009, n85010, n85011, n85012, n85013, n85015,
    n85016, n85017, n85018, n85019, n85020, n85021, n85022, n85024, n85025,
    n85026, n85027, n85028, n85029, n85030, n85031, n85033, n85034, n85035,
    n85036, n85037, n85038, n85039, n85040, n85042, n85043, n85044, n85045,
    n85046, n85047, n85048, n85049, n85051, n85052, n85053, n85054, n85055,
    n85056, n85057, n85058, n85059, n85060, n85061, n85062, n85063, n85064,
    n85065, n85066, n85067, n85068, n85069, n85070, n85072, n85073, n85074,
    n85075, n85076, n85077, n85078, n85079, n85081, n85082, n85083, n85084,
    n85085, n85086, n85087, n85088, n85090, n85091, n85092, n85093, n85094,
    n85095, n85096, n85097, n85099, n85100, n85101, n85102, n85103, n85104,
    n85105, n85106, n85108, n85109, n85110, n85111, n85112, n85113, n85114,
    n85115, n85117, n85118, n85119, n85120, n85121, n85122, n85123, n85124,
    n85126, n85127, n85128, n85129, n85130, n85131, n85132, n85133, n85135,
    n85136, n85137, n85138, n85139, n85140, n85141, n85142, n85143, n85144,
    n85146, n85147, n85148, n85149, n85150, n85151, n85153, n85154, n85155,
    n85156, n85157, n85158, n85159, n85160, n85162, n85163, n85164, n85165,
    n85166, n85167, n85168, n85170, n85171, n85172, n85173, n85174, n85175,
    n85176, n85178, n85179, n85180, n85181, n85183, n85184, n85185, n85186,
    n85187, n85188, n85189, n85190, n85191, n85192, n85193, n85194, n85195,
    n85197, n85198, n85199, n85200, n85201, n85202, n85203, n85204, n85205,
    n85206, n85207, n85208, n85209, n85211, n85212, n85213, n85214, n85215,
    n85216, n85217, n85218, n85219, n85220, n85221, n85222, n85224, n85225,
    n85226, n85227, n85228, n85230, n85231, n85232, n85233, n85234, n85235,
    n85236, n85237, n85238, n85239, n85240, n85241, n85242, n85243, n85244,
    n85245, n85246, n85247, n85248, n85249, n85250, n85251, n85252, n85253,
    n85254, n85255, n85256, n85257, n85258, n85259, n85260, n85261, n85262,
    n85263, n85264, n85265, n85266, n85267, n85268, n85269, n85270, n85271,
    n85272, n85273, n85274, n85275, n85276, n85277, n85278, n85279, n85280,
    n85281, n85282, n85283, n85284, n85285, n85286, n85287, n85288, n85289,
    n85290, n85291, n85292, n85293, n85294, n85295, n85296, n85297, n85298,
    n85299, n85300, n85301, n85302, n85303, n85304, n85305, n85306, n85307,
    n85308, n85309, n85310, n85311, n85312, n85313, n85314, n85315, n85316,
    n85317, n85318, n85319, n85320, n85321, n85322, n85323, n85324, n85325,
    n85326, n85327, n85328, n85329, n85330, n85331, n85332, n85333, n85334,
    n85335, n85336, n85337, n85338, n85339, n85340, n85341, n85342, n85343,
    n85344, n85345, n85346, n85347, n85348, n85349, n85350, n85351, n85352,
    n85353, n85354, n85355, n85356, n85357, n85358, n85359, n85360, n85361,
    n85362, n85363, n85364, n85365, n85366, n85367, n85368, n85369, n85370,
    n85371, n85372, n85373, n85374, n85375, n85376, n85377, n85378, n85379,
    n85380, n85381, n85382, n85383, n85384, n85385, n85386, n85387, n85388,
    n85389, n85390, n85391, n85392, n85393, n85394, n85395, n85396, n85397,
    n85398, n85399, n85400, n85401, n85402, n85403, n85404, n85406, n85407,
    n85408, n85409, n85410, n85411, n85412, n85413, n85414, n85415, n85416,
    n85417, n85418, n85419, n85420, n85421, n85422, n85423, n85424, n85425,
    n85426, n85427, n85428, n85429, n85430, n85431, n85432, n85433, n85434,
    n85435, n85436, n85437, n85438, n85439, n85440, n85441, n85442, n85443,
    n85444, n85445, n85446, n85447, n85448, n85449, n85450, n85451, n85452,
    n85453, n85454, n85455, n85456, n85457, n85458, n85459, n85460, n85461,
    n85462, n85463, n85464, n85465, n85466, n85467, n85468, n85469, n85470,
    n85471, n85472, n85473, n85474, n85475, n85476, n85477, n85478, n85479,
    n85480, n85481, n85482, n85483, n85484, n85485, n85486, n85487, n85488,
    n85489, n85490, n85491, n85492, n85493, n85494, n85495, n85496, n85497,
    n85498, n85499, n85500, n85501, n85502, n85503, n85504, n85505, n85506,
    n85507, n85508, n85509, n85510, n85511, n85512, n85514, n85515, n85516,
    n85517, n85518, n85519, n85520, n85521, n85522, n85523, n85524, n85525,
    n85526, n85527, n85528, n85529, n85530, n85531, n85532, n85533, n85534,
    n85535, n85536, n85537, n85538, n85539, n85540, n85541, n85542, n85543,
    n85544, n85545, n85546, n85547, n85548, n85549, n85550, n85551, n85552,
    n85553, n85554, n85555, n85556, n85557, n85558, n85559, n85560, n85561,
    n85562, n85563, n85564, n85565, n85566, n85567, n85568, n85569, n85570,
    n85571, n85572, n85573, n85574, n85575, n85576, n85577, n85578, n85579,
    n85580, n85581, n85582, n85583, n85584, n85585, n85586, n85587, n85588,
    n85589, n85590, n85591, n85592, n85593, n85594, n85595, n85596, n85597,
    n85598, n85599, n85600, n85601, n85602, n85603, n85604, n85605, n85606,
    n85607, n85608, n85609, n85610, n85611, n85612, n85613, n85614, n85615,
    n85616, n85617, n85618, n85619, n85620, n85621, n85622, n85623, n85624,
    n85625, n85626, n85627, n85628, n85629, n85630, n85631, n85632, n85633,
    n85635, n85636, n85637, n85638, n85639, n85640, n85641, n85642, n85643,
    n85644, n85645, n85646, n85647, n85648, n85649, n85650, n85651, n85652,
    n85653, n85654, n85655, n85656, n85657, n85658, n85659, n85660, n85661,
    n85662, n85663, n85664, n85665, n85666, n85667, n85668, n85669, n85670,
    n85671, n85672, n85673, n85674, n85675, n85676, n85677, n85678, n85679,
    n85680, n85681, n85682, n85683, n85684, n85685, n85686, n85687, n85688,
    n85689, n85690, n85691, n85692, n85693, n85694, n85695, n85696, n85697,
    n85698, n85699, n85700, n85701, n85702, n85703, n85704, n85705, n85706,
    n85707, n85708, n85709, n85710, n85711, n85712, n85713, n85714, n85715,
    n85716, n85717, n85718, n85719, n85720, n85721, n85722, n85723, n85724,
    n85725, n85726, n85727, n85728, n85729, n85730, n85731, n85732, n85733,
    n85734, n85735, n85736, n85737, n85738, n85739, n85740, n85741, n85742,
    n85743, n85744, n85745, n85746, n85747, n85748, n85749, n85750, n85751,
    n85752, n85753, n85754, n85755, n85756, n85757, n85758, n85759, n85760,
    n85761, n85762, n85763, n85764, n85766, n85767, n85768, n85769, n85770,
    n85771, n85772, n85773, n85774, n85775, n85776, n85777, n85778, n85779,
    n85780, n85781, n85782, n85783, n85784, n85785, n85786, n85787, n85788,
    n85789, n85790, n85791, n85792, n85793, n85794, n85795, n85796, n85797,
    n85798, n85799, n85800, n85801, n85802, n85803, n85804, n85805, n85806,
    n85807, n85808, n85809, n85810, n85811, n85812, n85813, n85814, n85815,
    n85816, n85817, n85818, n85819, n85820, n85821, n85822, n85823, n85824,
    n85825, n85826, n85827, n85828, n85829, n85830, n85831, n85832, n85833,
    n85834, n85835, n85836, n85837, n85838, n85839, n85840, n85841, n85842,
    n85843, n85844, n85845, n85846, n85847, n85848, n85849, n85850, n85851,
    n85852, n85853, n85854, n85855, n85856, n85857, n85858, n85859, n85860,
    n85861, n85862, n85863, n85864, n85865, n85866, n85867, n85868, n85869,
    n85870, n85871, n85872, n85873, n85874, n85875, n85876, n85877, n85878,
    n85879, n85880, n85881, n85882, n85883, n85884, n85885, n85886, n85887,
    n85888, n85889, n85890, n85891, n85892, n85893, n85894, n85895, n85896,
    n85897, n85898, n85899, n85900, n85902, n85903, n85904, n85905, n85906,
    n85907, n85908, n85909, n85910, n85911, n85912, n85913, n85914, n85915,
    n85916, n85917, n85918, n85919, n85920, n85921, n85922, n85923, n85924,
    n85925, n85926, n85927, n85928, n85929, n85930, n85931, n85932, n85933,
    n85934, n85935, n85936, n85937, n85938, n85939, n85940, n85941, n85942,
    n85943, n85944, n85945, n85946, n85947, n85948, n85949, n85950, n85951,
    n85952, n85953, n85954, n85955, n85956, n85957, n85958, n85959, n85960,
    n85961, n85962, n85963, n85964, n85965, n85966, n85967, n85968, n85969,
    n85970, n85971, n85972, n85973, n85974, n85975, n85976, n85977, n85978,
    n85979, n85980, n85981, n85982, n85983, n85984, n85985, n85986, n85987,
    n85988, n85989, n85990, n85991, n85992, n85993, n85994, n85995, n85996,
    n85997, n85998, n85999, n86000, n86001, n86002, n86003, n86004, n86005,
    n86006, n86007, n86008, n86009, n86010, n86011, n86012, n86013, n86014,
    n86015, n86016, n86017, n86018, n86019, n86020, n86021, n86022, n86023,
    n86024, n86025, n86026, n86027, n86028, n86029, n86030, n86031, n86032,
    n86033, n86035, n86036, n86037, n86038, n86039, n86040, n86041, n86042,
    n86043, n86044, n86045, n86046, n86047, n86048, n86049, n86050, n86051,
    n86052, n86053, n86054, n86055, n86056, n86057, n86058, n86059, n86060,
    n86061, n86062, n86063, n86064, n86065, n86066, n86067, n86068, n86069,
    n86070, n86071, n86072, n86073, n86074, n86075, n86076, n86077, n86078,
    n86079, n86080, n86081, n86082, n86083, n86084, n86085, n86086, n86087,
    n86088, n86089, n86090, n86091, n86092, n86093, n86094, n86095, n86096,
    n86097, n86098, n86099, n86100, n86101, n86102, n86103, n86104, n86105,
    n86106, n86107, n86108, n86109, n86110, n86111, n86112, n86113, n86114,
    n86115, n86116, n86117, n86118, n86119, n86120, n86121, n86122, n86123,
    n86124, n86125, n86126, n86127, n86128, n86129, n86130, n86131, n86132,
    n86133, n86134, n86135, n86136, n86137, n86138, n86139, n86140, n86141,
    n86142, n86143, n86144, n86145, n86146, n86147, n86148, n86149, n86150,
    n86151, n86152, n86153, n86154, n86155, n86156, n86157, n86158, n86159,
    n86160, n86161, n86162, n86163, n86164, n86166, n86167, n86168, n86169,
    n86170, n86171, n86172, n86173, n86174, n86175, n86176, n86177, n86178,
    n86179, n86180, n86181, n86182, n86183, n86184, n86185, n86186, n86187,
    n86188, n86189, n86190, n86191, n86192, n86193, n86194, n86195, n86196,
    n86197, n86198, n86199, n86200, n86201, n86202, n86203, n86204, n86205,
    n86206, n86207, n86208, n86209, n86210, n86211, n86212, n86213, n86214,
    n86215, n86216, n86217, n86218, n86219, n86220, n86221, n86222, n86223,
    n86224, n86225, n86226, n86227, n86228, n86229, n86230, n86231, n86232,
    n86233, n86234, n86235, n86236, n86237, n86238, n86239, n86240, n86241,
    n86242, n86243, n86244, n86245, n86246, n86247, n86248, n86249, n86250,
    n86251, n86252, n86253, n86254, n86255, n86256, n86257, n86258, n86259,
    n86260, n86261, n86262, n86264, n86265, n86266, n86267, n86268, n86269,
    n86270, n86271, n86272, n86273, n86274, n86275, n86276, n86277, n86278,
    n86279, n86280, n86281, n86282, n86283, n86284, n86285, n86286, n86287,
    n86288, n86289, n86290, n86291, n86292, n86293, n86294, n86295, n86296,
    n86297, n86298, n86299, n86300, n86301, n86302, n86303, n86304, n86305,
    n86306, n86307, n86308, n86309, n86310, n86311, n86312, n86313, n86314,
    n86315, n86316, n86317, n86318, n86319, n86320, n86321, n86322, n86323,
    n86324, n86325, n86326, n86327, n86328, n86329, n86330, n86331, n86332,
    n86333, n86334, n86335, n86336, n86337, n86338, n86339, n86340, n86341,
    n86342, n86343, n86344, n86345, n86346, n86347, n86348, n86349, n86350,
    n86351, n86352, n86354, n86355, n86356, n86357, n86358, n86359, n86360,
    n86361, n86362, n86363, n86364, n86365, n86366, n86367, n86368, n86369,
    n86370, n86371, n86372, n86373, n86374, n86375, n86376, n86377, n86378,
    n86379, n86380, n86381, n86382, n86383, n86384, n86385, n86386, n86387,
    n86388, n86389, n86390, n86391, n86392, n86393, n86394, n86395, n86396,
    n86397, n86398, n86399, n86400, n86401, n86402, n86403, n86404, n86405,
    n86406, n86407, n86408, n86409, n86410, n86411, n86412, n86413, n86414,
    n86415, n86416, n86417, n86418, n86419, n86420, n86421, n86422, n86423,
    n86424, n86425, n86426, n86427, n86428, n86429, n86430, n86431, n86432,
    n86433, n86434, n86435, n86437, n86438, n86439, n86440, n86441, n86442,
    n86443, n86444, n86445, n86446, n86447, n86448, n86449, n86450, n86451,
    n86452, n86453, n86454, n86455, n86456, n86457, n86458, n86459, n86460,
    n86461, n86462, n86463, n86464, n86465, n86466, n86467, n86468, n86469,
    n86470, n86471, n86472, n86473, n86474, n86475, n86476, n86477, n86478,
    n86479, n86480, n86481, n86482, n86483, n86484, n86485, n86486, n86487,
    n86488, n86489, n86490, n86491, n86492, n86493, n86494, n86495, n86496,
    n86497, n86498, n86499, n86500, n86501, n86502, n86503, n86504, n86505,
    n86506, n86507, n86508, n86509, n86510, n86511, n86513, n86514, n86515,
    n86516, n86517, n86518, n86519, n86520, n86521, n86522, n86523, n86524,
    n86525, n86526, n86527, n86528, n86529, n86530, n86531, n86532, n86533,
    n86534, n86535, n86536, n86537, n86538, n86539, n86540, n86541, n86542,
    n86543, n86544, n86545, n86546, n86547, n86548, n86549, n86550, n86551,
    n86552, n86553, n86554, n86555, n86556, n86557, n86558, n86559, n86560,
    n86561, n86562, n86563, n86564, n86565, n86566, n86567, n86568, n86569,
    n86570, n86571, n86572, n86573, n86574, n86575, n86576, n86577, n86578,
    n86579, n86580, n86581, n86582, n86583, n86585, n86586, n86587, n86588,
    n86589, n86590, n86591, n86592, n86593, n86594, n86595, n86596, n86597,
    n86598, n86599, n86600, n86601, n86602, n86603, n86604, n86605, n86606,
    n86607, n86608, n86609, n86610, n86611, n86612, n86613, n86614, n86615,
    n86616, n86617, n86618, n86619, n86620, n86621, n86622, n86623, n86624,
    n86625, n86626, n86627, n86628, n86629, n86630, n86631, n86632, n86633,
    n86634, n86635, n86636, n86637, n86638, n86639, n86640, n86641, n86642,
    n86643, n86644, n86645, n86646, n86647, n86648, n86649, n86650, n86651,
    n86652, n86653, n86654, n86655, n86656, n86657, n86658, n86659, n86660,
    n86661, n86663, n86664, n86665, n86666, n86667, n86668, n86669, n86670,
    n86671, n86672, n86673, n86674, n86675, n86676, n86677, n86678, n86679,
    n86680, n86681, n86682, n86683, n86684, n86685, n86686, n86687, n86688,
    n86689, n86690, n86691, n86692, n86693, n86694, n86695, n86696, n86697,
    n86698, n86699, n86700, n86701, n86702, n86703, n86704, n86705, n86706,
    n86707, n86708, n86709, n86710, n86711, n86712, n86713, n86714, n86715,
    n86716, n86717, n86718, n86719, n86720, n86721, n86722, n86723, n86724,
    n86725, n86726, n86727, n86728, n86729, n86730, n86731, n86732, n86733,
    n86734, n86735, n86736, n86738, n86739, n86740, n86741, n86742, n86743,
    n86744, n86745, n86746, n86747, n86748, n86749, n86750, n86751, n86752,
    n86753, n86754, n86755, n86756, n86757, n86758, n86759, n86760, n86761,
    n86762, n86763, n86764, n86765, n86766, n86767, n86768, n86769, n86770,
    n86771, n86772, n86773, n86774, n86775, n86776, n86777, n86778, n86779,
    n86780, n86781, n86782, n86783, n86784, n86785, n86786, n86787, n86788,
    n86789, n86790, n86791, n86792, n86793, n86794, n86795, n86796, n86797,
    n86798, n86799, n86800, n86801, n86802, n86803, n86804, n86805, n86806,
    n86807, n86808, n86809, n86811, n86812, n86813, n86814, n86815, n86816,
    n86817, n86818, n86819, n86820, n86821, n86822, n86823, n86824, n86825,
    n86826, n86827, n86828, n86829, n86830, n86831, n86832, n86833, n86834,
    n86835, n86836, n86837, n86838, n86839, n86840, n86841, n86842, n86843,
    n86844, n86845, n86846, n86847, n86848, n86849, n86850, n86851, n86852,
    n86853, n86854, n86855, n86856, n86857, n86858, n86859, n86860, n86861,
    n86862, n86863, n86864, n86865, n86866, n86867, n86868, n86869, n86870,
    n86871, n86872, n86873, n86874, n86875, n86876, n86877, n86878, n86879,
    n86880, n86881, n86882, n86883, n86884, n86885, n86886, n86887, n86889,
    n86890, n86891, n86892, n86893, n86894, n86895, n86896, n86897, n86898,
    n86899, n86900, n86901, n86902, n86903, n86904, n86905, n86906, n86907,
    n86908, n86909, n86910, n86911, n86912, n86913, n86914, n86915, n86916,
    n86917, n86918, n86919, n86920, n86921, n86922, n86923, n86924, n86925,
    n86926, n86927, n86928, n86929, n86930, n86931, n86932, n86933, n86934,
    n86935, n86936, n86937, n86938, n86939, n86940, n86941, n86942, n86943,
    n86944, n86945, n86946, n86947, n86948, n86949, n86950, n86951, n86952,
    n86953, n86954, n86955, n86956, n86957, n86958, n86959, n86961, n86962,
    n86963, n86964, n86965, n86966, n86967, n86968, n86969, n86970, n86971,
    n86972, n86973, n86974, n86975, n86976, n86977, n86978, n86979, n86980,
    n86981, n86982, n86983, n86984, n86985, n86986, n86987, n86988, n86989,
    n86990, n86991, n86992, n86993, n86994, n86995, n86996, n86997, n86998,
    n86999, n87000, n87001, n87002, n87003, n87004, n87005, n87006, n87007,
    n87008, n87009, n87010, n87011, n87012, n87013, n87014, n87015, n87016,
    n87017, n87018, n87019, n87020, n87021, n87022, n87023, n87024, n87025,
    n87026, n87027, n87028, n87029, n87030, n87031, n87032, n87033, n87034,
    n87035, n87036, n87037, n87038, n87040, n87041, n87042, n87043, n87044,
    n87045, n87046, n87047, n87048, n87049, n87050, n87051, n87052, n87053,
    n87054, n87055, n87056, n87057, n87058, n87059, n87060, n87061, n87062,
    n87063, n87064, n87065, n87066, n87067, n87068, n87069, n87070, n87071,
    n87072, n87073, n87074, n87075, n87076, n87077, n87078, n87079, n87080,
    n87081, n87082, n87083, n87084, n87085, n87086, n87087, n87088, n87089,
    n87090, n87091, n87092, n87093, n87094, n87095, n87096, n87097, n87098,
    n87099, n87100, n87101, n87102, n87103, n87104, n87105, n87106, n87107,
    n87108, n87109, n87111, n87112, n87113, n87114, n87115, n87116, n87117,
    n87118, n87119, n87120, n87121, n87122, n87123, n87124, n87125, n87126,
    n87127, n87128, n87129, n87130, n87131, n87132, n87133, n87134, n87135,
    n87136, n87137, n87138, n87139, n87140, n87141, n87142, n87143, n87144,
    n87145, n87146, n87147, n87148, n87149, n87150, n87151, n87152, n87153,
    n87154, n87155, n87156, n87157, n87158, n87159, n87160, n87161, n87162,
    n87163, n87164, n87165, n87166, n87167, n87168, n87169, n87170, n87171,
    n87172, n87173, n87174, n87175, n87176, n87177, n87178, n87179, n87180,
    n87181, n87182, n87183, n87184, n87185, n87186, n87187, n87189, n87190,
    n87191, n87192, n87193, n87194, n87195, n87196, n87197, n87198, n87199,
    n87200, n87201, n87202, n87203, n87204, n87205, n87206, n87207, n87208,
    n87209, n87210, n87211, n87212, n87213, n87214, n87215, n87216, n87217,
    n87218, n87219, n87220, n87221, n87222, n87223, n87224, n87225, n87226,
    n87227, n87228, n87229, n87230, n87231, n87232, n87233, n87234, n87235,
    n87236, n87237, n87238, n87239, n87240, n87241, n87242, n87243, n87244,
    n87245, n87246, n87247, n87248, n87249, n87250, n87251, n87252, n87253,
    n87254, n87255, n87256, n87257, n87258, n87259, n87260, n87261, n87262,
    n87263, n87265, n87266, n87267, n87268, n87269, n87270, n87271, n87272,
    n87273, n87274, n87275, n87276, n87277, n87278, n87279, n87280, n87281,
    n87282, n87283, n87284, n87285, n87286, n87287, n87288, n87289, n87290,
    n87291, n87292, n87293, n87294, n87295, n87296, n87297, n87298, n87299,
    n87300, n87301, n87302, n87303, n87304, n87305, n87306, n87307, n87308,
    n87309, n87310, n87311, n87312, n87313, n87314, n87315, n87316, n87317,
    n87318, n87319, n87320, n87321, n87322, n87323, n87324, n87325, n87326,
    n87327, n87328, n87329, n87330, n87331, n87332, n87333, n87334, n87335,
    n87336, n87338, n87339, n87340, n87341, n87342, n87343, n87344, n87345,
    n87346, n87347, n87348, n87349, n87350, n87351, n87352, n87353, n87354,
    n87355, n87356, n87357, n87358, n87359, n87360, n87361, n87362, n87363,
    n87364, n87365, n87366, n87367, n87368, n87369, n87370, n87371, n87372,
    n87373, n87374, n87375, n87376, n87377, n87378, n87379, n87380, n87381,
    n87382, n87383, n87384, n87385, n87386, n87387, n87388, n87389, n87390,
    n87391, n87392, n87393, n87394, n87395, n87396, n87397, n87398, n87399,
    n87400, n87401, n87402, n87403, n87404, n87405, n87406, n87407, n87408,
    n87409, n87410, n87411, n87412, n87413, n87415, n87416, n87417, n87418,
    n87419, n87420, n87421, n87422, n87423, n87424, n87425, n87426, n87427,
    n87428, n87429, n87430, n87431, n87432, n87433, n87434, n87435, n87436,
    n87437, n87438, n87439, n87440, n87441, n87442, n87443, n87444, n87445,
    n87446, n87447, n87448, n87449, n87450, n87451, n87452, n87453, n87454,
    n87455, n87456, n87457, n87458, n87459, n87460, n87461, n87462, n87463,
    n87464, n87465, n87466, n87467, n87468, n87469, n87470, n87471, n87472,
    n87473, n87474, n87475, n87476, n87477, n87478, n87479, n87480, n87481,
    n87482, n87483, n87484, n87485, n87486, n87487, n87488, n87489, n87490,
    n87492, n87493, n87494, n87495, n87496, n87497, n87498, n87499, n87500,
    n87501, n87502, n87503, n87504, n87505, n87506, n87507, n87508, n87509,
    n87510, n87511, n87512, n87513, n87514, n87515, n87516, n87517, n87518,
    n87519, n87520, n87521, n87522, n87523, n87524, n87525, n87526, n87527,
    n87528, n87529, n87530, n87531, n87532, n87533, n87534, n87535, n87536,
    n87537, n87538, n87539, n87540, n87541, n87542, n87543, n87544, n87545,
    n87546, n87547, n87548, n87549, n87550, n87551, n87552, n87553, n87554,
    n87555, n87556, n87557, n87558, n87559, n87560, n87561, n87562, n87563,
    n87564, n87566, n87567, n87568, n87569, n87570, n87571, n87572, n87573,
    n87574, n87575, n87576, n87577, n87578, n87579, n87580, n87581, n87582,
    n87583, n87584, n87585, n87586, n87587, n87588, n87589, n87590, n87591,
    n87592, n87593, n87594, n87595, n87596, n87597, n87598, n87599, n87600,
    n87601, n87602, n87603, n87604, n87605, n87606, n87607, n87608, n87609,
    n87610, n87611, n87612, n87613, n87614, n87615, n87616, n87617, n87618,
    n87619, n87620, n87621, n87622, n87623, n87624, n87625, n87626, n87627,
    n87628, n87629, n87630, n87631, n87632, n87633, n87634, n87635, n87636,
    n87637, n87638, n87639, n87640, n87641, n87642, n87644, n87645, n87646,
    n87647, n87648, n87649, n87650, n87651, n87652, n87653, n87654, n87655,
    n87656, n87657, n87658, n87659, n87660, n87661, n87662, n87663, n87664,
    n87665, n87666, n87667, n87668, n87669, n87670, n87671, n87672, n87673,
    n87674, n87675, n87676, n87677, n87678, n87679, n87680, n87681, n87682,
    n87683, n87684, n87685, n87686, n87687, n87688, n87689, n87690, n87691,
    n87692, n87693, n87694, n87695, n87696, n87697, n87698, n87699, n87700,
    n87701, n87702, n87703, n87704, n87705, n87706, n87707, n87708, n87709,
    n87710, n87711, n87712, n87713, n87714, n87715, n87716, n87717, n87719,
    n87720, n87721, n87722, n87723, n87724, n87725, n87726, n87727, n87728,
    n87729, n87730, n87731, n87732, n87733, n87734, n87735, n87736, n87737,
    n87738, n87739, n87740, n87741, n87742, n87743, n87744, n87745, n87746,
    n87747, n87748, n87749, n87750, n87751, n87752, n87753, n87754, n87755,
    n87756, n87757, n87758, n87759, n87760, n87761, n87762, n87763, n87764,
    n87765, n87766, n87767, n87768, n87769, n87770, n87771, n87772, n87773,
    n87774, n87775, n87776, n87777, n87778, n87779, n87780, n87781, n87782,
    n87783, n87784, n87785, n87786, n87787, n87788, n87790, n87791, n87792,
    n87793, n87794, n87795, n87796, n87797, n87798, n87799, n87800, n87801,
    n87802, n87803, n87804, n87805, n87806, n87807, n87808, n87809, n87810,
    n87811, n87812, n87813, n87814, n87815, n87816, n87817, n87818, n87819,
    n87820, n87821, n87822, n87823, n87824, n87825, n87826, n87827, n87828,
    n87829, n87830, n87831, n87832, n87833, n87834, n87835, n87836, n87837,
    n87838, n87839, n87840, n87841, n87842, n87843, n87844, n87845, n87846,
    n87847, n87848, n87849, n87850, n87851, n87852, n87853, n87854, n87855,
    n87856, n87857, n87858, n87859, n87860, n87861, n87862, n87863, n87864,
    n87865, n87866, n87867, n87868, n87870, n87871, n87872, n87873, n87874,
    n87875, n87876, n87877, n87878, n87879, n87880, n87881, n87882, n87883,
    n87884, n87885, n87886, n87887, n87888, n87889, n87890, n87891, n87892,
    n87893, n87894, n87895, n87896, n87897, n87898, n87899, n87900, n87901,
    n87902, n87903, n87904, n87905, n87906, n87907, n87908, n87909, n87910,
    n87911, n87912, n87913, n87914, n87915, n87916, n87917, n87918, n87919,
    n87920, n87921, n87922, n87923, n87924, n87925, n87926, n87927, n87928,
    n87929, n87930, n87931, n87932, n87933, n87934, n87935, n87936, n87937,
    n87938, n87939, n87941, n87942, n87943, n87944, n87945, n87946, n87947,
    n87948, n87949, n87950, n87951, n87952, n87953, n87954, n87955, n87956,
    n87957, n87958, n87959, n87960, n87961, n87962, n87963, n87964, n87965,
    n87966, n87967, n87968, n87969, n87970, n87971, n87972, n87973, n87974,
    n87975, n87976, n87977, n87978, n87979, n87980, n87981, n87982, n87983,
    n87984, n87985, n87986, n87987, n87988, n87989, n87990, n87991, n87992,
    n87993, n87994, n87995, n87996, n87997, n87998, n87999, n88000, n88001,
    n88002, n88003, n88004, n88005, n88006, n88007, n88008, n88009, n88010,
    n88011, n88013, n88014, n88015, n88016, n88017, n88018, n88019, n88020,
    n88021, n88022, n88023, n88024, n88025, n88026, n88027, n88028, n88029,
    n88030, n88031, n88032, n88033, n88034, n88035, n88036, n88037, n88038,
    n88039, n88040, n88041, n88042, n88043, n88044, n88045, n88046, n88047,
    n88048, n88049, n88050, n88051, n88052, n88053, n88054, n88055, n88056,
    n88057, n88058, n88059, n88060, n88061, n88062, n88063, n88064, n88065,
    n88066, n88067, n88068, n88069, n88070, n88071, n88072, n88073, n88074,
    n88075, n88076, n88077, n88078, n88079, n88080, n88081, n88082, n88083,
    n88084, n88085, n88086, n88087, n88088, n88089, n88090, n88091, n88093,
    n88094, n88095, n88096, n88097, n88098, n88099, n88100, n88101, n88102,
    n88103, n88104, n88105, n88106, n88107, n88108, n88109, n88110, n88111,
    n88112, n88113, n88114, n88115, n88116, n88117, n88118, n88119, n88120,
    n88121, n88122, n88123, n88124, n88126, n88127, n88128, n88129, n88130,
    n88131, n88132, n88133, n88134, n88135, n88136, n88137, n88138, n88139,
    n88141, n88142, n88143, n88144, n88145, n88146, n88147, n88148, n88149,
    n88150, n88151, n88152, n88153, n88154, n88155, n88156, n88157, n88159,
    n88160, n88161, n88162, n88163, n88164, n88165, n88166, n88167, n88168,
    n88169, n88170, n88171, n88172, n88173, n88174, n88175, n88176, n88177,
    n88178, n88179, n88181, n88182, n88183, n88184, n88185, n88186, n88187,
    n88188, n88189, n88190, n88191, n88192, n88193, n88194, n88195, n88196,
    n88197, n88198, n88199, n88200, n88201, n88202, n88204, n88205, n88206,
    n88207, n88208, n88209, n88210, n88211, n88212, n88213, n88214, n88215,
    n88216, n88217, n88218, n88219, n88220, n88221, n88222, n88223, n88224,
    n88225, n88227, n88228, n88229, n88230, n88231, n88232, n88233, n88234,
    n88235, n88236, n88237, n88238, n88239, n88240, n88241, n88242, n88243,
    n88244, n88245, n88246, n88247, n88248, n88250, n88251, n88252, n88253,
    n88254, n88255, n88256, n88257, n88258, n88259, n88260, n88261, n88262,
    n88263, n88264, n88265, n88266, n88267, n88268, n88269, n88270, n88271,
    n88273, n88274, n88275, n88276, n88277, n88278, n88279, n88280, n88281,
    n88282, n88283, n88284, n88285, n88286, n88287, n88288, n88289, n88290,
    n88291, n88292, n88293, n88294, n88296, n88297, n88298, n88299, n88300,
    n88301, n88302, n88303, n88304, n88305, n88306, n88307, n88308, n88309,
    n88310, n88311, n88312, n88313, n88314, n88315, n88316, n88317, n88319,
    n88320, n88321, n88322, n88323, n88324, n88325, n88326, n88327, n88328,
    n88329, n88330, n88331, n88332, n88333, n88334, n88335, n88336, n88337,
    n88338, n88339, n88340, n88342, n88343, n88344, n88345, n88346, n88347,
    n88348, n88349, n88350, n88351, n88352, n88353, n88354, n88355, n88356,
    n88357, n88358, n88359, n88360, n88361, n88362, n88363, n88365, n88366,
    n88367, n88368, n88369, n88370, n88371, n88372, n88373, n88374, n88375,
    n88376, n88377, n88378, n88379, n88380, n88381, n88382, n88383, n88384,
    n88385, n88386, n88388, n88389, n88390, n88391, n88392, n88393, n88394,
    n88395, n88396, n88397, n88398, n88399, n88400, n88401, n88402, n88403,
    n88404, n88405, n88406, n88407, n88408, n88409, n88411, n88412, n88413,
    n88414, n88415, n88416, n88417, n88418, n88419, n88420, n88421, n88422,
    n88423, n88424, n88425, n88426, n88427, n88428, n88429, n88430, n88431,
    n88432, n88434, n88435, n88436, n88437, n88438, n88439, n88440, n88441,
    n88442, n88443, n88444, n88445, n88446, n88447, n88448, n88449, n88450,
    n88451, n88452, n88453, n88454, n88455, n88457, n88458, n88459, n88460,
    n88461, n88462, n88463, n88464, n88465, n88466, n88467, n88468, n88469,
    n88470, n88471, n88472, n88473, n88474, n88475, n88476, n88477, n88478,
    n88480, n88481, n88482, n88483, n88484, n88485, n88486, n88487, n88488,
    n88489, n88490, n88491, n88492, n88493, n88494, n88495, n88496, n88497,
    n88498, n88499, n88500, n88501, n88503, n88504, n88505, n88506, n88507,
    n88508, n88509, n88510, n88511, n88512, n88513, n88514, n88515, n88516,
    n88517, n88518, n88519, n88520, n88521, n88522, n88523, n88524, n88526,
    n88527, n88528, n88529, n88530, n88531, n88532, n88533, n88534, n88535,
    n88536, n88537, n88538, n88539, n88540, n88541, n88542, n88543, n88544,
    n88545, n88546, n88547, n88549, n88550, n88551, n88552, n88553, n88554,
    n88555, n88556, n88557, n88558, n88559, n88560, n88561, n88562, n88563,
    n88564, n88565, n88566, n88567, n88568, n88569, n88570, n88572, n88573,
    n88574, n88575, n88576, n88577, n88578, n88579, n88580, n88581, n88582,
    n88583, n88584, n88585, n88586, n88587, n88588, n88589, n88590, n88591,
    n88592, n88593, n88595, n88596, n88597, n88598, n88599, n88600, n88601,
    n88602, n88603, n88604, n88605, n88606, n88607, n88608, n88609, n88610,
    n88611, n88612, n88613, n88614, n88615, n88616, n88618, n88619, n88620,
    n88621, n88622, n88623, n88624, n88625, n88626, n88627, n88628, n88629,
    n88630, n88631, n88632, n88633, n88634, n88635, n88636, n88637, n88638,
    n88639, n88641, n88642, n88643, n88644, n88645, n88646, n88647, n88648,
    n88649, n88650, n88651, n88652, n88653, n88654, n88655, n88656, n88657,
    n88658, n88659, n88660, n88661, n88662, n88664, n88665, n88666, n88667,
    n88668, n88669, n88670, n88671, n88672, n88673, n88674, n88675, n88676,
    n88677, n88678, n88679, n88680, n88681, n88682, n88683, n88684, n88685,
    n88687, n88688, n88689, n88690, n88691, n88692, n88693, n88694, n88695,
    n88696, n88697, n88698, n88699, n88700, n88701, n88702, n88703, n88704,
    n88705, n88706, n88707, n88708, n88710, n88711, n88712, n88713, n88714,
    n88715, n88716, n88717, n88718, n88719, n88720, n88721, n88722, n88723,
    n88724, n88725, n88726, n88727, n88728, n88729, n88730, n88731, n88733,
    n88734, n88735, n88736, n88737, n88738, n88739, n88740, n88741, n88742,
    n88743, n88744, n88745, n88746, n88747, n88748, n88749, n88750, n88751,
    n88752, n88753, n88754, n88756, n88757, n88758, n88759, n88760, n88761,
    n88762, n88763, n88764, n88765, n88766, n88767, n88768, n88769, n88770,
    n88771, n88772, n88773, n88774, n88775, n88776, n88777, n88779, n88780,
    n88781, n88782, n88783, n88784, n88785, n88786, n88787, n88788, n88789,
    n88790, n88791, n88792, n88793, n88794, n88795, n88796, n88797, n88798,
    n88799, n88800, n88802, n88803, n88804, n88805, n88806, n88807, n88808,
    n88809, n88810, n88811, n88812, n88813, n88814, n88815, n88816, n88817,
    n88818, n88819, n88820, n88821, n88822, n88823, n88825, n88826, n88827,
    n88828, n88829, n88830, n88831, n88832, n88833, n88834, n88835, n88836,
    n88837, n88838, n88839, n88840, n88841, n88842, n88843, n88844, n88846,
    n88847, n88848, n88849, n88850, n88851, n88852, n88853, n88854, n88855,
    n88856, n88857, n88858, n88859, n88860, n88862, n88863, n88864, n88865,
    n88866, n88867, n88868, n88869, n88870, n88871, n88872, n88873, n88874,
    n88876, n88877, n88878, n88879, n88880, n88881, n88882, n88883, n88884,
    n88885, n88886, n88887, n88888, n88889, n88890, n88892, n88893, n88894,
    n88895, n88896, n88897, n88898, n88899, n88900, n88901, n88902, n88903,
    n88904, n88905, n88907, n88908, n88909, n88910, n88911, n88912, n88913,
    n88914, n88915, n88916, n88917, n88918, n88919, n88920, n88921, n88923,
    n88924, n88925, n88926, n88927, n88928, n88929, n88930, n88931, n88932,
    n88933, n88935, n88936, n88937, n88938, n88939, n88940, n88941, n88942,
    n88943, n88944, n88945, n88946, n88947, n88948, n88949, n88950, n88952,
    n88953, n88954, n88955, n88957, n88958, n88959, n88960, n88962, n88963,
    n88964, n88965, n88967, n88968, n88969, n88970, n88972, n88973, n88974,
    n88975, n88977, n88978, n88979, n88980, n88982, n88983, n88984, n88985,
    n88987, n88988, n88989, n88990, n88992, n88993, n88994, n88996, n88997,
    n88998, n89000, n89001, n89002, n89004, n89005, n89006, n89008, n89009,
    n89010, n89012, n89013, n89014, n89016, n89017, n89018, n89020, n89021,
    n89022, n89024, n89025, n89026, n89028, n89029, n89030, n89032, n89033,
    n89034, n89036, n89037, n89038, n89040, n89041, n89042, n89044, n89045,
    n89046, n89048, n89049, n89050, n89052, n89053, n89054, n89055, n89056,
    n89057, n89058, n89059, n89060, n89061, n89063, n89064, n89065, n89066,
    n89068, n89069, n89070, n89071, n89073, n89074, n89075, n89076, n89078,
    n89079, n89080, n89081, n89083, n89084, n89085, n89086, n89088, n89089,
    n89090, n89091, n89093, n89094, n89095, n89096, n89098, n89099, n89100,
    n89101, n89103, n89104, n89105, n89106, n89108, n89109, n89110, n89111,
    n89113, n89114, n89115, n89116, n89118, n89119, n89120, n89121, n89123,
    n89124, n89125, n89126, n89128, n89129, n89130, n89131, n89133, n89134,
    n89135, n89136, n89138, n89139, n89140, n89141, n89142, n89144, n89145,
    n89146, n89147, n89149, n89150, n89151, n89152, n89154, n89155, n89156,
    n89157, n89159, n89160, n89161, n89162, n89164, n89165, n89166, n89167,
    n89169, n89170, n89171, n89172, n89174, n89175, n89176, n89177, n89179,
    n89180, n89181, n89182, n89184, n89185, n89186, n89187, n89189, n89190,
    n89191, n89192, n89194, n89195, n89196, n89197, n89199, n89200, n89201,
    n89202, n89204, n89205, n89206, n89207, n89209, n89210, n89211, n89212,
    n89215, n89216, n89217, n89218, n89219, n89220, n89221, n89222, n89223,
    n89224, n89225, n89226, n89228, n89229, n89230, n89231, n89232, n89233,
    n89234, n89235, n89236, n89238, n89239, n89240, n89241, n89242, n89243,
    n89244, n89245, n89246, n89247, n89249, n89250, n89251, n89252, n89253,
    n89254, n89255, n89256, n89257, n89258, n89260, n89261, n89262, n89263,
    n89264, n89265, n89266, n89267, n89268, n89269, n89271, n89272, n89273,
    n89274, n89275, n89276, n89277, n89278, n89279, n89280, n89282, n89283,
    n89284, n89285, n89286, n89287, n89288, n89289, n89290, n89291, n89293,
    n89294, n89295, n89296, n89297, n89298, n89299, n89300, n89301, n89302,
    n89304, n89305, n89306, n89307, n89308, n89309, n89310, n89311, n89312,
    n89313, n89314, n89315, n89316, n89317, n89318, n89319, n89320, n89321,
    n89322, n89323, n89324, n89325, n89326, n89327, n89328, n89329, n89330,
    n89331, n89332, n89333, n89334, n89335, n89336, n89337, n89338, n89339,
    n89340, n89341, n89342, n89343, n89344, n89345, n89346, n89347, n89348,
    n89349, n89350, n89351, n89352, n89353, n89354, n89355, n89356, n89357,
    n89358, n89359, n89360, n89361, n89362, n89363, n89364, n89365, n89367,
    n89368, n89369, n89370, n89371, n89372, n89373, n89374, n89375, n89376,
    n89377, n89378, n89379, n89380, n89381, n89382, n89383, n89384, n89385,
    n89386, n89387, n89388, n89389, n89390, n89391, n89392, n89393, n89394,
    n89395, n89396, n89397, n89398, n89399, n89400, n89401, n89402, n89403,
    n89404, n89405, n89406, n89407, n89409, n89410, n89411, n89412, n89413,
    n89414, n89415, n89416, n89417, n89418, n89419, n89420, n89421, n89422,
    n89423, n89424, n89425, n89426, n89427, n89428, n89429, n89430, n89431,
    n89432, n89433, n89434, n89435, n89436, n89437, n89438, n89439, n89440,
    n89441, n89442, n89443, n89444, n89445, n89446, n89447, n89448, n89449,
    n89451, n89452, n89453, n89454, n89455, n89456, n89457, n89458, n89459,
    n89460, n89461, n89462, n89463, n89464, n89465, n89466, n89467, n89468,
    n89469, n89470, n89471, n89472, n89473, n89474, n89475, n89476, n89477,
    n89478, n89479, n89480, n89481, n89482, n89483, n89484, n89485, n89486,
    n89487, n89488, n89489, n89490, n89491, n89493, n89494, n89495, n89496,
    n89497, n89498, n89499, n89500, n89501, n89502, n89503, n89504, n89505,
    n89506, n89507, n89508, n89509, n89510, n89511, n89512, n89513, n89514,
    n89515, n89516, n89517, n89518, n89519, n89520, n89521, n89522, n89523,
    n89524, n89525, n89526, n89527, n89528, n89529, n89530, n89531, n89532,
    n89533, n89535, n89536, n89537, n89538, n89539, n89540, n89541, n89542,
    n89543, n89544, n89545, n89546, n89547, n89548, n89549, n89550, n89551,
    n89552, n89553, n89554, n89555, n89556, n89557, n89558, n89559, n89560,
    n89561, n89562, n89563, n89564, n89565, n89566, n89567, n89568, n89569,
    n89570, n89571, n89572, n89573, n89574, n89575, n89577, n89578, n89579,
    n89580, n89581, n89582, n89583, n89584, n89585, n89586, n89587, n89588,
    n89589, n89590, n89591, n89592, n89593, n89594, n89595, n89596, n89597,
    n89598, n89599, n89600, n89601, n89602, n89603, n89604, n89605, n89606,
    n89607, n89608, n89609, n89610, n89611, n89612, n89613, n89614, n89615,
    n89616, n89617, n89619, n89620, n89621, n89622, n89623, n89624, n89625,
    n89626, n89627, n89628, n89629, n89630, n89631, n89632, n89633, n89634,
    n89635, n89636, n89637, n89638, n89639, n89640, n89641, n89642, n89643,
    n89644, n89645, n89646, n89647, n89648, n89649, n89650, n89651, n89652,
    n89653, n89654, n89655, n89656, n89657, n89658, n89659, n89661, n89662,
    n89663, n89664, n89665, n89666, n89667, n89668, n89669, n89670, n89671,
    n89672, n89673, n89674, n89675, n89676, n89677, n89678, n89679, n89680,
    n89681, n89682, n89683, n89684, n89685, n89686, n89687, n89688, n89689,
    n89690, n89691, n89692, n89693, n89694, n89695, n89696, n89697, n89698,
    n89699, n89700, n89701, n89702, n89703, n89704, n89705, n89706, n89707,
    n89708, n89709, n89710, n89711, n89712, n89713, n89714, n89715, n89716,
    n89717, n89718, n89719, n89720, n89721, n89722, n89723, n89724, n89725,
    n89726, n89727, n89728, n89729, n89730, n89732, n89733, n89734, n89735,
    n89736, n89737, n89738, n89739, n89740, n89741, n89742, n89743, n89744,
    n89745, n89746, n89747, n89748, n89749, n89750, n89751, n89752, n89753,
    n89754, n89755, n89756, n89757, n89758, n89759, n89760, n89761, n89762,
    n89763, n89764, n89765, n89766, n89767, n89768, n89769, n89770, n89771,
    n89772, n89773, n89774, n89776, n89777, n89778, n89779, n89780, n89781,
    n89782, n89783, n89784, n89785, n89786, n89787, n89788, n89789, n89790,
    n89791, n89792, n89793, n89794, n89795, n89796, n89797, n89798, n89799,
    n89800, n89801, n89802, n89803, n89804, n89805, n89806, n89807, n89808,
    n89809, n89810, n89811, n89812, n89813, n89814, n89815, n89816, n89817,
    n89818, n89820, n89821, n89822, n89823, n89824, n89825, n89826, n89827,
    n89828, n89829, n89830, n89831, n89832, n89833, n89834, n89835, n89836,
    n89837, n89838, n89839, n89840, n89841, n89842, n89843, n89844, n89845,
    n89846, n89847, n89848, n89849, n89850, n89851, n89852, n89853, n89854,
    n89855, n89856, n89857, n89858, n89859, n89860, n89861, n89862, n89864,
    n89865, n89866, n89867, n89868, n89869, n89870, n89871, n89872, n89873,
    n89874, n89875, n89876, n89877, n89878, n89879, n89880, n89881, n89882,
    n89883, n89884, n89885, n89886, n89887, n89888, n89889, n89890, n89891,
    n89892, n89893, n89894, n89895, n89896, n89897, n89898, n89899, n89900,
    n89901, n89902, n89903, n89904, n89905, n89906, n89908, n89909, n89910,
    n89911, n89912, n89913, n89914, n89915, n89916, n89917, n89918, n89919,
    n89920, n89921, n89922, n89923, n89924, n89925, n89926, n89927, n89928,
    n89929, n89930, n89931, n89932, n89933, n89934, n89935, n89936, n89937,
    n89938, n89939, n89940, n89941, n89942, n89943, n89944, n89945, n89946,
    n89947, n89948, n89949, n89950, n89952, n89953, n89954, n89955, n89956,
    n89957, n89958, n89959, n89960, n89961, n89962, n89963, n89964, n89965,
    n89966, n89967, n89968, n89969, n89970, n89971, n89972, n89973, n89974,
    n89975, n89976, n89977, n89978, n89979, n89980, n89981, n89982, n89983,
    n89984, n89985, n89986, n89987, n89988, n89989, n89990, n89991, n89992,
    n89993, n89994, n89996, n89997, n89998, n89999, n90000, n90001, n90002,
    n90003, n90004, n90005, n90006, n90007, n90008, n90009, n90010, n90011,
    n90012, n90013, n90014, n90015, n90016, n90017, n90018, n90019, n90020,
    n90021, n90022, n90023, n90024, n90025, n90026, n90027, n90028, n90029,
    n90030, n90031, n90032, n90033, n90034, n90035, n90036, n90037, n90038,
    n90039, n90040, n90041, n90042, n90043, n90044, n90045, n90046, n90047,
    n90048, n90049, n90050, n90051, n90052, n90053, n90054, n90055, n90056,
    n90057, n90058, n90059, n90060, n90061, n90062, n90063, n90064, n90065,
    n90066, n90067, n90068, n90069, n90070, n90071, n90072, n90073, n90074,
    n90075, n90076, n90077, n90078, n90079, n90080, n90081, n90082, n90083,
    n90084, n90085, n90086, n90087, n90088, n90089, n90090, n90091, n90092,
    n90094, n90095, n90096, n90097, n90098, n90099, n90100, n90101, n90102,
    n90103, n90104, n90105, n90106, n90107, n90108, n90109, n90110, n90111,
    n90112, n90113, n90114, n90115, n90116, n90117, n90118, n90119, n90120,
    n90121, n90122, n90123, n90124, n90125, n90126, n90127, n90128, n90129,
    n90130, n90131, n90132, n90133, n90134, n90135, n90136, n90137, n90138,
    n90139, n90140, n90142, n90143, n90144, n90145, n90146, n90147, n90148,
    n90149, n90150, n90151, n90152, n90153, n90154, n90155, n90156, n90157,
    n90158, n90159, n90160, n90161, n90162, n90163, n90164, n90165, n90166,
    n90167, n90168, n90169, n90170, n90171, n90172, n90173, n90174, n90175,
    n90176, n90177, n90178, n90179, n90180, n90181, n90182, n90183, n90184,
    n90185, n90186, n90187, n90188, n90190, n90191, n90192, n90193, n90194,
    n90195, n90196, n90197, n90198, n90199, n90200, n90201, n90202, n90203,
    n90204, n90205, n90206, n90207, n90208, n90209, n90210, n90211, n90212,
    n90213, n90214, n90215, n90216, n90217, n90218, n90219, n90220, n90221,
    n90222, n90223, n90224, n90225, n90226, n90227, n90228, n90229, n90230,
    n90231, n90232, n90233, n90234, n90235, n90236, n90238, n90239, n90240,
    n90241, n90242, n90243, n90244, n90245, n90246, n90247, n90248, n90249,
    n90250, n90251, n90252, n90253, n90254, n90255, n90256, n90257, n90258,
    n90259, n90260, n90261, n90262, n90263, n90264, n90265, n90266, n90267,
    n90268, n90269, n90270, n90271, n90272, n90273, n90274, n90275, n90276,
    n90277, n90278, n90279, n90280, n90281, n90282, n90283, n90284, n90286,
    n90287, n90288, n90289, n90290, n90291, n90292, n90293, n90294, n90295,
    n90296, n90297, n90298, n90299, n90300, n90301, n90302, n90303, n90304,
    n90305, n90306, n90307, n90308, n90309, n90310, n90311, n90312, n90313,
    n90314, n90315, n90316, n90317, n90318, n90319, n90320, n90321, n90322,
    n90323, n90324, n90325, n90326, n90327, n90328, n90329, n90330, n90331,
    n90332, n90334, n90335, n90336, n90337, n90338, n90339, n90340, n90341,
    n90342, n90343, n90344, n90345, n90346, n90347, n90348, n90349, n90350,
    n90351, n90352, n90353, n90354, n90355, n90356, n90357, n90358, n90359,
    n90360, n90361, n90362, n90363, n90364, n90365, n90366, n90367, n90368,
    n90369, n90370, n90371, n90372, n90373, n90374, n90375, n90376, n90377,
    n90378, n90379, n90380, n90382, n90383, n90384, n90385, n90386, n90387,
    n90388, n90389, n90390, n90391, n90392, n90393, n90394, n90395, n90396,
    n90397, n90398, n90399, n90400, n90401, n90402, n90403, n90404, n90405,
    n90406, n90407, n90408, n90409, n90410, n90411, n90412, n90413, n90414,
    n90415, n90416, n90417, n90418, n90419, n90420, n90421, n90422, n90423,
    n90424, n90425, n90426, n90427, n90428, n90430, n90431, n90432, n90433,
    n90434, n90435, n90436, n90437, n90439, n90440, n90441, n90442, n90443,
    n90444, n90445, n90446, n90448, n90449, n90450, n90451, n90452, n90453,
    n90454, n90456, n90457, n90458, n90459, n90460, n90461, n90462, n90463,
    n90465, n90466, n90467, n90468, n90469, n90470, n90471, n90472, n90473,
    n90475, n90476, n90477, n90478, n90479, n90480, n90481, n90482, n90484,
    n90485, n90486, n90487, n90488, n90489, n90490, n90491, n90492, n90494,
    n90495, n90496, n90497, n90498, n90499, n90500, n90501, n90503, n90504,
    n90505, n90506, n90507, n90508, n90509, n90510, n90511, n90513, n90514,
    n90515, n90516, n90517, n90518, n90519, n90520, n90522, n90523, n90524,
    n90525, n90526, n90527, n90528, n90529, n90530, n90532, n90533, n90534,
    n90535, n90536, n90537, n90538, n90539, n90541, n90542, n90543, n90544,
    n90545, n90546, n90547, n90548, n90549, n90551, n90552, n90553, n90554,
    n90555, n90556, n90557, n90558, n90560, n90561, n90562, n90563, n90564,
    n90565, n90566, n90567, n90568, n90570, n90571, n90572, n90573, n90574,
    n90575, n90576, n90577, n90579, n90580, n90581, n90582, n90583, n90584,
    n90585, n90586, n90587, n90589, n90590, n90591, n90592, n90593, n90594,
    n90595, n90596, n90598, n90599, n90600, n90601, n90602, n90603, n90604,
    n90605, n90606, n90608, n90609, n90610, n90611, n90612, n90613, n90614,
    n90615, n90617, n90618, n90619, n90620, n90621, n90622, n90623, n90624,
    n90625, n90627, n90628, n90629, n90630, n90631, n90632, n90633, n90634,
    n90636, n90637, n90638, n90639, n90640, n90641, n90642, n90643, n90644,
    n90646, n90647, n90648, n90649, n90650, n90651, n90652, n90653, n90655,
    n90656, n90657, n90658, n90659, n90660, n90661, n90662, n90663, n90665,
    n90666, n90667, n90668, n90669, n90670, n90671, n90672, n90674, n90675,
    n90676, n90677, n90678, n90679, n90680, n90681, n90682, n90684, n90685,
    n90686, n90687, n90688, n90689, n90690, n90691, n90693, n90694, n90695,
    n90696, n90697, n90698, n90699, n90700, n90701, n90703, n90704, n90705,
    n90706, n90707, n90708, n90709, n90710, n90712, n90713, n90714, n90715,
    n90716, n90717, n90718, n90719, n90720, n90722, n90723, n90724, n90725,
    n90726, n90727, n90728, n90729, n90731, n90732, n90733, n90734, n90735,
    n90736, n90738, n90739, n90740, n90741, n90742, n90743, n90744, n90745,
    n90746, n90747, n90748, n90749, n90750, n90751, n90752, n90753, n90754,
    n90755, n90756, n90757, n90758, n90759, n90760, n90761, n90762, n90763,
    n90764, n90765, n90766, n90767, n90768, n90769, n90770, n90771, n90772,
    n90773, n90774, n90775, n90776, n90777, n90778, n90779, n90781, n90782,
    n90783, n90784, n90785, n90786, n90787, n90788, n90789, n90790, n90791,
    n90792, n90793, n90794, n90795, n90796, n90797, n90798, n90799, n90800,
    n90801, n90802, n90804, n90805, n90806, n90807, n90808, n90809, n90810,
    n90811, n90812, n90813, n90814, n90815, n90816, n90817, n90818, n90819,
    n90820, n90821, n90822, n90823, n90824, n90825, n90826, n90827, n90828,
    n90829, n90830, n90831, n90832, n90834, n90835, n90836, n90837, n90838,
    n90839, n90840, n90841, n90842, n90843, n90844, n90845, n90846, n90847,
    n90848, n90849, n90850, n90851, n90852, n90853, n90854, n90855, n90856,
    n90857, n90858, n90859, n90860, n90861, n90862, n90863, n90865, n90866,
    n90867, n90868, n90869, n90870, n90871, n90872, n90873, n90874, n90875,
    n90876, n90877, n90878, n90879, n90880, n90881, n90882, n90883, n90884,
    n90885, n90886, n90887, n90888, n90889, n90890, n90891, n90892, n90893,
    n90894, n90895, n90896, n90897, n90898, n90899, n90900, n90902, n90903,
    n90904, n90905, n90906, n90907, n90908, n90909, n90910, n90911, n90912,
    n90913, n90914, n90915, n90916, n90917, n90918, n90919, n90920, n90921,
    n90922, n90923, n90924, n90925, n90926, n90927, n90928, n90929, n90930,
    n90931, n90933, n90934, n90935, n90936, n90937, n90938, n90939, n90940,
    n90941, n90942, n90943, n90944, n90945, n90946, n90947, n90948, n90949,
    n90950, n90951, n90952, n90953, n90954, n90955, n90956, n90957, n90958,
    n90959, n90961, n90962, n90963, n90964, n90965, n90966, n90967, n90968,
    n90969, n90970, n90971, n90972, n90973, n90974, n90975, n90976, n90977,
    n90978, n90979, n90980, n90981, n90982, n90983, n90984, n90985, n90987,
    n90988, n90989, n90990, n90991, n90992, n90993, n90994, n90995, n90996,
    n90997, n90998, n90999, n91000, n91001, n91002, n91003, n91004, n91005,
    n91006, n91007, n91008, n91009, n91010, n91011, n91012, n91013, n91015,
    n91016, n91017, n91018, n91019, n91020, n91021, n91022, n91023, n91024,
    n91025, n91026, n91027, n91028, n91029, n91030, n91031, n91032, n91033,
    n91034, n91035, n91036, n91037, n91038, n91039, n91041, n91042, n91043,
    n91044, n91045, n91046, n91047, n91048, n91049, n91050, n91051, n91052,
    n91053, n91054, n91055, n91056, n91057, n91058, n91059, n91060, n91061,
    n91062, n91063, n91064, n91065, n91066, n91067, n91069, n91070, n91071,
    n91072, n91073, n91074, n91075, n91076, n91077, n91078, n91079, n91080,
    n91081, n91082, n91083, n91084, n91085, n91086, n91087, n91088, n91089,
    n91090, n91091, n91092, n91093, n91095, n91096, n91097, n91098, n91099,
    n91100, n91101, n91102, n91103, n91104, n91105, n91106, n91107, n91108,
    n91109, n91110, n91111, n91112, n91113, n91114, n91115, n91116, n91117,
    n91118, n91119, n91120, n91121, n91123, n91124, n91125, n91126, n91127,
    n91128, n91129, n91130, n91131, n91132, n91133, n91134, n91135, n91136,
    n91137, n91138, n91139, n91140, n91141, n91142, n91143, n91144, n91145,
    n91146, n91147, n91149, n91150, n91151, n91152, n91153, n91154, n91155,
    n91156, n91157, n91158, n91159, n91160, n91161, n91162, n91163, n91164,
    n91165, n91166, n91167, n91168, n91169, n91170, n91171, n91172, n91173,
    n91174, n91175, n91177, n91178, n91179, n91180, n91181, n91182, n91183,
    n91184, n91185, n91186, n91187, n91188, n91189, n91190, n91191, n91192,
    n91193, n91194, n91195, n91196, n91197, n91198, n91199, n91200, n91201,
    n91203, n91204, n91205, n91206, n91207, n91208, n91209, n91210, n91211,
    n91212, n91213, n91214, n91215, n91216, n91217, n91218, n91219, n91220,
    n91221, n91222, n91223, n91224, n91225, n91226, n91227, n91228, n91229,
    n91231, n91232, n91233, n91234, n91235, n91236, n91237, n91238, n91239,
    n91240, n91241, n91242, n91243, n91244, n91245, n91246, n91247, n91248,
    n91249, n91250, n91251, n91252, n91253, n91254, n91255, n91257, n91258,
    n91259, n91260, n91261, n91262, n91263, n91264, n91265, n91266, n91267,
    n91268, n91269, n91270, n91271, n91272, n91273, n91274, n91275, n91276,
    n91277, n91278, n91279, n91280, n91281, n91282, n91283, n91285, n91286,
    n91287, n91288, n91289, n91290, n91291, n91292, n91293, n91294, n91295,
    n91296, n91297, n91298, n91299, n91300, n91301, n91302, n91303, n91304,
    n91305, n91306, n91307, n91308, n91309, n91311, n91312, n91313, n91314,
    n91315, n91316, n91317, n91318, n91319, n91320, n91321, n91322, n91323,
    n91324, n91325, n91326, n91327, n91328, n91329, n91330, n91331, n91332,
    n91333, n91334, n91335, n91336, n91338, n91339, n91340, n91341, n91342,
    n91343, n91344, n91345, n91346, n91347, n91348, n91349, n91350, n91351,
    n91352, n91353, n91354, n91355, n91356, n91357, n91358, n91359, n91360,
    n91361, n91363, n91364, n91365, n91366, n91367, n91368, n91369, n91370,
    n91371, n91372, n91373, n91374, n91375, n91376, n91377, n91378, n91379,
    n91380, n91381, n91382, n91383, n91384, n91385, n91386, n91387, n91388,
    n91390, n91391, n91392, n91393, n91394, n91395, n91396, n91397, n91398,
    n91399, n91400, n91401, n91402, n91403, n91404, n91405, n91406, n91407,
    n91408, n91409, n91410, n91411, n91412, n91413, n91415, n91416, n91417,
    n91418, n91419, n91420, n91421, n91422, n91423, n91424, n91425, n91426,
    n91427, n91428, n91429, n91430, n91431, n91432, n91433, n91434, n91435,
    n91436, n91437, n91438, n91439, n91440, n91442, n91443, n91444, n91445,
    n91446, n91447, n91448, n91449, n91450, n91451, n91452, n91453, n91454,
    n91455, n91456, n91457, n91458, n91459, n91460, n91461, n91462, n91463,
    n91464, n91465, n91467, n91468, n91469, n91470, n91471, n91472, n91473,
    n91474, n91475, n91476, n91477, n91478, n91479, n91480, n91481, n91482,
    n91483, n91484, n91485, n91486, n91487, n91488, n91489, n91490, n91491,
    n91492, n91494, n91495, n91496, n91497, n91498, n91499, n91500, n91501,
    n91502, n91503, n91504, n91505, n91506, n91507, n91508, n91509, n91510,
    n91511, n91512, n91513, n91514, n91515, n91516, n91517, n91519, n91520,
    n91521, n91522, n91523, n91524, n91525, n91526, n91527, n91528, n91529,
    n91530, n91531, n91532, n91533, n91534, n91535, n91536, n91537, n91538,
    n91539, n91540, n91541, n91542, n91543, n91544, n91546, n91547, n91548,
    n91549, n91550, n91551, n91552, n91553, n91554, n91555, n91556, n91557,
    n91558, n91559, n91560, n91561, n91562, n91563, n91564, n91565, n91566,
    n91567, n91568, n91569, n91571, n91572, n91573, n91574, n91575, n91576,
    n91577, n91578, n91579, n91580, n91581, n91582, n91583, n91584, n91585,
    n91586, n91587, n91588, n91589, n91590, n91591, n91592, n91593, n91594,
    n91596, n91597, n91598, n91599, n91600, n91601, n91602, n91603, n91604,
    n91605, n91606, n91607, n91608, n91609, n91610, n91611, n91612, n91613,
    n91614, n91615, n91616, n91617, n91618, n91619, n91621, n91622, n91623,
    n91624, n91625, n91626, n91627, n91628, n91629, n91630, n91631, n91632,
    n91633, n91634, n91635, n91636, n91637, n91638, n91639, n91640, n91641,
    n91642, n91643, n91644, n91645, n91646, n91647, n91648, n91649, n91650,
    n91651, n91652, n91653, n91654, n91655, n91656, n91657, n91658, n91660,
    n91661, n91662, n91663, n91664, n91665, n91666, n91667, n91669, n91670,
    n91671, n91673, n91674, n91675, n91677, n91678, n91680, n91681, n91682,
    n91684, n91685, n91687, n91688, n91689, n91690, n91692, n91693, n91694,
    n91695, n91696, n91697, n91698, n91699, n91700, n91701, n91702, n91703,
    n91704, n91705, n91706, n91708, n91709, n91710, n91712, n91713, n91715,
    n91716, n91717, n91719, n91721, n91722, n91723, n91724, n91725, n91727,
    n91728, n91729, n121, n126, n131, n136, n141, n146, n151, n156, n161,
    n166, n171, n176, n181, n186, n191, n196, n201, n206, n211, n216, n221,
    n226, n231, n236, n241, n246, n251, n256, n261, n266, n271, n276, n281,
    n286, n291, n296, n301, n306, n311, n316, n321, n326, n331, n336, n341,
    n346, n351, n356, n361, n366, n371, n376, n381, n386, n391, n396, n401,
    n406, n411, n416, n421, n426, n431, n436, n441, n446, n451, n456, n461,
    n466, n471, n476, n481, n486, n491, n496, n501, n506, n511, n516, n521,
    n526, n531, n536, n541, n546, n551, n556, n561, n566, n571, n576, n581,
    n586, n591, n596, n601, n606, n611, n616, n621, n626, n631, n636, n641,
    n646, n651, n656, n661, n666, n671, n676, n681, n686, n691, n696, n701,
    n706, n711, n716, n721, n726, n731, n736, n741, n746, n751, n756, n761,
    n766, n771, n776, n781, n786, n791, n796, n801, n806, n811, n816, n821,
    n826, n831, n836, n841, n846, n851, n856, n861, n866, n871, n876, n881,
    n886, n891, n896, n901, n906, n911, n916, n921, n926, n931, n936, n941,
    n946, n951, n956, n961, n966, n971, n976, n981, n986, n991, n996,
    n1001, n1006, n1011, n1016, n1021, n1026, n1031, n1036, n1041, n1046,
    n1051, n1056, n1061, n1066, n1071, n1076, n1081, n1086, n1091, n1096,
    n1101, n1106, n1111, n1116, n1121, n1126, n1131, n1136, n1141, n1146,
    n1151, n1156, n1161, n1166, n1171, n1176, n1181, n1186, n1191, n1196,
    n1201, n1206, n1211, n1216, n1221, n1226, n1231, n1236, n1241, n1246,
    n1251, n1256, n1261, n1266, n1271, n1276, n1281, n1286, n1291, n1296,
    n1301, n1306, n1311, n1316, n1321, n1326, n1331, n1336, n1341, n1346,
    n1351, n1356, n1361, n1366, n1371, n1376, n1381, n1386, n1391, n1396,
    n1401, n1406, n1411, n1416, n1421, n1426, n1431, n1436, n1441, n1446,
    n1451, n1456, n1461, n1466, n1471, n1476, n1481, n1486, n1491, n1496,
    n1501, n1506, n1511, n1516, n1521, n1526, n1531, n1536, n1541, n1546,
    n1551, n1556, n1561, n1566, n1571, n1576, n1581, n1586, n1591, n1596,
    n1601, n1606, n1611, n1616, n1621, n1626, n1631, n1636, n1641, n1646,
    n1651, n1656, n1661, n1666, n1671, n1676, n1681, n1686, n1691, n1696,
    n1701, n1706, n1711, n1716, n1721, n1726, n1731, n1736, n1741, n1746,
    n1751, n1756, n1761, n1766, n1771, n1776, n1781, n1786, n1791, n1796,
    n1801, n1806, n1811, n1816, n1821, n1826, n1831, n1836, n1841, n1846,
    n1851, n1856, n1861, n1866, n1871, n1876, n1881, n1886, n1891, n1896,
    n1901, n1906, n1911, n1916, n1921, n1926, n1931, n1936, n1941, n1946,
    n1951, n1956, n1961, n1966, n1971, n1976, n1981, n1986, n1991, n1996,
    n2001, n2006, n2011, n2016, n2021, n2026, n2031, n2036, n2041, n2046,
    n2051, n2056, n2061, n2066, n2071, n2076, n2081, n2086, n2091, n2096,
    n2101, n2106, n2111, n2116, n2121, n2126, n2131, n2136, n2141, n2146,
    n2151, n2156, n2161, n2166, n2171, n2176, n2181, n2186, n2191, n2196,
    n2201, n2206, n2211, n2216, n2221, n2226, n2231, n2236, n2241, n2246,
    n2251, n2256, n2261, n2266, n2271, n2276, n2281, n2286, n2291, n2296,
    n2301, n2306, n2311, n2316, n2321, n2326, n2331, n2336, n2341, n2346,
    n2351, n2356, n2361, n2366, n2371, n2376, n2381, n2386, n2391, n2396,
    n2401, n2406, n2411, n2416, n2421, n2426, n2431, n2436, n2441, n2446,
    n2451, n2456, n2461, n2466, n2471, n2476, n2481, n2486, n2491, n2496,
    n2501, n2506, n2511, n2516, n2521, n2526, n2531, n2536, n2541, n2546,
    n2551, n2556, n2561, n2566, n2571, n2576, n2581, n2586, n2591, n2596,
    n2601, n2606, n2611, n2616, n2621, n2626, n2631, n2636, n2641, n2646,
    n2651, n2656, n2661, n2666, n2671, n2676, n2681, n2686, n2691, n2696,
    n2701, n2706, n2711, n2716, n2721, n2726, n2731, n2736, n2741, n2746,
    n2751, n2756, n2761, n2766, n2771, n2776, n2781, n2786, n2791, n2796,
    n2801, n2806, n2811, n2816, n2821, n2826, n2831, n2836, n2841, n2846,
    n2851, n2856, n2861, n2866, n2871, n2876, n2881, n2886, n2891, n2896,
    n2901, n2906, n2911, n2916, n2921, n2926, n2931, n2936, n2941, n2946,
    n2951, n2956, n2961, n2966, n2971, n2976, n2981, n2986, n2991, n2996,
    n3001, n3006, n3011, n3016, n3021, n3026, n3031, n3036, n3041, n3046,
    n3051, n3056, n3061, n3066, n3071, n3076, n3081, n3086, n3091, n3096,
    n3101, n3106, n3111, n3116, n3121, n3126, n3131, n3136, n3141, n3146,
    n3151, n3156, n3161, n3166, n3171, n3176, n3181, n3186, n3191, n3196,
    n3201, n3206, n3211, n3216, n3221, n3226, n3231, n3236, n3241, n3246,
    n3251, n3256, n3261, n3266, n3271, n3276, n3281, n3286, n3291, n3296,
    n3301, n3306, n3311, n3316, n3321, n3326, n3331, n3336, n3341, n3346,
    n3351, n3356, n3361, n3366, n3371, n3376, n3381, n3386, n3391, n3396,
    n3401, n3406, n3411, n3416, n3421, n3426, n3431, n3436, n3441, n3446,
    n3451, n3456, n3461, n3466, n3471, n3476, n3481, n3486, n3491, n3496,
    n3501, n3506, n3511, n3516, n3521, n3526, n3531, n3536, n3541, n3546,
    n3551, n3556, n3561, n3566, n3571, n3576, n3581, n3586, n3591, n3596,
    n3601, n3606, n3611, n3616, n3621, n3626, n3631, n3636, n3641, n3646,
    n3651, n3656, n3661, n3666, n3671, n3676, n3681, n3686, n3691, n3696,
    n3701, n3706, n3711, n3716, n3721, n3726, n3731, n3736, n3741, n3746,
    n3751, n3756, n3761, n3766, n3771, n3776, n3781, n3786, n3791, n3796,
    n3801, n3806, n3811, n3816, n3821, n3826, n3831, n3836, n3841, n3846,
    n3851, n3856, n3861, n3866, n3871, n3876, n3881, n3886, n3891, n3896,
    n3901, n3906, n3911, n3916, n3921, n3926, n3931, n3936, n3941, n3946,
    n3951, n3956, n3961, n3966, n3971, n3976, n3981, n3986, n3991, n3996,
    n4001, n4006, n4011, n4016, n4021, n4026, n4031, n4036, n4041, n4046,
    n4051, n4056, n4061, n4066, n4071, n4076, n4081, n4086, n4091, n4096,
    n4101, n4106, n4111, n4116, n4121, n4126, n4131, n4136, n4141, n4146,
    n4151, n4156, n4161, n4166, n4171, n4176, n4181, n4186, n4191, n4196,
    n4201, n4206, n4211, n4216, n4221, n4226, n4231, n4236, n4241, n4246,
    n4251, n4256, n4261, n4266, n4271, n4276, n4281, n4286, n4291, n4296,
    n4301, n4306, n4311, n4316, n4321, n4326, n4331, n4336, n4341, n4346,
    n4351, n4356, n4361, n4366, n4371, n4376, n4381, n4386, n4391, n4396,
    n4401, n4406, n4411, n4416, n4421, n4426, n4431, n4436, n4441, n4446,
    n4451, n4456, n4461, n4466, n4471, n4476, n4481, n4486, n4491, n4496,
    n4501, n4506, n4511, n4516, n4521, n4526, n4531, n4536, n4541, n4546,
    n4551, n4556, n4561, n4566, n4571, n4576, n4581, n4586, n4591, n4596,
    n4601, n4606, n4611, n4616, n4621, n4626, n4631, n4636, n4641, n4646,
    n4651, n4656, n4661, n4666, n4671, n4676, n4681, n4686, n4691, n4696,
    n4701, n4706, n4711, n4716, n4721, n4726, n4731, n4736, n4741, n4746,
    n4751, n4756, n4761, n4766, n4771, n4776, n4781, n4786, n4791, n4796,
    n4801, n4806, n4811, n4816, n4821, n4826, n4831, n4836, n4841, n4846,
    n4851, n4856, n4861, n4866, n4871, n4876, n4881, n4886, n4891, n4896,
    n4901, n4906, n4911, n4916, n4921, n4926, n4931, n4936, n4941, n4946,
    n4951, n4956, n4961, n4966, n4971, n4976, n4981, n4986, n4991, n4996,
    n5001, n5006, n5011, n5016, n5021, n5026, n5031, n5036, n5041, n5046,
    n5051, n5056, n5061, n5066, n5071, n5076, n5081, n5086, n5091, n5096,
    n5101, n5106, n5111, n5116, n5121, n5126, n5131, n5136, n5141, n5146,
    n5151, n5156, n5161, n5166, n5171, n5176, n5181, n5186, n5191, n5196,
    n5201, n5206, n5211, n5216, n5221, n5226, n5231, n5236, n5241, n5246,
    n5251, n5256, n5261, n5266, n5271, n5276, n5281, n5286, n5291, n5296,
    n5301, n5306, n5311, n5316, n5321, n5326, n5331, n5336, n5341, n5346,
    n5351, n5356, n5361, n5366, n5371, n5376, n5381, n5386, n5391, n5396,
    n5401, n5406, n5411, n5416, n5421, n5426, n5431, n5436, n5441, n5446,
    n5451, n5456, n5461, n5466, n5471, n5476, n5481, n5486, n5491, n5496,
    n5501, n5506, n5511, n5516, n5521, n5526, n5531, n5536, n5541, n5546,
    n5551, n5556, n5561, n5566, n5571, n5576, n5581, n5586, n5591, n5596,
    n5601, n5606, n5611, n5616, n5621, n5626, n5631, n5636, n5641, n5646,
    n5651, n5656, n5661, n5666, n5671, n5676, n5681, n5686, n5691, n5696,
    n5701, n5706, n5711, n5716, n5721, n5726, n5731, n5736, n5741, n5746,
    n5751, n5756, n5761, n5766, n5771, n5776, n5781, n5786, n5791, n5796,
    n5801, n5806, n5811, n5816, n5821, n5826, n5831, n5836, n5841, n5846,
    n5851, n5856, n5861, n5866, n5871, n5876, n5881, n5886, n5891, n5896,
    n5901, n5906, n5911, n5916, n5921, n5926, n5931, n5936, n5941, n5946,
    n5951, n5956, n5961, n5966, n5971, n5976, n5981, n5986, n5991, n5996,
    n6001, n6006, n6011, n6016, n6021, n6026, n6031, n6036, n6041, n6046,
    n6051, n6056, n6061, n6066, n6071, n6076, n6081, n6086, n6091, n6096,
    n6101, n6106, n6111, n6116, n6121, n6126, n6131, n6136, n6141, n6146,
    n6151, n6156, n6161, n6166, n6171, n6176, n6181, n6186, n6191, n6196,
    n6201, n6206, n6211, n6216, n6221, n6226, n6231, n6236, n6241, n6246,
    n6251, n6256, n6261, n6266, n6271, n6276, n6281, n6286, n6291, n6296,
    n6301, n6306, n6311, n6316, n6321, n6326, n6331, n6336, n6341, n6346,
    n6351, n6356, n6361, n6366, n6371, n6376, n6381, n6386, n6391, n6396,
    n6401, n6406, n6411, n6416, n6421, n6426, n6431, n6436, n6441, n6446,
    n6451, n6456, n6461, n6466, n6471, n6476, n6481, n6486, n6491, n6496,
    n6501, n6506, n6511, n6516, n6521, n6526, n6531, n6536, n6541, n6546,
    n6551, n6556, n6561, n6566, n6571, n6576, n6581, n6586, n6591, n6596,
    n6601, n6606, n6611, n6616, n6621, n6626, n6631, n6636, n6641, n6646,
    n6651, n6656, n6661, n6666, n6671, n6676, n6681, n6686, n6691, n6696,
    n6701, n6706, n6711, n6716, n6721, n6726, n6731, n6736, n6741, n6746,
    n6751, n6756, n6761, n6766, n6771, n6776, n6781, n6786, n6791, n6796,
    n6801, n6806, n6811, n6816, n6821, n6826, n6831, n6836, n6841, n6846,
    n6851, n6856, n6861, n6866, n6871, n6876, n6881, n6886, n6891, n6896,
    n6901, n6906, n6911, n6916, n6921, n6926, n6931, n6936, n6941, n6946,
    n6951, n6956, n6961, n6966, n6971, n6976, n6981, n6986, n6991, n6996,
    n7001, n7006, n7011, n7016, n7021, n7026, n7031, n7036, n7041, n7046,
    n7051, n7056, n7061, n7066, n7071, n7076, n7081, n7086, n7091, n7096,
    n7101, n7106, n7111, n7116, n7121, n7126, n7131, n7136, n7141, n7146,
    n7151, n7156, n7161, n7166, n7171, n7176, n7181, n7186, n7191, n7196,
    n7201, n7206, n7211, n7216, n7221, n7226, n7231, n7236, n7241, n7246,
    n7251, n7256, n7261, n7266, n7271, n7276, n7281, n7286, n7291, n7296,
    n7301, n7306, n7311, n7316, n7321, n7326, n7331, n7336, n7341, n7346,
    n7351, n7356, n7361, n7366, n7371, n7376, n7381, n7386, n7391, n7396,
    n7401, n7406, n7411, n7416, n7421, n7426, n7431, n7436, n7441, n7446,
    n7451, n7456, n7461, n7466, n7471, n7476, n7481, n7486, n7491, n7496,
    n7501, n7506, n7511, n7516, n7521, n7526, n7531, n7536, n7541, n7546,
    n7551, n7556, n7561, n7566, n7571, n7576, n7581, n7586, n7591, n7596,
    n7601, n7606, n7611, n7616, n7621, n7626, n7631, n7636, n7641, n7646,
    n7651, n7656, n7661, n7666, n7671, n7676, n7681, n7686, n7691, n7696,
    n7701, n7706, n7711, n7716, n7721, n7726, n7731, n7736, n7741, n7746,
    n7751, n7756, n7761, n7766, n7771, n7776, n7781, n7786, n7791, n7796,
    n7801, n7806, n7811, n7816, n7821, n7826, n7831, n7836, n7841, n7846,
    n7851, n7856, n7861, n7866, n7871, n7876, n7881, n7886, n7891, n7896,
    n7901, n7906, n7911, n7916, n7921, n7926, n7931, n7936, n7941, n7946,
    n7951, n7956, n7961, n7966, n7971, n7976, n7981, n7986, n7991, n7996,
    n8001, n8006, n8011, n8016, n8021, n8026, n8031, n8036, n8041, n8046,
    n8051, n8056, n8061, n8066, n8071, n8076, n8081, n8086, n8091, n8096,
    n8101, n8106, n8111, n8116, n8121, n8126, n8131, n8136, n8141, n8146,
    n8151, n8156, n8161, n8166, n8171, n8176, n8181, n8186, n8191, n8196,
    n8201, n8206, n8211, n8216, n8221, n8226, n8231, n8236, n8241, n8246,
    n8251, n8256, n8261, n8266, n8271, n8276, n8281, n8286, n8291, n8296,
    n8301, n8306, n8311, n8316, n8321, n8326, n8331, n8336, n8341, n8346,
    n8351, n8356, n8361, n8366, n8371, n8376, n8381, n8386, n8391, n8396,
    n8401, n8406, n8411, n8416, n8421, n8426, n8431, n8436, n8441, n8446,
    n8451, n8456, n8461, n8466, n8471, n8476, n8481, n8486, n8491, n8496,
    n8501, n8506, n8511, n8516, n8521, n8526, n8531, n8536, n8541, n8546,
    n8551, n8556, n8561, n8566, n8571, n8576, n8581, n8586, n8591, n8596,
    n8601, n8606, n8611, n8616, n8621, n8626, n8631, n8636, n8641, n8646,
    n8651, n8656, n8661, n8666, n8671, n8676, n8681, n8686, n8691, n8696,
    n8701, n8706, n8711, n8716, n8721, n8726, n8731, n8736, n8741, n8746,
    n8751, n8756, n8761, n8766, n8771, n8776, n8781, n8786, n8791, n8796,
    n8801, n8806, n8811, n8816, n8821, n8826, n8831, n8836, n8841, n8846,
    n8851, n8856, n8861, n8866, n8871, n8876, n8881, n8886, n8891, n8896,
    n8901, n8906, n8911, n8916, n8921, n8926, n8931, n8936, n8941, n8946,
    n8951, n8956, n8961, n8966, n8971, n8976, n8981, n8986, n8991, n8996,
    n9001, n9006, n9011, n9016, n9021, n9026, n9031, n9036, n9041, n9046,
    n9051, n9056, n9061, n9066, n9071, n9076, n9081, n9086, n9091, n9096,
    n9101, n9106, n9111, n9116, n9121, n9126, n9131, n9136, n9141, n9146,
    n9151, n9156, n9161, n9166, n9171, n9176, n9181, n9186, n9191, n9196,
    n9201, n9206, n9211, n9216, n9221, n9226, n9231, n9236, n9241, n9246,
    n9251, n9256, n9261, n9266, n9271, n9276, n9281, n9286, n9291, n9296,
    n9301, n9306, n9311, n9316, n9321, n9326, n9331, n9336, n9341, n9346,
    n9351, n9356, n9361, n9366, n9371, n9376, n9381, n9386, n9391, n9396,
    n9401, n9406, n9411, n9416, n9421, n9426, n9431, n9436, n9441, n9446,
    n9451, n9456, n9461, n9466, n9471, n9476, n9481, n9486, n9491, n9496,
    n9501, n9506, n9511, n9516, n9521, n9526, n9531, n9536, n9541, n9546,
    n9551, n9556, n9561, n9566, n9571, n9576, n9581, n9586, n9591, n9596,
    n9601, n9606, n9611, n9616, n9621, n9626, n9631, n9636, n9641, n9646,
    n9651, n9656, n9661, n9666, n9671, n9676, n9681, n9686, n9691, n9696,
    n9701, n9706, n9711, n9716, n9721, n9726, n9731, n9736, n9741, n9746,
    n9751, n9756, n9761, n9766, n9771, n9776, n9781, n9786, n9791, n9796,
    n9801, n9806, n9811, n9816, n9821, n9826, n9831, n9836, n9841, n9846,
    n9851, n9856, n9861, n9866, n9871, n9876, n9881, n9886, n9891, n9896,
    n9901, n9906, n9911, n9916, n9921, n9926, n9931, n9936, n9941, n9946,
    n9951, n9956, n9961, n9966, n9971, n9976, n9981, n9986, n9991, n9996,
    n10001, n10006, n10011, n10016, n10021, n10026, n10031, n10036, n10041,
    n10046, n10051, n10056, n10061, n10066, n10071, n10076, n10081, n10086,
    n10091, n10096, n10101, n10106, n10111, n10116, n10121, n10126, n10131,
    n10136, n10141, n10146, n10151, n10156, n10161, n10166, n10171, n10176,
    n10181, n10186, n10191, n10196, n10201, n10206, n10211, n10216, n10221,
    n10226, n10231, n10236, n10241, n10246, n10251, n10256, n10261, n10266,
    n10271, n10276, n10281, n10286, n10291, n10296, n10301, n10306, n10311,
    n10316, n10321, n10326, n10331, n10336, n10341, n10346, n10351, n10356,
    n10361, n10366, n10371, n10376, n10381, n10386, n10391, n10396, n10401,
    n10406, n10411, n10416, n10421, n10426, n10431, n10436, n10441, n10446,
    n10451, n10456, n10461, n10466, n10471, n10476, n10481, n10486, n10491,
    n10496, n10501, n10506, n10511, n10516, n10521, n10526, n10531, n10536,
    n10541, n10546, n10551, n10556, n10561, n10566, n10571, n10576, n10581,
    n10586, n10591, n10596, n10601, n10606, n10611, n10616, n10621, n10626,
    n10631, n10636, n10641, n10646, n10651, n10656, n10661, n10666, n10671,
    n10676, n10681, n10686, n10691, n10696, n10701, n10706, n10711, n10716,
    n10721, n10726, n10731, n10736, n10741, n10746, n10751, n10756, n10761,
    n10766, n10771, n10776, n10781, n10786, n10791, n10796, n10801, n10806,
    n10811, n10816, n10821, n10826, n10831, n10836, n10841, n10846, n10851,
    n10856, n10861, n10866, n10871, n10876, n10881, n10886, n10891, n10896,
    n10901, n10906, n10911, n10916, n10921, n10926, n10931, n10936, n10941,
    n10946, n10951, n10956, n10961, n10966, n10971, n10976, n10981, n10986,
    n10991, n10996, n11001, n11006, n11011, n11016, n11021, n11026, n11031,
    n11036, n11041, n11046, n11051, n11056, n11061, n11066, n11071, n11076,
    n11081, n11086, n11091, n11096, n11101, n11106, n11111, n11116, n11121,
    n11126, n11131, n11136, n11141, n11146, n11151, n11156, n11161, n11166,
    n11171, n11176, n11181, n11186, n11191, n11196, n11201, n11206, n11211,
    n11216, n11221, n11226, n11231, n11236, n11241, n11246, n11251, n11256,
    n11261, n11266, n11271, n11276, n11281, n11286, n11291, n11296, n11301,
    n11306, n11311, n11316, n11321, n11326, n11331, n11336, n11341, n11346,
    n11351, n11356, n11361, n11366, n11371, n11376, n11381, n11386, n11391,
    n11396, n11401, n11406, n11411, n11416, n11421, n11426, n11431, n11436,
    n11441, n11446, n11451, n11456, n11461, n11466, n11471, n11476, n11481,
    n11486, n11491, n11496, n11501, n11506, n11511, n11516, n11521, n11526,
    n11531, n11536, n11541, n11546, n11551, n11556, n11561, n11566, n11571,
    n11576, n11581, n11586, n11591, n11596, n11601, n11606, n11611, n11616,
    n11621, n11626, n11631, n11636, n11641, n11646, n11651, n11656, n11661,
    n11666, n11671, n11676, n11681, n11686, n11691, n11696, n11701, n11706,
    n11711, n11716, n11721, n11726, n11731, n11736, n11741, n11746, n11751,
    n11756, n11761, n11766, n11771, n11776, n11781, n11786, n11791, n11796,
    n11801, n11806, n11811, n11816, n11821, n11826, n11831, n11836, n11841,
    n11846, n11851, n11856, n11861, n11866, n11871, n11876, n11881, n11886,
    n11891, n11896, n11901, n11906, n11911, n11916, n11921, n11926, n11931,
    n11936, n11941, n11946, n11951, n11956, n11961, n11966, n11971, n11976,
    n11981, n11986, n11991, n11996, n12001, n12006, n12011, n12016, n12021,
    n12026, n12031, n12036, n12041, n12046, n12051, n12056, n12061, n12066,
    n12071, n12076, n12081, n12086, n12091, n12096, n12101, n12106, n12111,
    n12116, n12121, n12126, n12131, n12136, n12141, n12146, n12151, n12156,
    n12161, n12166, n12171, n12176, n12181, n12186, n12191, n12196, n12201,
    n12206, n12211, n12216, n12221, n12226, n12231, n12236, n12241, n12246,
    n12251, n12256, n12261, n12266, n12271, n12276, n12281, n12286, n12291,
    n12296, n12301, n12306, n12311, n12316, n12321, n12326, n12331, n12336,
    n12341, n12346, n12351, n12356, n12361, n12366, n12371, n12376, n12381,
    n12386, n12391, n12396, n12401, n12406, n12411, n12416, n12421, n12426,
    n12431, n12436, n12441, n12446, n12451, n12456, n12461, n12466, n12471,
    n12476, n12481, n12486, n12491, n12496, n12501, n12506, n12511, n12516,
    n12521, n12526, n12531, n12536, n12541, n12546, n12551, n12556, n12561,
    n12566, n12571, n12576, n12581, n12586, n12591, n12596, n12601, n12606,
    n12611, n12616, n12621, n12626, n12631, n12636, n12641, n12646, n12651,
    n12656, n12661, n12666, n12671, n12676, n12681, n12686, n12691, n12696,
    n12701, n12706, n12711, n12716, n12721, n12726, n12731, n12736, n12741,
    n12746, n12751, n12756, n12761, n12766, n12771, n12776, n12781, n12786,
    n12791, n12796, n12801, n12806, n12811, n12816, n12821, n12826, n12831,
    n12836, n12841, n12846, n12851, n12856, n12861, n12866, n12871, n12876,
    n12881, n12886, n12891, n12896, n12901, n12906, n12911, n12916, n12921,
    n12926, n12931, n12936, n12941, n12946, n12951, n12956, n12961, n12966,
    n12971, n12976, n12981, n12986, n12991, n12996, n13001, n13006, n13011,
    n13016, n13021, n13026, n13031, n13036, n13041, n13046, n13051, n13056,
    n13061, n13066, n13071, n13076, n13081, n13086, n13091, n13096, n13101,
    n13106, n13111, n13116, n13121, n13126, n13131, n13136, n13141, n13146,
    n13151, n13156, n13161, n13166, n13171, n13176, n13181, n13186, n13191,
    n13196, n13201, n13206, n13211, n13216, n13221, n13226, n13231, n13236,
    n13241, n13246, n13251, n13256, n13261, n13266, n13271, n13276, n13281,
    n13286, n13291, n13296, n13301, n13306, n13311, n13316, n13321, n13326,
    n13331, n13336, n13341, n13346, n13351, n13356, n13361, n13366, n13371,
    n13376, n13381, n13386, n13391, n13396, n13401, n13406, n13411, n13416,
    n13421, n13426, n13431, n13436, n13441, n13446, n13451, n13456, n13461,
    n13466, n13471, n13476, n13481, n13486, n13491, n13496, n13501, n13506,
    n13511, n13516, n13521, n13526, n13531, n13536, n13541, n13546, n13551,
    n13556, n13561, n13566, n13571, n13576, n13581, n13586, n13591, n13596,
    n13601, n13606, n13611, n13616, n13621, n13626, n13631, n13636, n13641,
    n13646, n13651, n13656, n13661, n13666, n13671, n13676, n13681, n13686,
    n13691, n13696, n13701, n13706, n13711, n13716, n13721, n13726, n13731,
    n13736, n13741, n13746, n13751, n13756, n13761, n13766, n13771, n13776,
    n13781, n13786, n13791, n13796, n13801, n13806, n13811, n13816, n13821,
    n13826, n13831, n13836, n13841, n13846, n13851, n13856, n13861, n13866,
    n13871, n13876, n13881, n13886, n13891, n13896, n13901, n13906, n13911,
    n13916, n13921, n13926, n13931, n13936, n13941, n13946, n13951, n13956,
    n13961, n13966, n13971, n13976, n13981, n13986, n13991, n13996, n14001,
    n14006, n14011, n14016, n14021, n14026, n14031, n14036, n14041, n14046,
    n14051, n14056, n14061, n14066, n14071, n14076, n14081, n14086, n14091,
    n14096, n14101, n14106, n14111, n14116, n14121, n14126, n14131, n14136,
    n14141, n14146, n14151, n14156, n14161, n14166, n14171, n14176, n14181,
    n14186, n14191, n14196, n14201, n14206, n14211, n14216, n14221, n14226,
    n14231, n14236, n14241, n14246, n14251, n14256, n14261, n14266, n14271,
    n14276, n14281, n14286, n14291, n14296, n14301, n14306, n14311, n14316,
    n14321, n14326, n14331, n14336, n14341, n14346, n14351, n14356, n14361,
    n14366, n14371, n14376, n14381, n14386, n14391, n14396, n14401, n14406,
    n14411, n14416, n14421, n14426, n14431, n14436, n14441, n14446, n14451,
    n14456, n14461, n14466, n14471, n14476, n14481, n14486, n14491, n14496,
    n14501, n14506, n14511, n14516, n14521, n14526, n14531, n14536, n14541,
    n14546, n14551, n14556, n14561, n14566, n14571, n14576, n14581, n14586,
    n14591, n14596, n14601, n14606, n14611, n14616, n14621, n14626, n14631,
    n14636, n14641, n14646, n14651, n14656, n14661, n14666, n14671, n14676,
    n14681, n14686, n14691, n14696, n14701, n14706, n14711, n14716, n14721,
    n14726, n14731, n14736, n14741, n14746, n14751, n14756, n14761, n14766,
    n14771, n14776, n14781, n14786, n14791, n14796, n14801, n14806, n14811,
    n14816, n14821, n14826, n14831, n14836, n14841, n14846, n14851, n14856,
    n14861, n14866, n14871, n14876, n14881, n14886, n14891, n14896, n14901,
    n14906, n14911, n14916, n14921, n14926, n14931, n14936, n14941, n14946,
    n14951, n14956, n14961, n14966, n14971, n14976, n14981, n14986, n14991,
    n14996, n15001, n15006, n15011, n15016, n15021, n15026, n15031, n15036,
    n15041, n15046, n15051, n15056, n15061, n15066, n15071, n15076, n15081,
    n15086, n15091, n15096, n15101, n15106, n15111, n15116, n15121, n15126,
    n15131, n15136, n15141, n15146, n15151, n15156, n15161, n15166, n15171,
    n15176, n15181, n15186, n15191, n15196, n15201, n15206, n15211, n15216,
    n15221, n15226, n15231, n15236, n15241, n15246, n15251, n15256, n15261,
    n15266, n15271, n15276, n15281, n15286, n15291, n15296, n15301, n15306,
    n15311, n15316, n15321, n15326, n15331, n15336, n15341, n15346, n15351,
    n15356, n15361, n15366, n15371, n15376, n15381, n15386, n15391, n15396,
    n15401, n15406, n15411, n15416, n15421, n15426, n15431, n15436, n15441,
    n15446, n15451, n15456, n15461, n15466, n15471, n15476, n15481, n15486,
    n15491, n15496, n15501, n15506, n15511, n15516, n15521, n15526, n15531,
    n15536, n15541, n15546, n15551, n15556, n15561, n15566, n15571, n15576,
    n15581, n15586, n15591, n15596, n15601, n15606, n15611, n15616, n15621,
    n15626, n15631, n15636, n15641, n15646, n15651, n15656, n15661, n15666,
    n15671, n15676, n15681, n15686, n15691, n15696, n15701, n15706, n15711,
    n15716, n15721, n15726, n15731, n15736, n15741, n15746, n15751, n15756,
    n15761, n15766, n15771, n15776, n15781, n15786, n15791, n15796, n15801,
    n15806, n15811, n15816, n15821, n15826, n15831, n15836, n15841, n15846,
    n15851, n15856, n15861, n15866, n15871, n15876, n15881, n15886, n15891,
    n15896, n15901, n15906, n15911, n15916, n15921, n15926, n15931, n15936,
    n15941, n15946, n15951, n15956, n15961, n15966, n15971, n15976, n15981,
    n15986, n15991, n15996, n16001, n16006, n16011, n16016, n16021, n16026,
    n16031, n16036, n16041, n16046, n16051, n16056, n16061, n16066, n16071,
    n16076, n16081, n16086, n16091, n16096, n16101, n16106, n16111, n16116,
    n16121, n16126, n16131, n16136, n16141, n16146, n16151, n16156, n16161,
    n16166, n16171, n16176, n16181, n16186, n16191, n16196, n16201, n16206,
    n16211, n16216, n16221, n16226, n16231, n16236, n16241, n16246, n16251,
    n16256, n16261, n16266, n16271, n16276, n16281, n16286, n16291, n16296,
    n16301, n16306, n16311, n16316, n16321, n16326, n16331, n16336, n16341,
    n16346, n16351, n16356, n16361, n16366, n16371, n16376, n16381, n16386,
    n16391, n16396, n16401, n16406, n16411, n16416, n16421, n16426, n16431,
    n16436, n16441, n16446, n16451, n16456, n16461, n16466, n16471, n16476,
    n16481, n16486, n16491, n16496, n16501, n16506, n16511, n16516, n16521,
    n16526, n16531, n16536, n16541, n16546, n16551, n16556, n16561, n16566,
    n16571, n16576, n16581, n16586, n16591, n16596, n16601, n16606, n16611,
    n16616, n16621, n16626, n16631, n16636, n16641, n16646, n16651, n16656,
    n16661, n16666, n16671, n16676, n16681, n16686, n16691, n16696, n16701,
    n16706, n16711, n16716;
  assign n10021_1 = P3_ADDR_REG_13_ & P3_WR_REG;
  assign n10022 = P2_P3_DATAO_REG_30_ & ~P2_P3_DATAO_REG_31_;
  assign n10023 = P2_P1_DATAO_REG_30_ & ~P2_P1_DATAO_REG_31_;
  assign n10024 = P2_P2_DATAO_REG_30_ & ~P2_P2_DATAO_REG_31_;
  assign n10025 = ~n10022 & ~n10023;
  assign n10026_1 = ~n10024 & n10025;
  assign n10027 = P2_P3_ADDRESS_REG_13_ & n10026_1;
  assign n10028 = P2_P2_ADDRESS_REG_13_ & ~n10026_1;
  assign n10029 = ~n10027 & ~n10028;
  assign n10030 = ~P4_DATAO_REG_13_ & ~P4_DATAO_REG_20_;
  assign n10031_1 = ~P4_DATAO_REG_3_ & n10030;
  assign n10032 = ~P4_DATAO_REG_27_ & n10031_1;
  assign n10033 = ~P4_DATAO_REG_2_ & n10032;
  assign n10034 = ~P4_DATAO_REG_5_ & n10033;
  assign n10035 = ~P4_DATAO_REG_15_ & n10034;
  assign n10036_1 = ~P4_DATAO_REG_21_ & ~P4_DATAO_REG_26_;
  assign n10037 = ~P4_DATAO_REG_28_ & n10036_1;
  assign n10038 = ~P4_DATAO_REG_6_ & n10037;
  assign n10039 = ~P4_DATAO_REG_12_ & n10038;
  assign n10040 = ~P4_DATAO_REG_14_ & n10039;
  assign n10041_1 = ~P4_DATAO_REG_4_ & n10040;
  assign n10042 = ~P4_DATAO_REG_0_ & ~P4_DATAO_REG_16_;
  assign n10043 = ~P4_DATAO_REG_18_ & n10042;
  assign n10044 = ~P4_DATAO_REG_8_ & n10043;
  assign n10045 = ~P4_DATAO_REG_23_ & n10044;
  assign n10046_1 = ~P4_DATAO_REG_1_ & n10045;
  assign n10047 = ~P4_DATAO_REG_11_ & n10046_1;
  assign n10048 = ~P4_DATAO_REG_9_ & ~P4_DATAO_REG_17_;
  assign n10049 = ~P4_DATAO_REG_7_ & n10048;
  assign n10050 = ~P4_DATAO_REG_22_ & n10049;
  assign n10051_1 = ~P4_DATAO_REG_10_ & n10050;
  assign n10052 = ~P4_DATAO_REG_19_ & n10051_1;
  assign n10053 = ~P4_DATAO_REG_25_ & n10052;
  assign n10054 = ~P4_DATAO_REG_24_ & n10053;
  assign n10055 = n10035 & n10041_1;
  assign n10056_1 = n10047 & n10055;
  assign n10057 = n10054 & n10056_1;
  assign n10058 = P4_DATAO_REG_29_ & ~n10057;
  assign n10059 = ~P4_DATAO_REG_30_ & ~n10058;
  assign n10060 = ~P4_DATAO_REG_31_ & ~n10059;
  assign n10061_1 = ~P3_WR_REG & ~n10060;
  assign n10062 = ~n10029 & n10061_1;
  assign n10063 = ~P3_WR_REG & n10060;
  assign n10064 = P2_P1_ADDRESS_REG_13_ & n10063;
  assign n10065 = ~n10021_1 & ~n10062;
  assign n10066_1 = ~n10064 & n10065;
  assign n10067 = P4_ADDR_REG_3_ & P4_WR_REG;
  assign n10068 = P1_P3_DATAO_REG_30_ & ~P1_P3_DATAO_REG_31_;
  assign n10069 = P1_P1_DATAO_REG_30_ & ~P1_P1_DATAO_REG_31_;
  assign n10070 = P1_P2_DATAO_REG_30_ & ~P1_P2_DATAO_REG_31_;
  assign n10071_1 = ~n10068 & ~n10069;
  assign n10072 = ~n10070 & n10071_1;
  assign n10073 = P1_P3_ADDRESS_REG_3_ & n10072;
  assign n10074 = P1_P2_ADDRESS_REG_3_ & ~n10072;
  assign n10075 = ~n10073 & ~n10074;
  assign n10076_1 = ~P3_DATAO_REG_3_ & ~P3_DATAO_REG_20_;
  assign n10077 = ~P3_DATAO_REG_27_ & n10076_1;
  assign n10078 = ~P3_DATAO_REG_12_ & n10077;
  assign n10079 = ~P3_DATAO_REG_2_ & n10078;
  assign n10080 = ~P3_DATAO_REG_5_ & n10079;
  assign n10081_1 = ~P3_DATAO_REG_15_ & n10080;
  assign n10082 = ~P3_DATAO_REG_6_ & ~P3_DATAO_REG_13_;
  assign n10083 = ~P3_DATAO_REG_23_ & n10082;
  assign n10084 = ~P3_DATAO_REG_4_ & n10083;
  assign n10085 = ~P3_DATAO_REG_14_ & n10084;
  assign n10086_1 = ~P3_DATAO_REG_26_ & n10085;
  assign n10087 = ~P3_DATAO_REG_21_ & n10086_1;
  assign n10088 = ~P3_DATAO_REG_8_ & ~P3_DATAO_REG_16_;
  assign n10089 = ~P3_DATAO_REG_24_ & n10088;
  assign n10090 = ~P3_DATAO_REG_18_ & n10089;
  assign n10091_1 = ~P3_DATAO_REG_11_ & n10090;
  assign n10092 = ~P3_DATAO_REG_0_ & n10091_1;
  assign n10093 = ~P3_DATAO_REG_1_ & n10092;
  assign n10094 = ~P3_DATAO_REG_9_ & ~P3_DATAO_REG_17_;
  assign n10095 = ~P3_DATAO_REG_7_ & n10094;
  assign n10096_1 = ~P3_DATAO_REG_22_ & n10095;
  assign n10097 = ~P3_DATAO_REG_25_ & n10096_1;
  assign n10098 = ~P3_DATAO_REG_10_ & n10097;
  assign n10099 = ~P3_DATAO_REG_19_ & n10098;
  assign n10100 = n10081_1 & n10087;
  assign n10101_1 = n10093 & n10100;
  assign n10102 = n10099 & n10101_1;
  assign n10103 = P3_DATAO_REG_28_ & ~n10102;
  assign n10104 = ~P3_DATAO_REG_29_ & ~n10103;
  assign n10105 = ~P3_DATAO_REG_30_ & n10104;
  assign n10106_1 = ~P3_DATAO_REG_31_ & ~n10105;
  assign n10107 = ~P4_WR_REG & ~n10106_1;
  assign n10108 = ~n10075 & n10107;
  assign n10109 = ~P4_WR_REG & n10106_1;
  assign n10110 = P1_P1_ADDRESS_REG_3_ & n10109;
  assign n10111_1 = ~n10067 & ~n10108;
  assign n10112 = ~n10110 & n10111_1;
  assign n10113 = ~n10066_1 & ~n10112;
  assign n10114 = P3_ADDR_REG_12_ & P3_WR_REG;
  assign n10115 = P2_P3_ADDRESS_REG_12_ & n10026_1;
  assign n10116_1 = P2_P2_ADDRESS_REG_12_ & ~n10026_1;
  assign n10117 = ~n10115 & ~n10116_1;
  assign n10118 = n10061_1 & ~n10117;
  assign n10119 = P2_P1_ADDRESS_REG_12_ & n10063;
  assign n10120 = ~n10114 & ~n10118;
  assign n10121_1 = ~n10119 & n10120;
  assign n10122 = ~n10112 & ~n10121_1;
  assign n10123 = P3_ADDR_REG_10_ & P3_WR_REG;
  assign n10124 = P2_P3_ADDRESS_REG_10_ & n10026_1;
  assign n10125 = P2_P2_ADDRESS_REG_10_ & ~n10026_1;
  assign n10126_1 = ~n10124 & ~n10125;
  assign n10127 = n10061_1 & ~n10126_1;
  assign n10128 = P2_P1_ADDRESS_REG_10_ & n10063;
  assign n10129 = ~n10123 & ~n10127;
  assign n10130 = ~n10128 & n10129;
  assign n10131_1 = P4_ADDR_REG_4_ & P4_WR_REG;
  assign n10132 = P1_P3_ADDRESS_REG_4_ & n10072;
  assign n10133 = P1_P2_ADDRESS_REG_4_ & ~n10072;
  assign n10134 = ~n10132 & ~n10133;
  assign n10135 = n10107 & ~n10134;
  assign n10136_1 = P1_P1_ADDRESS_REG_4_ & n10109;
  assign n10137 = ~n10131_1 & ~n10135;
  assign n10138 = ~n10136_1 & n10137;
  assign n10139 = ~n10130 & ~n10138;
  assign n10140 = P3_ADDR_REG_8_ & P3_WR_REG;
  assign n10141_1 = P2_P3_ADDRESS_REG_8_ & n10026_1;
  assign n10142 = P2_P2_ADDRESS_REG_8_ & ~n10026_1;
  assign n10143 = ~n10141_1 & ~n10142;
  assign n10144 = n10061_1 & ~n10143;
  assign n10145 = P2_P1_ADDRESS_REG_8_ & n10063;
  assign n10146_1 = ~n10140 & ~n10144;
  assign n10147 = ~n10145 & n10146_1;
  assign n10148 = P4_ADDR_REG_5_ & P4_WR_REG;
  assign n10149 = P1_P3_ADDRESS_REG_5_ & n10072;
  assign n10150 = P1_P2_ADDRESS_REG_5_ & ~n10072;
  assign n10151_1 = ~n10149 & ~n10150;
  assign n10152 = n10107 & ~n10151_1;
  assign n10153 = P1_P1_ADDRESS_REG_5_ & n10109;
  assign n10154 = ~n10148 & ~n10152;
  assign n10155 = ~n10153 & n10154;
  assign n10156_1 = ~n10147 & ~n10155;
  assign n10157 = P3_ADDR_REG_5_ & P3_WR_REG;
  assign n10158 = P2_P3_ADDRESS_REG_5_ & n10026_1;
  assign n10159 = P2_P2_ADDRESS_REG_5_ & ~n10026_1;
  assign n10160 = ~n10158 & ~n10159;
  assign n10161_1 = n10061_1 & ~n10160;
  assign n10162 = P2_P1_ADDRESS_REG_5_ & n10063;
  assign n10163 = ~n10157 & ~n10161_1;
  assign n10164 = ~n10162 & n10163;
  assign n10165 = P4_ADDR_REG_7_ & P4_WR_REG;
  assign n10166_1 = P1_P3_ADDRESS_REG_7_ & n10072;
  assign n10167 = P1_P2_ADDRESS_REG_7_ & ~n10072;
  assign n10168 = ~n10166_1 & ~n10167;
  assign n10169 = n10107 & ~n10168;
  assign n10170 = P1_P1_ADDRESS_REG_7_ & n10109;
  assign n10171_1 = ~n10165 & ~n10169;
  assign n10172 = ~n10170 & n10171_1;
  assign n10173 = ~n10164 & ~n10172;
  assign n10174 = P3_ADDR_REG_4_ & P3_WR_REG;
  assign n10175 = P2_P3_ADDRESS_REG_4_ & n10026_1;
  assign n10176_1 = P2_P2_ADDRESS_REG_4_ & ~n10026_1;
  assign n10177 = ~n10175 & ~n10176_1;
  assign n10178 = n10061_1 & ~n10177;
  assign n10179 = P2_P1_ADDRESS_REG_4_ & n10063;
  assign n10180 = ~n10174 & ~n10178;
  assign n10181_1 = ~n10179 & n10180;
  assign n10182 = ~n10172 & ~n10181_1;
  assign n10183 = P4_ADDR_REG_8_ & P4_WR_REG;
  assign n10184 = P1_P3_ADDRESS_REG_8_ & n10072;
  assign n10185 = P1_P2_ADDRESS_REG_8_ & ~n10072;
  assign n10186_1 = ~n10184 & ~n10185;
  assign n10187 = n10107 & ~n10186_1;
  assign n10188 = P1_P1_ADDRESS_REG_8_ & n10109;
  assign n10189 = ~n10183 & ~n10187;
  assign n10190 = ~n10188 & n10189;
  assign n10191_1 = P3_ADDR_REG_2_ & P3_WR_REG;
  assign n10192 = P2_P3_ADDRESS_REG_2_ & n10026_1;
  assign n10193 = P2_P2_ADDRESS_REG_2_ & ~n10026_1;
  assign n10194 = ~n10192 & ~n10193;
  assign n10195 = n10061_1 & ~n10194;
  assign n10196_1 = P2_P1_ADDRESS_REG_2_ & n10063;
  assign n10197 = ~n10191_1 & ~n10195;
  assign n10198 = ~n10196_1 & n10197;
  assign n10199 = ~n10190 & ~n10198;
  assign n10200 = P4_ADDR_REG_9_ & P4_WR_REG;
  assign n10201_1 = P1_P3_ADDRESS_REG_9_ & n10072;
  assign n10202 = P1_P2_ADDRESS_REG_9_ & ~n10072;
  assign n10203 = ~n10201_1 & ~n10202;
  assign n10204 = n10107 & ~n10203;
  assign n10205 = P1_P1_ADDRESS_REG_9_ & n10109;
  assign n10206_1 = ~n10200 & ~n10204;
  assign n10207 = ~n10205 & n10206_1;
  assign n10208 = P3_ADDR_REG_1_ & P3_WR_REG;
  assign n10209 = P2_P1_ADDRESS_REG_1_ & n10060;
  assign n10210 = P2_P3_ADDRESS_REG_1_ & n10026_1;
  assign n10211_1 = P2_P2_ADDRESS_REG_1_ & ~n10026_1;
  assign n10212 = ~n10210 & ~n10211_1;
  assign n10213 = ~n10060 & ~n10212;
  assign n10214 = ~n10209 & ~n10213;
  assign n10215 = ~P3_WR_REG & ~n10214;
  assign n10216_1 = ~n10208 & ~n10215;
  assign n10217 = P3_ADDR_REG_0_ & P3_WR_REG;
  assign n10218 = P2_P1_ADDRESS_REG_0_ & n10060;
  assign n10219 = P2_P3_ADDRESS_REG_0_ & n10026_1;
  assign n10220 = P2_P2_ADDRESS_REG_0_ & ~n10026_1;
  assign n10221_1 = ~n10219 & ~n10220;
  assign n10222 = ~n10060 & ~n10221_1;
  assign n10223 = ~n10218 & ~n10222;
  assign n10224 = ~P3_WR_REG & ~n10223;
  assign n10225 = ~n10217 & ~n10224;
  assign n10226_1 = ~n10216_1 & n10225;
  assign n10227 = P4_ADDR_REG_10_ & P4_WR_REG;
  assign n10228 = P1_P3_ADDRESS_REG_10_ & n10072;
  assign n10229 = P1_P2_ADDRESS_REG_10_ & ~n10072;
  assign n10230 = ~n10228 & ~n10229;
  assign n10231_1 = n10107 & ~n10230;
  assign n10232 = P1_P1_ADDRESS_REG_10_ & n10109;
  assign n10233 = ~n10227 & ~n10231_1;
  assign n10234 = ~n10232 & n10233;
  assign n10235 = ~n10216_1 & n10234;
  assign n10236_1 = ~n10226_1 & ~n10235;
  assign n10237 = ~n10207 & ~n10236_1;
  assign n10238 = n10216_1 & ~n10225;
  assign n10239 = n10207 & ~n10225;
  assign n10240 = ~n10238 & ~n10239;
  assign n10241_1 = ~n10234 & ~n10240;
  assign n10242 = ~n10237 & ~n10241_1;
  assign n10243 = n10199 & ~n10242;
  assign n10244 = ~n10216_1 & ~n10225;
  assign n10245 = ~n10190 & ~n10207;
  assign n10246_1 = n10244 & n10245;
  assign n10247 = ~n10199 & n10242;
  assign n10248 = n10246_1 & ~n10247;
  assign n10249 = ~n10243 & ~n10248;
  assign n10250 = P3_ADDR_REG_3_ & P3_WR_REG;
  assign n10251_1 = P2_P3_ADDRESS_REG_3_ & n10026_1;
  assign n10252 = P2_P2_ADDRESS_REG_3_ & ~n10026_1;
  assign n10253 = ~n10251_1 & ~n10252;
  assign n10254 = n10061_1 & ~n10253;
  assign n10255 = P2_P1_ADDRESS_REG_3_ & n10063;
  assign n10256_1 = ~n10250 & ~n10254;
  assign n10257 = ~n10255 & n10256_1;
  assign n10258 = ~n10190 & ~n10257;
  assign n10259 = ~n10198 & ~n10207;
  assign n10260 = P4_ADDR_REG_11_ & P4_WR_REG;
  assign n10261_1 = P1_P3_ADDRESS_REG_11_ & n10072;
  assign n10262 = P1_P2_ADDRESS_REG_11_ & ~n10072;
  assign n10263 = ~n10261_1 & ~n10262;
  assign n10264 = n10107 & ~n10263;
  assign n10265 = P1_P1_ADDRESS_REG_11_ & n10109;
  assign n10266_1 = ~n10260 & ~n10264;
  assign n10267 = ~n10265 & n10266_1;
  assign n10268 = ~n10216_1 & n10267;
  assign n10269 = ~n10226_1 & ~n10268;
  assign n10270 = ~n10234 & ~n10269;
  assign n10271_1 = ~n10225 & n10234;
  assign n10272 = ~n10238 & ~n10271_1;
  assign n10273 = ~n10267 & ~n10272;
  assign n10274 = ~n10270 & ~n10273;
  assign n10275 = n10259 & ~n10274;
  assign n10276_1 = ~n10259 & n10274;
  assign n10277 = ~n10207 & ~n10234;
  assign n10278 = n10244 & n10277;
  assign n10279 = ~n10275 & ~n10276_1;
  assign n10280 = ~n10278 & n10279;
  assign n10281_1 = n10278 & ~n10279;
  assign n10282 = ~n10280 & ~n10281_1;
  assign n10283 = n10258 & ~n10282;
  assign n10284 = ~n10258 & n10282;
  assign n10285 = ~n10283 & ~n10284;
  assign n10286_1 = n10249 & ~n10285;
  assign n10287 = ~n10258 & ~n10282;
  assign n10288 = ~n10249 & n10287;
  assign n10289 = ~n10249 & n10258;
  assign n10290 = n10282 & n10289;
  assign n10291_1 = ~n10286_1 & ~n10288;
  assign n10292 = ~n10290 & n10291_1;
  assign n10293 = n10182 & n10292;
  assign n10294 = ~n10182 & ~n10292;
  assign n10295 = ~n10172 & ~n10257;
  assign n10296_1 = ~n10172 & ~n10190;
  assign n10297 = n10244 & n10296_1;
  assign n10298 = ~n10172 & ~n10198;
  assign n10299 = n10297 & n10298;
  assign n10300 = ~n10297 & ~n10298;
  assign n10301_1 = n10190 & ~n10225;
  assign n10302 = ~n10238 & ~n10301_1;
  assign n10303 = ~n10207 & ~n10302;
  assign n10304 = n10207 & ~n10216_1;
  assign n10305 = ~n10226_1 & ~n10304;
  assign n10306_1 = ~n10190 & ~n10305;
  assign n10307 = ~n10303 & ~n10306_1;
  assign n10308 = ~n10300 & ~n10307;
  assign n10309 = ~n10299 & ~n10308;
  assign n10310 = n10295 & ~n10309;
  assign n10311_1 = ~n10243 & ~n10247;
  assign n10312 = ~n10246_1 & n10311_1;
  assign n10313 = n10246_1 & ~n10311_1;
  assign n10314 = ~n10312 & ~n10313;
  assign n10315 = n10295 & ~n10314;
  assign n10316_1 = ~n10309 & ~n10314;
  assign n10317 = ~n10310 & ~n10315;
  assign n10318 = ~n10316_1 & n10317;
  assign n10319 = ~n10294 & ~n10318;
  assign n10320 = ~n10293 & ~n10319;
  assign n10321_1 = n10173 & ~n10320;
  assign n10322 = ~n10249 & ~n10282;
  assign n10323 = ~n10283 & ~n10289;
  assign n10324 = ~n10322 & n10323;
  assign n10325 = ~n10181_1 & ~n10190;
  assign n10326_1 = ~n10276_1 & n10278;
  assign n10327 = ~n10275 & ~n10326_1;
  assign n10328 = ~n10207 & ~n10257;
  assign n10329 = ~n10198 & ~n10234;
  assign n10330 = P4_ADDR_REG_12_ & P4_WR_REG;
  assign n10331_1 = P1_P3_ADDRESS_REG_12_ & n10072;
  assign n10332 = P1_P2_ADDRESS_REG_12_ & ~n10072;
  assign n10333 = ~n10331_1 & ~n10332;
  assign n10334 = n10107 & ~n10333;
  assign n10335 = P1_P1_ADDRESS_REG_12_ & n10109;
  assign n10336_1 = ~n10330 & ~n10334;
  assign n10337 = ~n10335 & n10336_1;
  assign n10338 = ~n10216_1 & n10337;
  assign n10339 = ~n10226_1 & ~n10338;
  assign n10340 = ~n10267 & ~n10339;
  assign n10341_1 = ~n10225 & n10267;
  assign n10342 = ~n10238 & ~n10341_1;
  assign n10343 = ~n10337 & ~n10342;
  assign n10344 = ~n10340 & ~n10343;
  assign n10345 = n10329 & ~n10344;
  assign n10346_1 = ~n10329 & n10344;
  assign n10347 = ~n10234 & ~n10267;
  assign n10348 = n10244 & n10347;
  assign n10349 = ~n10345 & ~n10346_1;
  assign n10350 = ~n10348 & n10349;
  assign n10351_1 = n10348 & ~n10349;
  assign n10352 = ~n10350 & ~n10351_1;
  assign n10353 = n10328 & ~n10352;
  assign n10354 = ~n10328 & n10352;
  assign n10355 = ~n10353 & ~n10354;
  assign n10356_1 = n10327 & ~n10355;
  assign n10357 = ~n10328 & ~n10352;
  assign n10358 = ~n10327 & n10357;
  assign n10359 = ~n10327 & n10328;
  assign n10360 = n10352 & n10359;
  assign n10361_1 = ~n10356_1 & ~n10358;
  assign n10362 = ~n10360 & n10361_1;
  assign n10363 = n10325 & ~n10362;
  assign n10364 = ~n10325 & n10362;
  assign n10365 = ~n10363 & ~n10364;
  assign n10366_1 = n10324 & ~n10365;
  assign n10367 = n10325 & n10362;
  assign n10368 = ~n10325 & ~n10362;
  assign n10369 = ~n10367 & ~n10368;
  assign n10370 = ~n10324 & ~n10369;
  assign n10371_1 = ~n10366_1 & ~n10370;
  assign n10372 = n10173 & ~n10371_1;
  assign n10373 = ~n10320 & ~n10371_1;
  assign n10374 = ~n10321_1 & ~n10372;
  assign n10375 = ~n10373 & n10374;
  assign n10376_1 = P3_ADDR_REG_6_ & P3_WR_REG;
  assign n10377 = P2_P3_ADDRESS_REG_6_ & n10026_1;
  assign n10378 = P2_P2_ADDRESS_REG_6_ & ~n10026_1;
  assign n10379 = ~n10377 & ~n10378;
  assign n10380 = n10061_1 & ~n10379;
  assign n10381_1 = P2_P1_ADDRESS_REG_6_ & n10063;
  assign n10382 = ~n10376_1 & ~n10380;
  assign n10383 = ~n10381_1 & n10382;
  assign n10384 = ~n10172 & ~n10383;
  assign n10385 = ~n10327 & ~n10352;
  assign n10386_1 = ~n10353 & ~n10359;
  assign n10387 = ~n10385 & n10386_1;
  assign n10388 = ~n10181_1 & ~n10207;
  assign n10389 = ~n10346_1 & n10348;
  assign n10390 = ~n10345 & ~n10389;
  assign n10391_1 = ~n10234 & ~n10257;
  assign n10392 = ~n10198 & ~n10267;
  assign n10393 = P4_ADDR_REG_13_ & P4_WR_REG;
  assign n10394 = P1_P3_ADDRESS_REG_13_ & n10072;
  assign n10395 = P1_P2_ADDRESS_REG_13_ & ~n10072;
  assign n10396_1 = ~n10394 & ~n10395;
  assign n10397 = n10107 & ~n10396_1;
  assign n10398 = P1_P1_ADDRESS_REG_13_ & n10109;
  assign n10399 = ~n10393 & ~n10397;
  assign n10400 = ~n10398 & n10399;
  assign n10401_1 = ~n10216_1 & n10400;
  assign n10402 = ~n10226_1 & ~n10401_1;
  assign n10403 = ~n10337 & ~n10402;
  assign n10404 = ~n10225 & n10337;
  assign n10405 = ~n10238 & ~n10404;
  assign n10406_1 = ~n10400 & ~n10405;
  assign n10407 = ~n10403 & ~n10406_1;
  assign n10408 = n10392 & ~n10407;
  assign n10409 = ~n10392 & n10407;
  assign n10410 = ~n10267 & ~n10337;
  assign n10411_1 = n10244 & n10410;
  assign n10412 = ~n10408 & ~n10409;
  assign n10413 = ~n10411_1 & n10412;
  assign n10414 = n10411_1 & ~n10412;
  assign n10415 = ~n10413 & ~n10414;
  assign n10416_1 = n10391_1 & ~n10415;
  assign n10417 = ~n10391_1 & n10415;
  assign n10418 = ~n10416_1 & ~n10417;
  assign n10419 = n10390 & ~n10418;
  assign n10420 = ~n10391_1 & ~n10415;
  assign n10421_1 = ~n10390 & n10420;
  assign n10422 = ~n10390 & n10391_1;
  assign n10423 = n10415 & n10422;
  assign n10424 = ~n10419 & ~n10421_1;
  assign n10425 = ~n10423 & n10424;
  assign n10426_1 = n10388 & ~n10425;
  assign n10427 = ~n10388 & n10425;
  assign n10428 = ~n10426_1 & ~n10427;
  assign n10429 = n10387 & ~n10428;
  assign n10430 = n10388 & n10425;
  assign n10431_1 = ~n10388 & ~n10425;
  assign n10432 = ~n10430 & ~n10431_1;
  assign n10433 = ~n10387 & ~n10432;
  assign n10434 = ~n10429 & ~n10433;
  assign n10435 = ~n10164 & ~n10190;
  assign n10436_1 = ~n10324 & ~n10368;
  assign n10437 = ~n10367 & ~n10436_1;
  assign n10438 = n10435 & ~n10437;
  assign n10439 = ~n10435 & n10437;
  assign n10440 = ~n10438 & ~n10439;
  assign n10441_1 = n10434 & ~n10440;
  assign n10442 = ~n10435 & ~n10437;
  assign n10443 = ~n10434 & n10442;
  assign n10444 = ~n10434 & n10435;
  assign n10445 = n10437 & n10444;
  assign n10446_1 = ~n10441_1 & ~n10443;
  assign n10447 = ~n10445 & n10446_1;
  assign n10448 = n10384 & ~n10447;
  assign n10449 = ~n10384 & n10447;
  assign n10450 = ~n10448 & ~n10449;
  assign n10451_1 = n10375 & ~n10450;
  assign n10452 = n10384 & n10447;
  assign n10453 = ~n10384 & ~n10447;
  assign n10454 = ~n10452 & ~n10453;
  assign n10455 = ~n10375 & ~n10454;
  assign n10456_1 = ~n10451_1 & ~n10455;
  assign n10457 = P4_ADDR_REG_6_ & P4_WR_REG;
  assign n10458 = P1_P3_ADDRESS_REG_6_ & n10072;
  assign n10459 = P1_P2_ADDRESS_REG_6_ & ~n10072;
  assign n10460 = ~n10458 & ~n10459;
  assign n10461_1 = n10107 & ~n10460;
  assign n10462 = P1_P1_ADDRESS_REG_6_ & n10109;
  assign n10463 = ~n10457 & ~n10461_1;
  assign n10464 = ~n10462 & n10463;
  assign n10465 = P3_ADDR_REG_7_ & P3_WR_REG;
  assign n10466_1 = P2_P3_ADDRESS_REG_7_ & n10026_1;
  assign n10467 = P2_P2_ADDRESS_REG_7_ & ~n10026_1;
  assign n10468 = ~n10466_1 & ~n10467;
  assign n10469 = n10061_1 & ~n10468;
  assign n10470 = P2_P1_ADDRESS_REG_7_ & n10063;
  assign n10471_1 = ~n10465 & ~n10469;
  assign n10472 = ~n10470 & n10471_1;
  assign n10473 = ~n10464 & ~n10472;
  assign n10474 = ~n10383 & ~n10464;
  assign n10475 = ~n10173 & n10371_1;
  assign n10476_1 = ~n10372 & ~n10475;
  assign n10477 = n10320 & ~n10476_1;
  assign n10478 = ~n10173 & ~n10371_1;
  assign n10479 = ~n10320 & n10478;
  assign n10480 = n10321_1 & n10371_1;
  assign n10481_1 = ~n10477 & ~n10479;
  assign n10482 = ~n10480 & n10481_1;
  assign n10483 = n10474 & n10482;
  assign n10484 = ~n10474 & ~n10482;
  assign n10485 = ~n10164 & ~n10464;
  assign n10486_1 = n10182 & ~n10292;
  assign n10487 = ~n10182 & n10292;
  assign n10488 = ~n10486_1 & ~n10487;
  assign n10489 = n10318 & ~n10488;
  assign n10490 = ~n10293 & ~n10294;
  assign n10491_1 = ~n10318 & ~n10490;
  assign n10492 = ~n10489 & ~n10491_1;
  assign n10493 = n10485 & ~n10492;
  assign n10494 = ~n10295 & n10314;
  assign n10495 = ~n10315 & ~n10494;
  assign n10496_1 = n10309 & ~n10495;
  assign n10497 = ~n10295 & ~n10314;
  assign n10498 = ~n10309 & n10497;
  assign n10499 = n10310 & n10314;
  assign n10500 = ~n10496_1 & ~n10498;
  assign n10501_1 = ~n10499 & n10500;
  assign n10502 = ~n10181_1 & ~n10464;
  assign n10503 = n10501_1 & n10502;
  assign n10504 = ~n10501_1 & ~n10502;
  assign n10505 = ~n10257 & ~n10464;
  assign n10506_1 = n10298 & ~n10307;
  assign n10507 = ~n10298 & n10307;
  assign n10508 = ~n10506_1 & ~n10507;
  assign n10509 = ~n10297 & n10508;
  assign n10510 = n10297 & n10507;
  assign n10511_1 = n10299 & ~n10307;
  assign n10512 = ~n10509 & ~n10510;
  assign n10513 = ~n10511_1 & n10512;
  assign n10514 = n10505 & ~n10513;
  assign n10515 = ~n10172 & ~n10464;
  assign n10516_1 = n10244 & n10515;
  assign n10517 = ~n10198 & ~n10464;
  assign n10518 = n10516_1 & n10517;
  assign n10519 = ~n10516_1 & ~n10517;
  assign n10520 = n10172 & ~n10225;
  assign n10521_1 = ~n10238 & ~n10520;
  assign n10522 = ~n10190 & ~n10521_1;
  assign n10523 = n10190 & ~n10216_1;
  assign n10524 = ~n10226_1 & ~n10523;
  assign n10525 = ~n10172 & ~n10524;
  assign n10526_1 = ~n10522 & ~n10525;
  assign n10527 = ~n10519 & ~n10526_1;
  assign n10528 = ~n10518 & ~n10527;
  assign n10529 = n10505 & ~n10528;
  assign n10530 = ~n10513 & ~n10528;
  assign n10531_1 = ~n10514 & ~n10529;
  assign n10532 = ~n10530 & n10531_1;
  assign n10533 = ~n10504 & ~n10532;
  assign n10534 = ~n10503 & ~n10533;
  assign n10535 = n10485 & ~n10534;
  assign n10536_1 = ~n10492 & ~n10534;
  assign n10537 = ~n10493 & ~n10535;
  assign n10538 = ~n10536_1 & n10537;
  assign n10539 = ~n10484 & ~n10538;
  assign n10540 = ~n10483 & ~n10539;
  assign n10541_1 = n10473 & ~n10540;
  assign n10542 = ~n10473 & n10540;
  assign n10543 = ~n10541_1 & ~n10542;
  assign n10544 = n10456_1 & ~n10543;
  assign n10545 = ~n10473 & ~n10540;
  assign n10546_1 = ~n10456_1 & n10545;
  assign n10547 = ~n10456_1 & n10473;
  assign n10548 = n10540 & n10547;
  assign n10549 = ~n10544 & ~n10546_1;
  assign n10550 = ~n10548 & n10549;
  assign n10551_1 = n10156_1 & n10550;
  assign n10552 = ~n10156_1 & ~n10550;
  assign n10553 = ~n10155 & ~n10472;
  assign n10554 = ~n10485 & n10534;
  assign n10555 = ~n10535 & ~n10554;
  assign n10556_1 = n10492 & ~n10555;
  assign n10557 = ~n10485 & ~n10534;
  assign n10558 = ~n10492 & n10557;
  assign n10559 = n10493 & n10534;
  assign n10560 = ~n10556_1 & ~n10558;
  assign n10561_1 = ~n10559 & n10560;
  assign n10562 = ~n10155 & ~n10383;
  assign n10563 = n10561_1 & n10562;
  assign n10564 = ~n10561_1 & ~n10562;
  assign n10565 = ~n10155 & ~n10164;
  assign n10566_1 = ~n10155 & ~n10181_1;
  assign n10567 = ~n10155 & ~n10257;
  assign n10568 = n10517 & ~n10526_1;
  assign n10569 = ~n10517 & n10526_1;
  assign n10570 = ~n10568 & ~n10569;
  assign n10571_1 = ~n10516_1 & n10570;
  assign n10572 = n10516_1 & n10569;
  assign n10573 = n10518 & ~n10526_1;
  assign n10574 = ~n10571_1 & ~n10572;
  assign n10575 = ~n10573 & n10574;
  assign n10576_1 = n10567 & ~n10575;
  assign n10577 = ~n10155 & ~n10464;
  assign n10578 = n10244 & n10577;
  assign n10579 = ~n10155 & ~n10198;
  assign n10580 = n10578 & n10579;
  assign n10581_1 = ~n10578 & ~n10579;
  assign n10582 = ~n10225 & n10464;
  assign n10583 = ~n10238 & ~n10582;
  assign n10584 = ~n10172 & ~n10583;
  assign n10585 = n10172 & ~n10216_1;
  assign n10586_1 = ~n10226_1 & ~n10585;
  assign n10587 = ~n10464 & ~n10586_1;
  assign n10588 = ~n10584 & ~n10587;
  assign n10589 = ~n10581_1 & ~n10588;
  assign n10590 = ~n10580 & ~n10589;
  assign n10591_1 = n10567 & ~n10590;
  assign n10592 = ~n10575 & ~n10590;
  assign n10593 = ~n10576_1 & ~n10591_1;
  assign n10594 = ~n10592 & n10593;
  assign n10595 = n10566_1 & ~n10594;
  assign n10596_1 = ~n10505 & n10513;
  assign n10597 = ~n10514 & ~n10596_1;
  assign n10598 = n10528 & ~n10597;
  assign n10599 = ~n10505 & ~n10513;
  assign n10600 = ~n10528 & n10599;
  assign n10601_1 = n10513 & n10529;
  assign n10602 = ~n10598 & ~n10600;
  assign n10603 = ~n10601_1 & n10602;
  assign n10604 = ~n10566_1 & n10594;
  assign n10605 = n10603 & ~n10604;
  assign n10606_1 = ~n10595 & ~n10605;
  assign n10607 = n10565 & ~n10606_1;
  assign n10608 = ~n10501_1 & n10502;
  assign n10609 = n10501_1 & ~n10502;
  assign n10610 = ~n10608 & ~n10609;
  assign n10611_1 = n10532 & ~n10610;
  assign n10612 = ~n10503 & ~n10504;
  assign n10613 = ~n10532 & ~n10612;
  assign n10614 = ~n10611_1 & ~n10613;
  assign n10615 = n10565 & ~n10614;
  assign n10616_1 = ~n10606_1 & ~n10614;
  assign n10617 = ~n10607 & ~n10615;
  assign n10618 = ~n10616_1 & n10617;
  assign n10619 = ~n10564 & ~n10618;
  assign n10620 = ~n10563 & ~n10619;
  assign n10621_1 = n10553 & ~n10620;
  assign n10622 = n10474 & ~n10482;
  assign n10623 = ~n10474 & n10482;
  assign n10624 = ~n10622 & ~n10623;
  assign n10625 = n10538 & ~n10624;
  assign n10626_1 = ~n10483 & ~n10484;
  assign n10627 = ~n10538 & ~n10626_1;
  assign n10628 = ~n10625 & ~n10627;
  assign n10629 = n10553 & ~n10628;
  assign n10630 = ~n10620 & ~n10628;
  assign n10631_1 = ~n10621_1 & ~n10629;
  assign n10632 = ~n10630 & n10631_1;
  assign n10633 = ~n10552 & ~n10632;
  assign n10634 = ~n10551_1 & ~n10633;
  assign n10635 = P3_ADDR_REG_9_ & P3_WR_REG;
  assign n10636_1 = P2_P3_ADDRESS_REG_9_ & n10026_1;
  assign n10637 = P2_P2_ADDRESS_REG_9_ & ~n10026_1;
  assign n10638 = ~n10636_1 & ~n10637;
  assign n10639 = n10061_1 & ~n10638;
  assign n10640 = P2_P1_ADDRESS_REG_9_ & n10063;
  assign n10641_1 = ~n10635 & ~n10639;
  assign n10642 = ~n10640 & n10641_1;
  assign n10643 = ~n10155 & ~n10642;
  assign n10644 = ~n10147 & ~n10464;
  assign n10645 = ~n10456_1 & ~n10540;
  assign n10646_1 = ~n10541_1 & ~n10547;
  assign n10647 = ~n10645 & n10646_1;
  assign n10648 = n10644 & ~n10647;
  assign n10649 = ~n10644 & n10647;
  assign n10650 = ~n10375 & ~n10453;
  assign n10651_1 = ~n10452 & ~n10650;
  assign n10652 = ~n10172 & ~n10472;
  assign n10653 = ~n10190 & ~n10383;
  assign n10654 = ~n10434 & ~n10437;
  assign n10655 = ~n10438 & ~n10444;
  assign n10656_1 = ~n10654 & n10655;
  assign n10657 = n10653 & ~n10656_1;
  assign n10658 = ~n10653 & n10656_1;
  assign n10659 = ~n10387 & ~n10431_1;
  assign n10660 = ~n10430 & ~n10659;
  assign n10661_1 = ~n10164 & ~n10207;
  assign n10662 = ~n10390 & ~n10415;
  assign n10663 = ~n10416_1 & ~n10422;
  assign n10664 = ~n10662 & n10663;
  assign n10665 = ~n10181_1 & ~n10234;
  assign n10666_1 = ~n10409 & n10411_1;
  assign n10667 = ~n10408 & ~n10666_1;
  assign n10668 = ~n10257 & ~n10267;
  assign n10669 = ~n10198 & ~n10337;
  assign n10670 = P4_ADDR_REG_14_ & P4_WR_REG;
  assign n10671_1 = P1_P3_ADDRESS_REG_14_ & n10072;
  assign n10672 = P1_P2_ADDRESS_REG_14_ & ~n10072;
  assign n10673 = ~n10671_1 & ~n10672;
  assign n10674 = n10107 & ~n10673;
  assign n10675 = P1_P1_ADDRESS_REG_14_ & n10109;
  assign n10676_1 = ~n10670 & ~n10674;
  assign n10677 = ~n10675 & n10676_1;
  assign n10678 = ~n10216_1 & n10677;
  assign n10679 = ~n10226_1 & ~n10678;
  assign n10680 = ~n10400 & ~n10679;
  assign n10681_1 = ~n10225 & n10400;
  assign n10682 = ~n10238 & ~n10681_1;
  assign n10683 = ~n10677 & ~n10682;
  assign n10684 = ~n10680 & ~n10683;
  assign n10685 = n10669 & ~n10684;
  assign n10686_1 = ~n10669 & n10684;
  assign n10687 = ~n10337 & ~n10400;
  assign n10688 = n10244 & n10687;
  assign n10689 = ~n10685 & ~n10686_1;
  assign n10690 = ~n10688 & n10689;
  assign n10691_1 = n10688 & ~n10689;
  assign n10692 = ~n10690 & ~n10691_1;
  assign n10693 = n10668 & ~n10692;
  assign n10694 = ~n10668 & n10692;
  assign n10695 = ~n10693 & ~n10694;
  assign n10696_1 = n10667 & ~n10695;
  assign n10697 = ~n10668 & ~n10692;
  assign n10698 = ~n10667 & n10697;
  assign n10699 = ~n10667 & n10668;
  assign n10700 = n10692 & n10699;
  assign n10701_1 = ~n10696_1 & ~n10698;
  assign n10702 = ~n10700 & n10701_1;
  assign n10703 = n10665 & ~n10702;
  assign n10704 = ~n10665 & n10702;
  assign n10705 = ~n10703 & ~n10704;
  assign n10706_1 = n10664 & ~n10705;
  assign n10707 = n10665 & n10702;
  assign n10708 = ~n10665 & ~n10702;
  assign n10709 = ~n10707 & ~n10708;
  assign n10710 = ~n10664 & ~n10709;
  assign n10711_1 = ~n10706_1 & ~n10710;
  assign n10712 = n10661_1 & ~n10711_1;
  assign n10713 = ~n10661_1 & n10711_1;
  assign n10714 = ~n10712 & ~n10713;
  assign n10715 = n10660 & ~n10714;
  assign n10716_1 = ~n10661_1 & ~n10711_1;
  assign n10717 = ~n10660 & n10716_1;
  assign n10718 = ~n10660 & n10661_1;
  assign n10719 = n10711_1 & n10718;
  assign n10720 = ~n10715 & ~n10717;
  assign n10721_1 = ~n10719 & n10720;
  assign n10722 = ~n10657 & ~n10658;
  assign n10723 = ~n10721_1 & n10722;
  assign n10724 = n10721_1 & ~n10722;
  assign n10725 = ~n10723 & ~n10724;
  assign n10726_1 = n10652 & ~n10725;
  assign n10727 = ~n10652 & n10725;
  assign n10728 = ~n10726_1 & ~n10727;
  assign n10729 = n10651_1 & ~n10728;
  assign n10730 = ~n10652 & ~n10725;
  assign n10731_1 = ~n10651_1 & n10730;
  assign n10732 = ~n10651_1 & n10652;
  assign n10733 = n10725 & n10732;
  assign n10734 = ~n10729 & ~n10731_1;
  assign n10735 = ~n10733 & n10734;
  assign n10736_1 = ~n10648 & ~n10649;
  assign n10737 = ~n10735 & n10736_1;
  assign n10738 = n10735 & ~n10736_1;
  assign n10739 = ~n10737 & ~n10738;
  assign n10740 = n10643 & ~n10739;
  assign n10741_1 = ~n10643 & n10739;
  assign n10742 = ~n10740 & ~n10741_1;
  assign n10743 = n10634 & ~n10742;
  assign n10744 = ~n10643 & ~n10739;
  assign n10745 = ~n10634 & n10744;
  assign n10746_1 = ~n10634 & n10643;
  assign n10747 = n10739 & n10746_1;
  assign n10748 = ~n10743 & ~n10745;
  assign n10749 = ~n10747 & n10748;
  assign n10750 = n10139 & n10749;
  assign n10751_1 = ~n10139 & ~n10749;
  assign n10752 = ~n10138 & ~n10642;
  assign n10753 = ~n10553 & n10628;
  assign n10754 = ~n10629 & ~n10753;
  assign n10755 = n10620 & ~n10754;
  assign n10756_1 = ~n10553 & ~n10628;
  assign n10757 = ~n10620 & n10756_1;
  assign n10758 = n10621_1 & n10628;
  assign n10759 = ~n10755 & ~n10757;
  assign n10760 = ~n10758 & n10759;
  assign n10761_1 = ~n10138 & ~n10147;
  assign n10762 = n10760 & n10761_1;
  assign n10763 = ~n10760 & ~n10761_1;
  assign n10764 = ~n10138 & ~n10472;
  assign n10765 = ~n10565 & n10614;
  assign n10766_1 = ~n10615 & ~n10765;
  assign n10767 = n10606_1 & ~n10766_1;
  assign n10768 = ~n10565 & ~n10614;
  assign n10769 = ~n10606_1 & n10768;
  assign n10770 = n10607 & n10614;
  assign n10771_1 = ~n10767 & ~n10769;
  assign n10772 = ~n10770 & n10771_1;
  assign n10773 = ~n10138 & ~n10383;
  assign n10774 = n10772 & n10773;
  assign n10775 = ~n10772 & ~n10773;
  assign n10776_1 = ~n10138 & ~n10164;
  assign n10777 = n10566_1 & ~n10603;
  assign n10778 = ~n10566_1 & n10603;
  assign n10779 = ~n10777 & ~n10778;
  assign n10780 = n10594 & ~n10779;
  assign n10781_1 = ~n10566_1 & ~n10603;
  assign n10782 = ~n10594 & n10781_1;
  assign n10783 = n10595 & n10603;
  assign n10784 = ~n10780 & ~n10782;
  assign n10785 = ~n10783 & n10784;
  assign n10786_1 = n10776_1 & ~n10785;
  assign n10787 = ~n10138 & ~n10181_1;
  assign n10788 = ~n10138 & ~n10257;
  assign n10789 = n10579 & ~n10588;
  assign n10790 = ~n10579 & n10588;
  assign n10791_1 = ~n10789 & ~n10790;
  assign n10792 = ~n10578 & n10791_1;
  assign n10793 = n10578 & n10790;
  assign n10794 = n10580 & ~n10588;
  assign n10795 = ~n10792 & ~n10793;
  assign n10796_1 = ~n10794 & n10795;
  assign n10797 = n10788 & ~n10796_1;
  assign n10798 = ~n10138 & ~n10155;
  assign n10799 = n10244 & n10798;
  assign n10800 = ~n10138 & ~n10198;
  assign n10801_1 = n10799 & n10800;
  assign n10802 = ~n10799 & ~n10800;
  assign n10803 = n10155 & ~n10225;
  assign n10804 = ~n10238 & ~n10803;
  assign n10805 = ~n10464 & ~n10804;
  assign n10806_1 = ~n10216_1 & n10464;
  assign n10807 = ~n10226_1 & ~n10806_1;
  assign n10808 = ~n10155 & ~n10807;
  assign n10809 = ~n10805 & ~n10808;
  assign n10810 = ~n10802 & ~n10809;
  assign n10811_1 = ~n10801_1 & ~n10810;
  assign n10812 = n10788 & ~n10811_1;
  assign n10813 = ~n10796_1 & ~n10811_1;
  assign n10814 = ~n10797 & ~n10812;
  assign n10815 = ~n10813 & n10814;
  assign n10816_1 = n10787 & ~n10815;
  assign n10817 = ~n10567 & n10575;
  assign n10818 = ~n10576_1 & ~n10817;
  assign n10819 = n10590 & ~n10818;
  assign n10820 = ~n10567 & ~n10575;
  assign n10821_1 = ~n10590 & n10820;
  assign n10822 = n10575 & n10591_1;
  assign n10823 = ~n10819 & ~n10821_1;
  assign n10824 = ~n10822 & n10823;
  assign n10825 = ~n10787 & n10815;
  assign n10826_1 = n10824 & ~n10825;
  assign n10827 = ~n10816_1 & ~n10826_1;
  assign n10828 = n10776_1 & ~n10827;
  assign n10829 = ~n10785 & ~n10827;
  assign n10830 = ~n10786_1 & ~n10828;
  assign n10831_1 = ~n10829 & n10830;
  assign n10832 = ~n10775 & ~n10831_1;
  assign n10833 = ~n10774 & ~n10832;
  assign n10834 = n10764 & ~n10833;
  assign n10835 = ~n10561_1 & n10562;
  assign n10836_1 = n10561_1 & ~n10562;
  assign n10837 = ~n10835 & ~n10836_1;
  assign n10838 = n10618 & ~n10837;
  assign n10839 = ~n10563 & ~n10564;
  assign n10840 = ~n10618 & ~n10839;
  assign n10841_1 = ~n10838 & ~n10840;
  assign n10842 = n10764 & ~n10841_1;
  assign n10843 = ~n10833 & ~n10841_1;
  assign n10844 = ~n10834 & ~n10842;
  assign n10845 = ~n10843 & n10844;
  assign n10846_1 = ~n10763 & ~n10845;
  assign n10847 = ~n10762 & ~n10846_1;
  assign n10848 = n10752 & ~n10847;
  assign n10849 = n10156_1 & ~n10550;
  assign n10850 = ~n10156_1 & n10550;
  assign n10851_1 = ~n10849 & ~n10850;
  assign n10852 = n10632 & ~n10851_1;
  assign n10853 = ~n10551_1 & ~n10552;
  assign n10854 = ~n10632 & ~n10853;
  assign n10855 = ~n10852 & ~n10854;
  assign n10856_1 = n10752 & ~n10855;
  assign n10857 = ~n10847 & ~n10855;
  assign n10858 = ~n10848 & ~n10856_1;
  assign n10859 = ~n10857 & n10858;
  assign n10860 = ~n10751_1 & ~n10859;
  assign n10861_1 = ~n10750 & ~n10860;
  assign n10862 = P3_ADDR_REG_11_ & P3_WR_REG;
  assign n10863 = P2_P3_ADDRESS_REG_11_ & n10026_1;
  assign n10864 = P2_P2_ADDRESS_REG_11_ & ~n10026_1;
  assign n10865 = ~n10863 & ~n10864;
  assign n10866_1 = n10061_1 & ~n10865;
  assign n10867 = P2_P1_ADDRESS_REG_11_ & n10063;
  assign n10868 = ~n10862 & ~n10866_1;
  assign n10869 = ~n10867 & n10868;
  assign n10870 = ~n10138 & ~n10869;
  assign n10871_1 = ~n10634 & ~n10739;
  assign n10872 = ~n10740 & ~n10746_1;
  assign n10873 = ~n10871_1 & n10872;
  assign n10874 = ~n10130 & ~n10155;
  assign n10875 = ~n10649 & n10735;
  assign n10876_1 = ~n10648 & ~n10875;
  assign n10877 = ~n10464 & ~n10642;
  assign n10878 = ~n10651_1 & ~n10725;
  assign n10879 = ~n10726_1 & ~n10732;
  assign n10880 = ~n10878 & n10879;
  assign n10881_1 = ~n10147 & ~n10172;
  assign n10882 = ~n10658 & n10721_1;
  assign n10883 = ~n10657 & ~n10882;
  assign n10884 = ~n10190 & ~n10472;
  assign n10885 = ~n10660 & ~n10711_1;
  assign n10886_1 = ~n10712 & ~n10718;
  assign n10887 = ~n10885 & n10886_1;
  assign n10888 = ~n10207 & ~n10383;
  assign n10889 = ~n10664 & ~n10708;
  assign n10890 = ~n10707 & ~n10889;
  assign n10891_1 = ~n10164 & ~n10234;
  assign n10892 = ~n10667 & ~n10692;
  assign n10893 = ~n10693 & ~n10699;
  assign n10894 = ~n10892 & n10893;
  assign n10895 = ~n10181_1 & ~n10267;
  assign n10896_1 = ~n10686_1 & n10688;
  assign n10897 = ~n10685 & ~n10896_1;
  assign n10898 = ~n10257 & ~n10337;
  assign n10899 = ~n10198 & ~n10400;
  assign n10900 = P4_ADDR_REG_15_ & P4_WR_REG;
  assign n10901_1 = P1_P3_ADDRESS_REG_15_ & n10072;
  assign n10902 = P1_P2_ADDRESS_REG_15_ & ~n10072;
  assign n10903 = ~n10901_1 & ~n10902;
  assign n10904 = n10107 & ~n10903;
  assign n10905 = P1_P1_ADDRESS_REG_15_ & n10109;
  assign n10906_1 = ~n10900 & ~n10904;
  assign n10907 = ~n10905 & n10906_1;
  assign n10908 = ~n10216_1 & n10907;
  assign n10909 = ~n10226_1 & ~n10908;
  assign n10910 = ~n10677 & ~n10909;
  assign n10911_1 = ~n10225 & n10677;
  assign n10912 = ~n10238 & ~n10911_1;
  assign n10913 = ~n10907 & ~n10912;
  assign n10914 = ~n10910 & ~n10913;
  assign n10915 = n10899 & ~n10914;
  assign n10916_1 = ~n10899 & n10914;
  assign n10917 = ~n10400 & ~n10677;
  assign n10918 = n10244 & n10917;
  assign n10919 = ~n10915 & ~n10916_1;
  assign n10920 = ~n10918 & n10919;
  assign n10921_1 = n10918 & ~n10919;
  assign n10922 = ~n10920 & ~n10921_1;
  assign n10923 = n10898 & ~n10922;
  assign n10924 = ~n10898 & n10922;
  assign n10925 = ~n10923 & ~n10924;
  assign n10926_1 = n10897 & ~n10925;
  assign n10927 = ~n10898 & ~n10922;
  assign n10928 = ~n10897 & n10927;
  assign n10929 = ~n10897 & n10898;
  assign n10930 = n10922 & n10929;
  assign n10931_1 = ~n10926_1 & ~n10928;
  assign n10932 = ~n10930 & n10931_1;
  assign n10933 = n10895 & ~n10932;
  assign n10934 = ~n10895 & n10932;
  assign n10935 = ~n10933 & ~n10934;
  assign n10936_1 = n10894 & ~n10935;
  assign n10937 = n10895 & n10932;
  assign n10938 = ~n10895 & ~n10932;
  assign n10939 = ~n10937 & ~n10938;
  assign n10940 = ~n10894 & ~n10939;
  assign n10941_1 = ~n10936_1 & ~n10940;
  assign n10942 = n10891_1 & ~n10941_1;
  assign n10943 = ~n10891_1 & n10941_1;
  assign n10944 = ~n10942 & ~n10943;
  assign n10945 = n10890 & ~n10944;
  assign n10946_1 = ~n10891_1 & ~n10941_1;
  assign n10947 = ~n10890 & n10946_1;
  assign n10948 = ~n10890 & n10891_1;
  assign n10949 = n10941_1 & n10948;
  assign n10950 = ~n10945 & ~n10947;
  assign n10951_1 = ~n10949 & n10950;
  assign n10952 = n10888 & ~n10951_1;
  assign n10953 = ~n10888 & n10951_1;
  assign n10954 = ~n10952 & ~n10953;
  assign n10955 = n10887 & ~n10954;
  assign n10956_1 = n10888 & n10951_1;
  assign n10957 = ~n10888 & ~n10951_1;
  assign n10958 = ~n10956_1 & ~n10957;
  assign n10959 = ~n10887 & ~n10958;
  assign n10960 = ~n10955 & ~n10959;
  assign n10961_1 = n10884 & ~n10960;
  assign n10962 = ~n10884 & n10960;
  assign n10963 = ~n10961_1 & ~n10962;
  assign n10964 = n10883 & ~n10963;
  assign n10965 = ~n10884 & ~n10960;
  assign n10966_1 = ~n10883 & n10965;
  assign n10967 = ~n10883 & n10884;
  assign n10968 = n10960 & n10967;
  assign n10969 = ~n10964 & ~n10966_1;
  assign n10970 = ~n10968 & n10969;
  assign n10971_1 = n10881_1 & ~n10970;
  assign n10972 = ~n10881_1 & n10970;
  assign n10973 = ~n10971_1 & ~n10972;
  assign n10974 = n10880 & ~n10973;
  assign n10975 = n10881_1 & n10970;
  assign n10976_1 = ~n10881_1 & ~n10970;
  assign n10977 = ~n10975 & ~n10976_1;
  assign n10978 = ~n10880 & ~n10977;
  assign n10979 = ~n10974 & ~n10978;
  assign n10980 = n10877 & ~n10979;
  assign n10981_1 = ~n10877 & n10979;
  assign n10982 = ~n10980 & ~n10981_1;
  assign n10983 = n10876_1 & ~n10982;
  assign n10984 = ~n10877 & ~n10979;
  assign n10985 = ~n10876_1 & n10984;
  assign n10986_1 = ~n10876_1 & n10877;
  assign n10987 = n10979 & n10986_1;
  assign n10988 = ~n10983 & ~n10985;
  assign n10989 = ~n10987 & n10988;
  assign n10990 = n10874 & ~n10989;
  assign n10991_1 = ~n10874 & n10989;
  assign n10992 = ~n10990 & ~n10991_1;
  assign n10993 = n10873 & ~n10992;
  assign n10994 = n10874 & n10989;
  assign n10995 = ~n10874 & ~n10989;
  assign n10996_1 = ~n10994 & ~n10995;
  assign n10997 = ~n10873 & ~n10996_1;
  assign n10998 = ~n10993 & ~n10997;
  assign n10999 = n10870 & ~n10998;
  assign n11000 = ~n10870 & n10998;
  assign n11001_1 = ~n10999 & ~n11000;
  assign n11002 = n10861_1 & ~n11001_1;
  assign n11003 = ~n10870 & ~n10998;
  assign n11004 = ~n10861_1 & n11003;
  assign n11005 = ~n10861_1 & n10870;
  assign n11006_1 = n10998 & n11005;
  assign n11007 = ~n11002 & ~n11004;
  assign n11008 = ~n11006_1 & n11007;
  assign n11009 = n10122 & n11008;
  assign n11010 = ~n10122 & ~n11008;
  assign n11011_1 = ~n10112 & ~n10869;
  assign n11012 = ~n10752 & n10855;
  assign n11013 = ~n10856_1 & ~n11012;
  assign n11014 = n10847 & ~n11013;
  assign n11015 = ~n10752 & ~n10855;
  assign n11016_1 = ~n10847 & n11015;
  assign n11017 = n10848 & n10855;
  assign n11018 = ~n11014 & ~n11016_1;
  assign n11019 = ~n11017 & n11018;
  assign n11020 = ~n10112 & ~n10130;
  assign n11021_1 = n11019 & n11020;
  assign n11022 = ~n11019 & ~n11020;
  assign n11023 = ~n10112 & ~n10642;
  assign n11024 = ~n10764 & n10841_1;
  assign n11025 = ~n10842 & ~n11024;
  assign n11026_1 = n10833 & ~n11025;
  assign n11027 = ~n10764 & ~n10841_1;
  assign n11028 = ~n10833 & n11027;
  assign n11029 = n10834 & n10841_1;
  assign n11030 = ~n11026_1 & ~n11028;
  assign n11031_1 = ~n11029 & n11030;
  assign n11032 = ~n10112 & ~n10147;
  assign n11033 = n11031_1 & n11032;
  assign n11034 = ~n11031_1 & ~n11032;
  assign n11035 = ~n10112 & ~n10472;
  assign n11036_1 = ~n10112 & ~n10383;
  assign n11037 = ~n10112 & ~n10164;
  assign n11038 = n10787 & ~n10824;
  assign n11039 = ~n10787 & n10824;
  assign n11040 = ~n11038 & ~n11039;
  assign n11041_1 = n10815 & ~n11040;
  assign n11042 = ~n10787 & ~n10824;
  assign n11043 = ~n10815 & n11042;
  assign n11044 = n10816_1 & n10824;
  assign n11045 = ~n11041_1 & ~n11043;
  assign n11046_1 = ~n11044 & n11045;
  assign n11047 = n11037 & ~n11046_1;
  assign n11048 = ~n10112 & ~n10181_1;
  assign n11049 = ~n10112 & ~n10257;
  assign n11050 = n10800 & ~n10809;
  assign n11051_1 = ~n10800 & n10809;
  assign n11052 = ~n11050 & ~n11051_1;
  assign n11053 = ~n10799 & n11052;
  assign n11054 = n10799 & n11051_1;
  assign n11055 = n10801_1 & ~n10809;
  assign n11056_1 = ~n11053 & ~n11054;
  assign n11057 = ~n11055 & n11056_1;
  assign n11058 = n11049 & ~n11057;
  assign n11059 = ~n10112 & ~n10138;
  assign n11060 = n10244 & n11059;
  assign n11061_1 = ~n10112 & ~n10198;
  assign n11062 = n11060 & n11061_1;
  assign n11063 = ~n11060 & ~n11061_1;
  assign n11064 = n10138 & ~n10225;
  assign n11065 = ~n10238 & ~n11064;
  assign n11066_1 = ~n10155 & ~n11065;
  assign n11067 = n10155 & ~n10216_1;
  assign n11068 = ~n10226_1 & ~n11067;
  assign n11069 = ~n10138 & ~n11068;
  assign n11070 = ~n11066_1 & ~n11069;
  assign n11071_1 = ~n11063 & ~n11070;
  assign n11072 = ~n11062 & ~n11071_1;
  assign n11073 = n11049 & ~n11072;
  assign n11074 = ~n11057 & ~n11072;
  assign n11075 = ~n11058 & ~n11073;
  assign n11076_1 = ~n11074 & n11075;
  assign n11077 = n11048 & ~n11076_1;
  assign n11078 = ~n10788 & n10796_1;
  assign n11079 = ~n10797 & ~n11078;
  assign n11080 = n10811_1 & ~n11079;
  assign n11081_1 = ~n10788 & ~n10796_1;
  assign n11082 = ~n10811_1 & n11081_1;
  assign n11083 = n10796_1 & n10812;
  assign n11084 = ~n11080 & ~n11082;
  assign n11085 = ~n11083 & n11084;
  assign n11086_1 = ~n11048 & n11076_1;
  assign n11087 = n11085 & ~n11086_1;
  assign n11088 = ~n11077 & ~n11087;
  assign n11089 = n11037 & ~n11088;
  assign n11090 = ~n11046_1 & ~n11088;
  assign n11091_1 = ~n11047 & ~n11089;
  assign n11092 = ~n11090 & n11091_1;
  assign n11093 = n11036_1 & ~n11092;
  assign n11094 = ~n10776_1 & n10785;
  assign n11095 = ~n10786_1 & ~n11094;
  assign n11096_1 = n10827 & ~n11095;
  assign n11097 = ~n10776_1 & ~n10785;
  assign n11098 = ~n10827 & n11097;
  assign n11099 = n10785 & n10828;
  assign n11100 = ~n11096_1 & ~n11098;
  assign n11101_1 = ~n11099 & n11100;
  assign n11102 = ~n11036_1 & n11092;
  assign n11103 = n11101_1 & ~n11102;
  assign n11104 = ~n11093 & ~n11103;
  assign n11105 = n11035 & ~n11104;
  assign n11106_1 = ~n10772 & n10773;
  assign n11107 = n10772 & ~n10773;
  assign n11108 = ~n11106_1 & ~n11107;
  assign n11109 = n10831_1 & ~n11108;
  assign n11110 = ~n10774 & ~n10775;
  assign n11111_1 = ~n10831_1 & ~n11110;
  assign n11112 = ~n11109 & ~n11111_1;
  assign n11113 = n11035 & ~n11112;
  assign n11114 = ~n11104 & ~n11112;
  assign n11115 = ~n11105 & ~n11113;
  assign n11116_1 = ~n11114 & n11115;
  assign n11117 = ~n11034 & ~n11116_1;
  assign n11118 = ~n11033 & ~n11117;
  assign n11119 = n11023 & ~n11118;
  assign n11120 = ~n10760 & n10761_1;
  assign n11121_1 = n10760 & ~n10761_1;
  assign n11122 = ~n11120 & ~n11121_1;
  assign n11123 = n10845 & ~n11122;
  assign n11124 = ~n10762 & ~n10763;
  assign n11125 = ~n10845 & ~n11124;
  assign n11126_1 = ~n11123 & ~n11125;
  assign n11127 = n11023 & ~n11126_1;
  assign n11128 = ~n11118 & ~n11126_1;
  assign n11129 = ~n11119 & ~n11127;
  assign n11130 = ~n11128 & n11129;
  assign n11131_1 = ~n11022 & ~n11130;
  assign n11132 = ~n11021_1 & ~n11131_1;
  assign n11133 = n11011_1 & ~n11132;
  assign n11134 = n10139 & ~n10749;
  assign n11135 = ~n10139 & n10749;
  assign n11136_1 = ~n11134 & ~n11135;
  assign n11137 = n10859 & ~n11136_1;
  assign n11138 = ~n10750 & ~n10751_1;
  assign n11139 = ~n10859 & ~n11138;
  assign n11140 = ~n11137 & ~n11139;
  assign n11141_1 = n11011_1 & ~n11140;
  assign n11142 = ~n11132 & ~n11140;
  assign n11143 = ~n11133 & ~n11141_1;
  assign n11144 = ~n11142 & n11143;
  assign n11145 = ~n11010 & ~n11144;
  assign n11146_1 = ~n11009 & ~n11145;
  assign n11147 = n10113 & ~n11146_1;
  assign n11148 = ~n10121_1 & ~n10138;
  assign n11149 = ~n10861_1 & ~n10998;
  assign n11150 = ~n10999 & ~n11005;
  assign n11151_1 = ~n11149 & n11150;
  assign n11152 = n11148 & ~n11151_1;
  assign n11153 = ~n11148 & n11151_1;
  assign n11154 = ~n10873 & ~n10995;
  assign n11155 = ~n10994 & ~n11154;
  assign n11156_1 = ~n10155 & ~n10869;
  assign n11157 = ~n10876_1 & ~n10979;
  assign n11158 = ~n10980 & ~n10986_1;
  assign n11159 = ~n11157 & n11158;
  assign n11160 = ~n10130 & ~n10464;
  assign n11161_1 = ~n10883 & ~n10960;
  assign n11162 = ~n10961_1 & ~n10967;
  assign n11163 = ~n11161_1 & n11162;
  assign n11164 = ~n10147 & ~n10190;
  assign n11165 = ~n10887 & ~n10957;
  assign n11166_1 = ~n10956_1 & ~n11165;
  assign n11167 = ~n10207 & ~n10472;
  assign n11168 = ~n10890 & ~n10941_1;
  assign n11169 = ~n10942 & ~n10948;
  assign n11170 = ~n11168 & n11169;
  assign n11171_1 = ~n10234 & ~n10383;
  assign n11172 = ~n10894 & ~n10938;
  assign n11173 = ~n10937 & ~n11172;
  assign n11174 = ~n10164 & ~n10267;
  assign n11175 = ~n10897 & ~n10922;
  assign n11176_1 = ~n10923 & ~n10929;
  assign n11177 = ~n11175 & n11176_1;
  assign n11178 = ~n10181_1 & ~n10337;
  assign n11179 = ~n10916_1 & n10918;
  assign n11180 = ~n10915 & ~n11179;
  assign n11181_1 = ~n10257 & ~n10400;
  assign n11182 = ~n10198 & ~n10677;
  assign n11183 = P4_ADDR_REG_16_ & P4_WR_REG;
  assign n11184 = P1_P3_ADDRESS_REG_16_ & n10072;
  assign n11185 = P1_P2_ADDRESS_REG_16_ & ~n10072;
  assign n11186_1 = ~n11184 & ~n11185;
  assign n11187 = n10107 & ~n11186_1;
  assign n11188 = P1_P1_ADDRESS_REG_16_ & n10109;
  assign n11189 = ~n11183 & ~n11187;
  assign n11190 = ~n11188 & n11189;
  assign n11191_1 = ~n10216_1 & n11190;
  assign n11192 = ~n10226_1 & ~n11191_1;
  assign n11193 = ~n10907 & ~n11192;
  assign n11194 = ~n10225 & n10907;
  assign n11195 = ~n10238 & ~n11194;
  assign n11196_1 = ~n11190 & ~n11195;
  assign n11197 = ~n11193 & ~n11196_1;
  assign n11198 = n11182 & ~n11197;
  assign n11199 = ~n11182 & n11197;
  assign n11200 = ~n10677 & ~n10907;
  assign n11201_1 = n10244 & n11200;
  assign n11202 = ~n11198 & ~n11199;
  assign n11203 = ~n11201_1 & n11202;
  assign n11204 = n11201_1 & ~n11202;
  assign n11205 = ~n11203 & ~n11204;
  assign n11206_1 = n11181_1 & ~n11205;
  assign n11207 = ~n11181_1 & n11205;
  assign n11208 = ~n11206_1 & ~n11207;
  assign n11209 = n11180 & ~n11208;
  assign n11210 = ~n11181_1 & ~n11205;
  assign n11211_1 = ~n11180 & n11210;
  assign n11212 = ~n11180 & n11181_1;
  assign n11213 = n11205 & n11212;
  assign n11214 = ~n11209 & ~n11211_1;
  assign n11215 = ~n11213 & n11214;
  assign n11216_1 = n11178 & ~n11215;
  assign n11217 = ~n11178 & n11215;
  assign n11218 = ~n11216_1 & ~n11217;
  assign n11219 = n11177 & ~n11218;
  assign n11220 = n11178 & n11215;
  assign n11221_1 = ~n11178 & ~n11215;
  assign n11222 = ~n11220 & ~n11221_1;
  assign n11223 = ~n11177 & ~n11222;
  assign n11224 = ~n11219 & ~n11223;
  assign n11225 = n11174 & ~n11224;
  assign n11226_1 = ~n11174 & n11224;
  assign n11227 = ~n11225 & ~n11226_1;
  assign n11228 = n11173 & ~n11227;
  assign n11229 = ~n11174 & ~n11224;
  assign n11230 = ~n11173 & n11229;
  assign n11231_1 = ~n11173 & n11174;
  assign n11232 = n11224 & n11231_1;
  assign n11233 = ~n11228 & ~n11230;
  assign n11234 = ~n11232 & n11233;
  assign n11235 = n11171_1 & ~n11234;
  assign n11236_1 = ~n11171_1 & n11234;
  assign n11237 = ~n11235 & ~n11236_1;
  assign n11238 = n11170 & ~n11237;
  assign n11239 = n11171_1 & n11234;
  assign n11240 = ~n11171_1 & ~n11234;
  assign n11241_1 = ~n11239 & ~n11240;
  assign n11242 = ~n11170 & ~n11241_1;
  assign n11243 = ~n11238 & ~n11242;
  assign n11244 = n11167 & ~n11243;
  assign n11245 = ~n11167 & n11243;
  assign n11246_1 = ~n11244 & ~n11245;
  assign n11247 = n11166_1 & ~n11246_1;
  assign n11248 = ~n11167 & ~n11243;
  assign n11249 = ~n11166_1 & n11248;
  assign n11250 = ~n11166_1 & n11167;
  assign n11251_1 = n11243 & n11250;
  assign n11252 = ~n11247 & ~n11249;
  assign n11253 = ~n11251_1 & n11252;
  assign n11254 = n11164 & ~n11253;
  assign n11255 = ~n11164 & n11253;
  assign n11256_1 = ~n11254 & ~n11255;
  assign n11257 = n11163 & ~n11256_1;
  assign n11258 = n11164 & n11253;
  assign n11259 = ~n11164 & ~n11253;
  assign n11260 = ~n11258 & ~n11259;
  assign n11261_1 = ~n11163 & ~n11260;
  assign n11262 = ~n11257 & ~n11261_1;
  assign n11263 = ~n10172 & ~n10642;
  assign n11264 = ~n10880 & ~n10976_1;
  assign n11265 = ~n10975 & ~n11264;
  assign n11266_1 = n11263 & ~n11265;
  assign n11267 = ~n11263 & n11265;
  assign n11268 = ~n11266_1 & ~n11267;
  assign n11269 = n11262 & ~n11268;
  assign n11270 = ~n11263 & ~n11265;
  assign n11271_1 = ~n11262 & n11270;
  assign n11272 = ~n11262 & n11263;
  assign n11273 = n11265 & n11272;
  assign n11274 = ~n11269 & ~n11271_1;
  assign n11275 = ~n11273 & n11274;
  assign n11276_1 = n11160 & ~n11275;
  assign n11277 = ~n11160 & n11275;
  assign n11278 = ~n11276_1 & ~n11277;
  assign n11279 = n11159 & ~n11278;
  assign n11280 = n11160 & n11275;
  assign n11281_1 = ~n11160 & ~n11275;
  assign n11282 = ~n11280 & ~n11281_1;
  assign n11283 = ~n11159 & ~n11282;
  assign n11284 = ~n11279 & ~n11283;
  assign n11285 = n11156_1 & ~n11284;
  assign n11286_1 = ~n11156_1 & n11284;
  assign n11287 = ~n11285 & ~n11286_1;
  assign n11288 = n11155 & ~n11287;
  assign n11289 = ~n11156_1 & ~n11284;
  assign n11290 = ~n11155 & n11289;
  assign n11291_1 = ~n11155 & n11156_1;
  assign n11292 = n11284 & n11291_1;
  assign n11293 = ~n11288 & ~n11290;
  assign n11294 = ~n11292 & n11293;
  assign n11295 = ~n11152 & ~n11153;
  assign n11296_1 = ~n11294 & n11295;
  assign n11297 = n11294 & ~n11295;
  assign n11298 = ~n11296_1 & ~n11297;
  assign n11299 = n10113 & ~n11298;
  assign n11300 = ~n11146_1 & ~n11298;
  assign n11301_1 = ~n11147 & ~n11299;
  assign n11302 = ~n11300 & n11301_1;
  assign n11303 = P3_ADDR_REG_14_ & P3_WR_REG;
  assign n11304 = P2_P3_ADDRESS_REG_14_ & n10026_1;
  assign n11305 = P2_P2_ADDRESS_REG_14_ & ~n10026_1;
  assign n11306_1 = ~n11304 & ~n11305;
  assign n11307 = n10061_1 & ~n11306_1;
  assign n11308 = P2_P1_ADDRESS_REG_14_ & n10063;
  assign n11309 = ~n11303 & ~n11307;
  assign n11310 = ~n11308 & n11309;
  assign n11311_1 = ~n10112 & ~n11310;
  assign n11312 = ~n11153 & n11294;
  assign n11313 = ~n11152 & ~n11312;
  assign n11314 = ~n10066_1 & ~n10138;
  assign n11315 = ~n11155 & ~n11284;
  assign n11316_1 = ~n11285 & ~n11291_1;
  assign n11317 = ~n11315 & n11316_1;
  assign n11318 = ~n10121_1 & ~n10155;
  assign n11319 = ~n11159 & ~n11281_1;
  assign n11320 = ~n11280 & ~n11319;
  assign n11321_1 = ~n10464 & ~n10869;
  assign n11322 = ~n11262 & ~n11265;
  assign n11323 = ~n11266_1 & ~n11272;
  assign n11324 = ~n11322 & n11323;
  assign n11325 = ~n10130 & ~n10172;
  assign n11326_1 = ~n11163 & ~n11259;
  assign n11327 = ~n11258 & ~n11326_1;
  assign n11328 = ~n10190 & ~n10642;
  assign n11329 = ~n11166_1 & ~n11243;
  assign n11330 = ~n11244 & ~n11250;
  assign n11331_1 = ~n11329 & n11330;
  assign n11332 = ~n10147 & ~n10207;
  assign n11333 = ~n11170 & ~n11240;
  assign n11334 = ~n11239 & ~n11333;
  assign n11335 = ~n10234 & ~n10472;
  assign n11336_1 = ~n11173 & ~n11224;
  assign n11337 = ~n11225 & ~n11231_1;
  assign n11338 = ~n11336_1 & n11337;
  assign n11339 = ~n10267 & ~n10383;
  assign n11340 = ~n11180 & ~n11205;
  assign n11341_1 = ~n11206_1 & ~n11212;
  assign n11342 = ~n11340 & n11341_1;
  assign n11343 = ~n10181_1 & ~n10400;
  assign n11344 = ~n11199 & n11201_1;
  assign n11345 = ~n11198 & ~n11344;
  assign n11346_1 = ~n10257 & ~n10677;
  assign n11347 = ~n10198 & ~n10907;
  assign n11348 = P4_ADDR_REG_17_ & P4_WR_REG;
  assign n11349 = P1_P3_ADDRESS_REG_17_ & n10072;
  assign n11350 = P1_P2_ADDRESS_REG_17_ & ~n10072;
  assign n11351_1 = ~n11349 & ~n11350;
  assign n11352 = n10107 & ~n11351_1;
  assign n11353 = P1_P1_ADDRESS_REG_17_ & n10109;
  assign n11354 = ~n11348 & ~n11352;
  assign n11355 = ~n11353 & n11354;
  assign n11356_1 = ~n10216_1 & n11355;
  assign n11357 = ~n10226_1 & ~n11356_1;
  assign n11358 = ~n11190 & ~n11357;
  assign n11359 = ~n10225 & n11190;
  assign n11360 = ~n10238 & ~n11359;
  assign n11361_1 = ~n11355 & ~n11360;
  assign n11362 = ~n11358 & ~n11361_1;
  assign n11363 = n11347 & ~n11362;
  assign n11364 = ~n11347 & n11362;
  assign n11365 = ~n10907 & ~n11190;
  assign n11366_1 = n10244 & n11365;
  assign n11367 = ~n11363 & ~n11364;
  assign n11368 = ~n11366_1 & n11367;
  assign n11369 = n11366_1 & ~n11367;
  assign n11370 = ~n11368 & ~n11369;
  assign n11371_1 = n11346_1 & ~n11370;
  assign n11372 = ~n11346_1 & n11370;
  assign n11373 = ~n11371_1 & ~n11372;
  assign n11374 = n11345 & ~n11373;
  assign n11375 = ~n11346_1 & ~n11370;
  assign n11376_1 = ~n11345 & n11375;
  assign n11377 = ~n11345 & n11346_1;
  assign n11378 = n11370 & n11377;
  assign n11379 = ~n11374 & ~n11376_1;
  assign n11380 = ~n11378 & n11379;
  assign n11381_1 = n11343 & ~n11380;
  assign n11382 = ~n11343 & n11380;
  assign n11383 = ~n11381_1 & ~n11382;
  assign n11384 = n11342 & ~n11383;
  assign n11385 = n11343 & n11380;
  assign n11386_1 = ~n11343 & ~n11380;
  assign n11387 = ~n11385 & ~n11386_1;
  assign n11388 = ~n11342 & ~n11387;
  assign n11389 = ~n11384 & ~n11388;
  assign n11390 = ~n10164 & ~n10337;
  assign n11391_1 = ~n11177 & ~n11221_1;
  assign n11392 = ~n11220 & ~n11391_1;
  assign n11393 = n11390 & ~n11392;
  assign n11394 = ~n11390 & n11392;
  assign n11395 = ~n11393 & ~n11394;
  assign n11396_1 = n11389 & ~n11395;
  assign n11397 = ~n11390 & ~n11392;
  assign n11398 = ~n11389 & n11397;
  assign n11399 = ~n11389 & n11390;
  assign n11400 = n11392 & n11399;
  assign n11401_1 = ~n11396_1 & ~n11398;
  assign n11402 = ~n11400 & n11401_1;
  assign n11403 = n11339 & ~n11402;
  assign n11404 = ~n11339 & n11402;
  assign n11405 = ~n11403 & ~n11404;
  assign n11406_1 = n11338 & ~n11405;
  assign n11407 = n11339 & n11402;
  assign n11408 = ~n11339 & ~n11402;
  assign n11409 = ~n11407 & ~n11408;
  assign n11410 = ~n11338 & ~n11409;
  assign n11411_1 = ~n11406_1 & ~n11410;
  assign n11412 = n11335 & ~n11411_1;
  assign n11413 = ~n11335 & n11411_1;
  assign n11414 = ~n11412 & ~n11413;
  assign n11415 = n11334 & ~n11414;
  assign n11416_1 = ~n11335 & ~n11411_1;
  assign n11417 = ~n11334 & n11416_1;
  assign n11418 = ~n11334 & n11335;
  assign n11419 = n11411_1 & n11418;
  assign n11420 = ~n11415 & ~n11417;
  assign n11421_1 = ~n11419 & n11420;
  assign n11422 = n11332 & ~n11421_1;
  assign n11423 = ~n11332 & n11421_1;
  assign n11424 = ~n11422 & ~n11423;
  assign n11425 = n11331_1 & ~n11424;
  assign n11426_1 = n11332 & n11421_1;
  assign n11427 = ~n11332 & ~n11421_1;
  assign n11428 = ~n11426_1 & ~n11427;
  assign n11429 = ~n11331_1 & ~n11428;
  assign n11430 = ~n11425 & ~n11429;
  assign n11431_1 = n11328 & ~n11430;
  assign n11432 = ~n11328 & n11430;
  assign n11433 = ~n11431_1 & ~n11432;
  assign n11434 = n11327 & ~n11433;
  assign n11435 = ~n11328 & ~n11430;
  assign n11436_1 = ~n11327 & n11435;
  assign n11437 = ~n11327 & n11328;
  assign n11438 = n11430 & n11437;
  assign n11439 = ~n11434 & ~n11436_1;
  assign n11440 = ~n11438 & n11439;
  assign n11441_1 = n11325 & ~n11440;
  assign n11442 = ~n11325 & n11440;
  assign n11443 = ~n11441_1 & ~n11442;
  assign n11444 = n11324 & ~n11443;
  assign n11445 = n11325 & n11440;
  assign n11446_1 = ~n11325 & ~n11440;
  assign n11447 = ~n11445 & ~n11446_1;
  assign n11448 = ~n11324 & ~n11447;
  assign n11449 = ~n11444 & ~n11448;
  assign n11450 = n11321_1 & ~n11449;
  assign n11451_1 = ~n11321_1 & n11449;
  assign n11452 = ~n11450 & ~n11451_1;
  assign n11453 = n11320 & ~n11452;
  assign n11454 = ~n11321_1 & ~n11449;
  assign n11455 = ~n11320 & n11454;
  assign n11456_1 = ~n11320 & n11321_1;
  assign n11457 = n11449 & n11456_1;
  assign n11458 = ~n11453 & ~n11455;
  assign n11459 = ~n11457 & n11458;
  assign n11460 = n11318 & ~n11459;
  assign n11461_1 = ~n11318 & n11459;
  assign n11462 = ~n11460 & ~n11461_1;
  assign n11463 = n11317 & ~n11462;
  assign n11464 = n11318 & n11459;
  assign n11465 = ~n11318 & ~n11459;
  assign n11466_1 = ~n11464 & ~n11465;
  assign n11467 = ~n11317 & ~n11466_1;
  assign n11468 = ~n11463 & ~n11467;
  assign n11469 = n11314 & ~n11468;
  assign n11470 = ~n11314 & n11468;
  assign n11471_1 = ~n11469 & ~n11470;
  assign n11472 = n11313 & ~n11471_1;
  assign n11473 = ~n11314 & ~n11468;
  assign n11474 = ~n11313 & n11473;
  assign n11475 = ~n11313 & n11314;
  assign n11476_1 = n11468 & n11475;
  assign n11477 = ~n11472 & ~n11474;
  assign n11478 = ~n11476_1 & n11477;
  assign n11479 = n11311_1 & ~n11478;
  assign n11480 = ~n11311_1 & n11478;
  assign n11481_1 = ~n11479 & ~n11480;
  assign n11482 = n11302 & ~n11481_1;
  assign n11483 = n11311_1 & n11478;
  assign n11484 = ~n11311_1 & ~n11478;
  assign n11485 = ~n11483 & ~n11484;
  assign n11486_1 = ~n11302 & ~n11485;
  assign n11487 = ~n11482 & ~n11486_1;
  assign n11488 = P3_ADDR_REG_15_ & P3_WR_REG;
  assign n11489 = P2_P3_ADDRESS_REG_15_ & n10026_1;
  assign n11490 = P2_P2_ADDRESS_REG_15_ & ~n10026_1;
  assign n11491_1 = ~n11489 & ~n11490;
  assign n11492 = n10061_1 & ~n11491_1;
  assign n11493 = P2_P1_ADDRESS_REG_15_ & n10063;
  assign n11494 = ~n11488 & ~n11492;
  assign n11495 = ~n11493 & n11494;
  assign n11496_1 = P4_ADDR_REG_2_ & P4_WR_REG;
  assign n11497 = P1_P3_ADDRESS_REG_2_ & n10072;
  assign n11498 = P1_P2_ADDRESS_REG_2_ & ~n10072;
  assign n11499 = ~n11497 & ~n11498;
  assign n11500 = n10107 & ~n11499;
  assign n11501_1 = P1_P1_ADDRESS_REG_2_ & n10109;
  assign n11502 = ~n11496_1 & ~n11500;
  assign n11503 = ~n11501_1 & n11502;
  assign n11504 = ~n11495 & ~n11503;
  assign n11505 = ~n11310 & ~n11503;
  assign n11506_1 = ~n10113 & n11298;
  assign n11507 = ~n11299 & ~n11506_1;
  assign n11508 = n11146_1 & ~n11507;
  assign n11509 = ~n10113 & ~n11298;
  assign n11510 = ~n11146_1 & n11509;
  assign n11511_1 = n11147 & n11298;
  assign n11512 = ~n11508 & ~n11510;
  assign n11513 = ~n11511_1 & n11512;
  assign n11514 = n11505 & n11513;
  assign n11515 = ~n11505 & ~n11513;
  assign n11516_1 = ~n10066_1 & ~n11503;
  assign n11517 = ~n11011_1 & n11140;
  assign n11518 = ~n11141_1 & ~n11517;
  assign n11519 = n11132 & ~n11518;
  assign n11520 = ~n11011_1 & ~n11140;
  assign n11521_1 = ~n11132 & n11520;
  assign n11522 = n11133 & n11140;
  assign n11523 = ~n11519 & ~n11521_1;
  assign n11524 = ~n11522 & n11523;
  assign n11525 = ~n10121_1 & ~n11503;
  assign n11526_1 = n11524 & n11525;
  assign n11527 = ~n11524 & ~n11525;
  assign n11528 = ~n10869 & ~n11503;
  assign n11529 = ~n10130 & ~n11503;
  assign n11530 = ~n10642 & ~n11503;
  assign n11531_1 = ~n11035 & n11112;
  assign n11532 = ~n11113 & ~n11531_1;
  assign n11533 = n11104 & ~n11532;
  assign n11534 = ~n11035 & ~n11112;
  assign n11535 = ~n11104 & n11534;
  assign n11536_1 = n11105 & n11112;
  assign n11537 = ~n11533 & ~n11535;
  assign n11538 = ~n11536_1 & n11537;
  assign n11539 = ~n10147 & ~n11503;
  assign n11540 = n11538 & n11539;
  assign n11541_1 = ~n11538 & ~n11539;
  assign n11542 = ~n10472 & ~n11503;
  assign n11543 = ~n10383 & ~n11503;
  assign n11544 = ~n10164 & ~n11503;
  assign n11545 = n11048 & ~n11085;
  assign n11546_1 = ~n11048 & n11085;
  assign n11547 = ~n11545 & ~n11546_1;
  assign n11548 = n11076_1 & ~n11547;
  assign n11549 = ~n11048 & ~n11085;
  assign n11550 = ~n11076_1 & n11549;
  assign n11551_1 = n11077 & n11085;
  assign n11552 = ~n11548 & ~n11550;
  assign n11553 = ~n11551_1 & n11552;
  assign n11554 = n11544 & ~n11553;
  assign n11555 = ~n11049 & n11057;
  assign n11556_1 = ~n11058 & ~n11555;
  assign n11557 = n11072 & ~n11556_1;
  assign n11558 = ~n11049 & ~n11057;
  assign n11559 = ~n11072 & n11558;
  assign n11560 = n11057 & n11073;
  assign n11561_1 = ~n11557 & ~n11559;
  assign n11562 = ~n11560 & n11561_1;
  assign n11563 = ~n10181_1 & ~n11503;
  assign n11564 = n11562 & n11563;
  assign n11565 = ~n11562 & ~n11563;
  assign n11566_1 = ~n10257 & ~n11503;
  assign n11567 = ~n10198 & ~n11503;
  assign n11568 = n10112 & ~n10225;
  assign n11569 = ~n10238 & ~n11568;
  assign n11570 = ~n10138 & ~n11569;
  assign n11571_1 = n10138 & ~n10216_1;
  assign n11572 = ~n10226_1 & ~n11571_1;
  assign n11573 = ~n10112 & ~n11572;
  assign n11574 = ~n11570 & ~n11573;
  assign n11575 = n11567 & ~n11574;
  assign n11576_1 = ~n10112 & ~n11503;
  assign n11577 = n10244 & n11576_1;
  assign n11578 = ~n11567 & n11574;
  assign n11579 = n11577 & ~n11578;
  assign n11580 = ~n11575 & ~n11579;
  assign n11581_1 = n11566_1 & ~n11580;
  assign n11582 = n11061_1 & ~n11070;
  assign n11583 = ~n11061_1 & n11070;
  assign n11584 = ~n11582 & ~n11583;
  assign n11585 = ~n11060 & n11584;
  assign n11586_1 = n11060 & n11583;
  assign n11587 = n11062 & ~n11070;
  assign n11588 = ~n11585 & ~n11586_1;
  assign n11589 = ~n11587 & n11588;
  assign n11590 = n11566_1 & ~n11589;
  assign n11591_1 = ~n11580 & ~n11589;
  assign n11592 = ~n11581_1 & ~n11590;
  assign n11593 = ~n11591_1 & n11592;
  assign n11594 = ~n11565 & ~n11593;
  assign n11595 = ~n11564 & ~n11594;
  assign n11596_1 = n11544 & ~n11595;
  assign n11597 = ~n11553 & ~n11595;
  assign n11598 = ~n11554 & ~n11596_1;
  assign n11599 = ~n11597 & n11598;
  assign n11600 = n11543 & ~n11599;
  assign n11601_1 = ~n11037 & n11046_1;
  assign n11602 = ~n11047 & ~n11601_1;
  assign n11603 = n11088 & ~n11602;
  assign n11604 = ~n11037 & ~n11046_1;
  assign n11605 = ~n11088 & n11604;
  assign n11606_1 = n11046_1 & n11089;
  assign n11607 = ~n11603 & ~n11605;
  assign n11608 = ~n11606_1 & n11607;
  assign n11609 = ~n11543 & n11599;
  assign n11610 = n11608 & ~n11609;
  assign n11611_1 = ~n11600 & ~n11610;
  assign n11612 = n11542 & ~n11611_1;
  assign n11613 = n11036_1 & ~n11101_1;
  assign n11614 = ~n11036_1 & n11101_1;
  assign n11615 = ~n11613 & ~n11614;
  assign n11616_1 = n11092 & ~n11615;
  assign n11617 = ~n11036_1 & ~n11101_1;
  assign n11618 = ~n11092 & n11617;
  assign n11619 = n11093 & n11101_1;
  assign n11620 = ~n11616_1 & ~n11618;
  assign n11621_1 = ~n11619 & n11620;
  assign n11622 = n11542 & ~n11621_1;
  assign n11623 = ~n11611_1 & ~n11621_1;
  assign n11624 = ~n11612 & ~n11622;
  assign n11625 = ~n11623 & n11624;
  assign n11626_1 = ~n11541_1 & ~n11625;
  assign n11627 = ~n11540 & ~n11626_1;
  assign n11628 = n11530 & ~n11627;
  assign n11629 = ~n11031_1 & n11032;
  assign n11630 = n11031_1 & ~n11032;
  assign n11631_1 = ~n11629 & ~n11630;
  assign n11632 = n11116_1 & ~n11631_1;
  assign n11633 = ~n11033 & ~n11034;
  assign n11634 = ~n11116_1 & ~n11633;
  assign n11635 = ~n11632 & ~n11634;
  assign n11636_1 = n11530 & ~n11635;
  assign n11637 = ~n11627 & ~n11635;
  assign n11638 = ~n11628 & ~n11636_1;
  assign n11639 = ~n11637 & n11638;
  assign n11640 = n11529 & ~n11639;
  assign n11641_1 = ~n11023 & n11126_1;
  assign n11642 = ~n11127 & ~n11641_1;
  assign n11643 = n11118 & ~n11642;
  assign n11644 = ~n11023 & ~n11126_1;
  assign n11645 = ~n11118 & n11644;
  assign n11646_1 = n11119 & n11126_1;
  assign n11647 = ~n11643 & ~n11645;
  assign n11648 = ~n11646_1 & n11647;
  assign n11649 = ~n11529 & n11639;
  assign n11650 = n11648 & ~n11649;
  assign n11651_1 = ~n11640 & ~n11650;
  assign n11652 = n11528 & ~n11651_1;
  assign n11653 = ~n11019 & n11020;
  assign n11654 = n11019 & ~n11020;
  assign n11655 = ~n11653 & ~n11654;
  assign n11656_1 = n11130 & ~n11655;
  assign n11657 = ~n11021_1 & ~n11022;
  assign n11658 = ~n11130 & ~n11657;
  assign n11659 = ~n11656_1 & ~n11658;
  assign n11660 = n11528 & ~n11659;
  assign n11661_1 = ~n11651_1 & ~n11659;
  assign n11662 = ~n11652 & ~n11660;
  assign n11663 = ~n11661_1 & n11662;
  assign n11664 = ~n11527 & ~n11663;
  assign n11665 = ~n11526_1 & ~n11664;
  assign n11666_1 = n11516_1 & ~n11665;
  assign n11667 = n10122 & ~n11008;
  assign n11668 = ~n10122 & n11008;
  assign n11669 = ~n11667 & ~n11668;
  assign n11670 = n11144 & ~n11669;
  assign n11671_1 = ~n11009 & ~n11010;
  assign n11672 = ~n11144 & ~n11671_1;
  assign n11673 = ~n11670 & ~n11672;
  assign n11674 = n11516_1 & ~n11673;
  assign n11675 = ~n11665 & ~n11673;
  assign n11676_1 = ~n11666_1 & ~n11674;
  assign n11677 = ~n11675 & n11676_1;
  assign n11678 = ~n11515 & ~n11677;
  assign n11679 = ~n11514 & ~n11678;
  assign n11680 = n11504 & ~n11679;
  assign n11681_1 = ~n11504 & n11679;
  assign n11682 = ~n11680 & ~n11681_1;
  assign n11683 = n11487 & ~n11682;
  assign n11684 = ~n11504 & ~n11679;
  assign n11685 = ~n11487 & n11684;
  assign n11686_1 = ~n11487 & n11504;
  assign n11687 = n11679 & n11686_1;
  assign n11688 = ~n11683 & ~n11685;
  assign n11689 = ~n11687 & n11688;
  assign n11690 = P3_ADDR_REG_16_ & P3_WR_REG;
  assign n11691_1 = P2_P3_ADDRESS_REG_16_ & n10026_1;
  assign n11692 = P2_P2_ADDRESS_REG_16_ & ~n10026_1;
  assign n11693 = ~n11691_1 & ~n11692;
  assign n11694 = n10061_1 & ~n11693;
  assign n11695 = P2_P1_ADDRESS_REG_16_ & n10063;
  assign n11696_1 = ~n11690 & ~n11694;
  assign n11697 = ~n11695 & n11696_1;
  assign n11698 = P4_ADDR_REG_1_ & P4_WR_REG;
  assign n11699 = P1_P1_ADDRESS_REG_1_ & n10106_1;
  assign n11700 = P1_P3_ADDRESS_REG_1_ & n10072;
  assign n11701_1 = P1_P2_ADDRESS_REG_1_ & ~n10072;
  assign n11702 = ~n11700 & ~n11701_1;
  assign n11703 = ~n10106_1 & ~n11702;
  assign n11704 = ~n11699 & ~n11703;
  assign n11705 = ~P4_WR_REG & ~n11704;
  assign n11706_1 = ~n11698 & ~n11705;
  assign n11707 = ~n11697 & ~n11706_1;
  assign n11708 = n11689 & n11707;
  assign n11709 = ~n11689 & ~n11707;
  assign n11710 = ~n11495 & ~n11706_1;
  assign n11711_1 = ~n11310 & ~n11706_1;
  assign n11712 = ~n10066_1 & ~n11706_1;
  assign n11713 = ~n11524 & n11525;
  assign n11714 = n11524 & ~n11525;
  assign n11715 = ~n11713 & ~n11714;
  assign n11716_1 = n11663 & ~n11715;
  assign n11717 = ~n11526_1 & ~n11527;
  assign n11718 = ~n11663 & ~n11717;
  assign n11719 = ~n11716_1 & ~n11718;
  assign n11720 = n11712 & ~n11719;
  assign n11721_1 = ~n11528 & n11659;
  assign n11722 = ~n11660 & ~n11721_1;
  assign n11723 = n11651_1 & ~n11722;
  assign n11724 = ~n11528 & ~n11659;
  assign n11725 = ~n11651_1 & n11724;
  assign n11726_1 = n11652 & n11659;
  assign n11727 = ~n11723 & ~n11725;
  assign n11728 = ~n11726_1 & n11727;
  assign n11729 = ~n10121_1 & ~n11706_1;
  assign n11730 = n11728 & n11729;
  assign n11731_1 = ~n11728 & ~n11729;
  assign n11732 = ~n10869 & ~n11706_1;
  assign n11733 = ~n10130 & ~n11706_1;
  assign n11734 = ~n10642 & ~n11706_1;
  assign n11735 = ~n10147 & ~n11706_1;
  assign n11736_1 = ~n10472 & ~n11706_1;
  assign n11737 = ~n11544 & n11595;
  assign n11738 = ~n11596_1 & ~n11737;
  assign n11739 = n11553 & ~n11738;
  assign n11740 = ~n11544 & ~n11595;
  assign n11741_1 = ~n11553 & n11740;
  assign n11742 = n11554 & n11595;
  assign n11743 = ~n11739 & ~n11741_1;
  assign n11744 = ~n11742 & n11743;
  assign n11745 = ~n10383 & ~n11706_1;
  assign n11746_1 = n11744 & n11745;
  assign n11747 = ~n11744 & ~n11745;
  assign n11748 = ~n10164 & ~n11706_1;
  assign n11749 = ~n11566_1 & n11589;
  assign n11750 = ~n11590 & ~n11749;
  assign n11751_1 = n11580 & ~n11750;
  assign n11752 = ~n11566_1 & ~n11589;
  assign n11753 = ~n11580 & n11752;
  assign n11754 = n11581_1 & n11589;
  assign n11755 = ~n11751_1 & ~n11753;
  assign n11756_1 = ~n11754 & n11755;
  assign n11757 = ~n10181_1 & ~n11706_1;
  assign n11758 = n11756_1 & n11757;
  assign n11759 = ~n11756_1 & ~n11757;
  assign n11760 = ~n10257 & ~n11706_1;
  assign n11761_1 = ~n10198 & ~n11706_1;
  assign n11762 = ~n10225 & n11503;
  assign n11763 = ~n10238 & ~n11762;
  assign n11764 = ~n10112 & ~n11763;
  assign n11765 = n10112 & ~n10216_1;
  assign n11766_1 = ~n10226_1 & ~n11765;
  assign n11767 = ~n11503 & ~n11766_1;
  assign n11768 = ~n11764 & ~n11767;
  assign n11769 = n11761_1 & ~n11768;
  assign n11770 = ~n11503 & ~n11706_1;
  assign n11771_1 = n10244 & n11770;
  assign n11772 = ~n11761_1 & n11768;
  assign n11773 = n11771_1 & ~n11772;
  assign n11774 = ~n11769 & ~n11773;
  assign n11775 = n11760 & ~n11774;
  assign n11776_1 = ~n11575 & ~n11578;
  assign n11777 = ~n11577 & n11776_1;
  assign n11778 = n11577 & ~n11776_1;
  assign n11779 = ~n11777 & ~n11778;
  assign n11780 = n11760 & ~n11779;
  assign n11781_1 = ~n11774 & ~n11779;
  assign n11782 = ~n11775 & ~n11780;
  assign n11783 = ~n11781_1 & n11782;
  assign n11784 = ~n11759 & ~n11783;
  assign n11785 = ~n11758 & ~n11784;
  assign n11786_1 = n11748 & ~n11785;
  assign n11787 = ~n11562 & n11563;
  assign n11788 = n11562 & ~n11563;
  assign n11789 = ~n11787 & ~n11788;
  assign n11790 = n11593 & ~n11789;
  assign n11791_1 = ~n11564 & ~n11565;
  assign n11792 = ~n11593 & ~n11791_1;
  assign n11793 = ~n11790 & ~n11792;
  assign n11794 = n11748 & ~n11793;
  assign n11795 = ~n11785 & ~n11793;
  assign n11796_1 = ~n11786_1 & ~n11794;
  assign n11797 = ~n11795 & n11796_1;
  assign n11798 = ~n11747 & ~n11797;
  assign n11799 = ~n11746_1 & ~n11798;
  assign n11800 = n11736_1 & ~n11799;
  assign n11801_1 = ~n11600 & ~n11609;
  assign n11802 = ~n11608 & n11801_1;
  assign n11803 = n11608 & ~n11801_1;
  assign n11804 = ~n11802 & ~n11803;
  assign n11805 = n11736_1 & ~n11804;
  assign n11806_1 = ~n11799 & ~n11804;
  assign n11807 = ~n11800 & ~n11805;
  assign n11808 = ~n11806_1 & n11807;
  assign n11809 = n11735 & ~n11808;
  assign n11810 = ~n11542 & n11611_1;
  assign n11811_1 = ~n11612 & ~n11810;
  assign n11812 = n11621_1 & ~n11811_1;
  assign n11813 = ~n11542 & ~n11611_1;
  assign n11814 = ~n11621_1 & n11813;
  assign n11815 = n11611_1 & n11622;
  assign n11816_1 = ~n11812 & ~n11814;
  assign n11817 = ~n11815 & n11816_1;
  assign n11818 = ~n11735 & n11808;
  assign n11819 = n11817 & ~n11818;
  assign n11820 = ~n11809 & ~n11819;
  assign n11821_1 = n11734 & ~n11820;
  assign n11822 = ~n11538 & n11539;
  assign n11823 = n11538 & ~n11539;
  assign n11824 = ~n11822 & ~n11823;
  assign n11825 = n11625 & ~n11824;
  assign n11826_1 = ~n11540 & ~n11541_1;
  assign n11827 = ~n11625 & ~n11826_1;
  assign n11828 = ~n11825 & ~n11827;
  assign n11829 = n11734 & ~n11828;
  assign n11830 = ~n11820 & ~n11828;
  assign n11831_1 = ~n11821_1 & ~n11829;
  assign n11832 = ~n11830 & n11831_1;
  assign n11833 = n11733 & ~n11832;
  assign n11834 = ~n11530 & n11635;
  assign n11835 = ~n11636_1 & ~n11834;
  assign n11836_1 = n11627 & ~n11835;
  assign n11837 = ~n11530 & ~n11635;
  assign n11838 = ~n11627 & n11837;
  assign n11839 = n11628 & n11635;
  assign n11840 = ~n11836_1 & ~n11838;
  assign n11841_1 = ~n11839 & n11840;
  assign n11842 = ~n11733 & n11832;
  assign n11843 = n11841_1 & ~n11842;
  assign n11844 = ~n11833 & ~n11843;
  assign n11845 = n11732 & ~n11844;
  assign n11846_1 = ~n11640 & ~n11649;
  assign n11847 = ~n11648 & n11846_1;
  assign n11848 = n11648 & ~n11846_1;
  assign n11849 = ~n11847 & ~n11848;
  assign n11850 = n11732 & ~n11849;
  assign n11851_1 = ~n11844 & ~n11849;
  assign n11852 = ~n11845 & ~n11850;
  assign n11853 = ~n11851_1 & n11852;
  assign n11854 = ~n11731_1 & ~n11853;
  assign n11855 = ~n11730 & ~n11854;
  assign n11856_1 = n11712 & ~n11855;
  assign n11857 = ~n11719 & ~n11855;
  assign n11858 = ~n11720 & ~n11856_1;
  assign n11859 = ~n11857 & n11858;
  assign n11860 = n11711_1 & ~n11859;
  assign n11861_1 = ~n11516_1 & n11673;
  assign n11862 = ~n11674 & ~n11861_1;
  assign n11863 = n11665 & ~n11862;
  assign n11864 = ~n11516_1 & ~n11673;
  assign n11865 = ~n11665 & n11864;
  assign n11866_1 = n11666_1 & n11673;
  assign n11867 = ~n11863 & ~n11865;
  assign n11868 = ~n11866_1 & n11867;
  assign n11869 = ~n11711_1 & n11859;
  assign n11870 = n11868 & ~n11869;
  assign n11871_1 = ~n11860 & ~n11870;
  assign n11872 = n11710 & ~n11871_1;
  assign n11873 = n11505 & ~n11513;
  assign n11874 = ~n11505 & n11513;
  assign n11875 = ~n11873 & ~n11874;
  assign n11876_1 = n11677 & ~n11875;
  assign n11877 = ~n11514 & ~n11515;
  assign n11878 = ~n11677 & ~n11877;
  assign n11879 = ~n11876_1 & ~n11878;
  assign n11880 = n11710 & ~n11879;
  assign n11881_1 = ~n11871_1 & ~n11879;
  assign n11882 = ~n11872 & ~n11880;
  assign n11883 = ~n11881_1 & n11882;
  assign n11884 = ~n11709 & ~n11883;
  assign n11885 = ~n11708 & ~n11884;
  assign n11886_1 = P3_ADDR_REG_17_ & P3_WR_REG;
  assign n11887 = P2_P3_ADDRESS_REG_17_ & n10026_1;
  assign n11888 = P2_P2_ADDRESS_REG_17_ & ~n10026_1;
  assign n11889 = ~n11887 & ~n11888;
  assign n11890 = n10061_1 & ~n11889;
  assign n11891_1 = P2_P1_ADDRESS_REG_17_ & n10063;
  assign n11892 = ~n11886_1 & ~n11890;
  assign n11893 = ~n11891_1 & n11892;
  assign n11894 = ~n11706_1 & ~n11893;
  assign n11895 = P3_ADDR_REG_18_ & P3_WR_REG;
  assign n11896_1 = P2_P3_ADDRESS_REG_18_ & n10026_1;
  assign n11897 = P2_P2_ADDRESS_REG_18_ & ~n10026_1;
  assign n11898 = ~n11896_1 & ~n11897;
  assign n11899 = n10061_1 & ~n11898;
  assign n11900 = P2_P1_ADDRESS_REG_18_ & n10063;
  assign n11901_1 = ~n11895 & ~n11899;
  assign n11902 = ~n11900 & n11901_1;
  assign n11903 = P4_ADDR_REG_0_ & P4_WR_REG;
  assign n11904 = P1_P1_ADDRESS_REG_0_ & n10106_1;
  assign n11905 = P1_P3_ADDRESS_REG_0_ & n10072;
  assign n11906_1 = P1_P2_ADDRESS_REG_0_ & ~n10072;
  assign n11907 = ~n11905 & ~n11906_1;
  assign n11908 = ~n10106_1 & ~n11907;
  assign n11909 = ~n11904 & ~n11908;
  assign n11910 = ~P4_WR_REG & ~n11909;
  assign n11911_1 = ~n11903 & ~n11910;
  assign n11912 = ~n11902 & ~n11911_1;
  assign n11913 = n11894 & ~n11912;
  assign n11914 = ~n11894 & n11912;
  assign n11915 = ~n11913 & ~n11914;
  assign n11916_1 = ~n11487 & ~n11679;
  assign n11917 = ~n11680 & ~n11686_1;
  assign n11918 = ~n11916_1 & n11917;
  assign n11919 = ~n11302 & ~n11484;
  assign n11920 = ~n11483 & ~n11919;
  assign n11921_1 = ~n11503 & ~n11697;
  assign n11922 = ~n10112 & ~n11495;
  assign n11923 = n11921_1 & ~n11922;
  assign n11924 = ~n11921_1 & n11922;
  assign n11925 = ~n11923 & ~n11924;
  assign n11926_1 = ~n11313 & ~n11468;
  assign n11927 = ~n11469 & ~n11475;
  assign n11928 = ~n11926_1 & n11927;
  assign n11929 = ~n11320 & ~n11449;
  assign n11930 = ~n11450 & ~n11456_1;
  assign n11931_1 = ~n11929 & n11930;
  assign n11932 = ~n10066_1 & ~n10155;
  assign n11933 = ~n11324 & ~n11446_1;
  assign n11934 = ~n11445 & ~n11933;
  assign n11935 = ~n11327 & ~n11430;
  assign n11936_1 = ~n11431_1 & ~n11437;
  assign n11937 = ~n11935 & n11936_1;
  assign n11938 = ~n11331_1 & ~n11427;
  assign n11939 = ~n11426_1 & ~n11938;
  assign n11940 = ~n11334 & ~n11411_1;
  assign n11941_1 = ~n11412 & ~n11418;
  assign n11942 = ~n11940 & n11941_1;
  assign n11943 = ~n10207 & ~n10642;
  assign n11944 = ~n10147 & ~n10234;
  assign n11945 = n11943 & ~n11944;
  assign n11946_1 = ~n11943 & n11944;
  assign n11947 = ~n11945 & ~n11946_1;
  assign n11948 = ~n11338 & ~n11408;
  assign n11949 = ~n11407 & ~n11948;
  assign n11950 = ~n11342 & ~n11386_1;
  assign n11951_1 = ~n11385 & ~n11950;
  assign n11952 = ~n10337 & ~n10383;
  assign n11953 = ~n11345 & ~n11370;
  assign n11954 = ~n11371_1 & ~n11377;
  assign n11955 = ~n11953 & n11954;
  assign n11956_1 = ~n11364 & n11366_1;
  assign n11957 = ~n11363 & ~n11956_1;
  assign n11958 = ~n11190 & ~n11355;
  assign n11959 = n10244 & n11958;
  assign n11960 = P4_ADDR_REG_18_ & P4_WR_REG;
  assign n11961_1 = P1_P3_ADDRESS_REG_18_ & n10072;
  assign n11962 = P1_P2_ADDRESS_REG_18_ & ~n10072;
  assign n11963 = ~n11961_1 & ~n11962;
  assign n11964 = n10107 & ~n11963;
  assign n11965 = P1_P1_ADDRESS_REG_18_ & n10109;
  assign n11966_1 = ~n11960 & ~n11964;
  assign n11967 = ~n11965 & n11966_1;
  assign n11968 = ~n10216_1 & n11967;
  assign n11969 = ~n10226_1 & ~n11968;
  assign n11970 = ~n11355 & ~n11969;
  assign n11971_1 = ~n10225 & n11355;
  assign n11972 = ~n10238 & ~n11971_1;
  assign n11973 = ~n11967 & ~n11972;
  assign n11974 = ~n11970 & ~n11973;
  assign n11975 = n10198 & n11974;
  assign n11976_1 = ~n10198 & ~n11974;
  assign n11977 = ~n11975 & ~n11976_1;
  assign n11978 = n11959 & ~n11977;
  assign n11979 = ~n10198 & ~n11190;
  assign n11980 = ~n11974 & n11979;
  assign n11981_1 = n11974 & ~n11979;
  assign n11982 = ~n11980 & ~n11981_1;
  assign n11983 = ~n11959 & n11982;
  assign n11984 = ~n11978 & ~n11983;
  assign n11985 = ~n10257 & ~n10907;
  assign n11986_1 = ~n11984 & ~n11985;
  assign n11987 = n11984 & n11985;
  assign n11988 = ~n11986_1 & ~n11987;
  assign n11989 = n11957 & n11988;
  assign n11990 = ~n11957 & ~n11988;
  assign n11991_1 = ~n11989 & ~n11990;
  assign n11992 = n11955 & n11991_1;
  assign n11993 = ~n11955 & ~n11991_1;
  assign n11994 = ~n11992 & ~n11993;
  assign n11995 = ~n10181_1 & ~n10677;
  assign n11996_1 = ~n10164 & ~n10400;
  assign n11997 = n11995 & ~n11996_1;
  assign n11998 = ~n11995 & n11996_1;
  assign n11999 = ~n11997 & ~n11998;
  assign n12000 = ~n11994 & n11999;
  assign n12001_1 = n11994 & ~n11999;
  assign n12002 = ~n12000 & ~n12001_1;
  assign n12003 = n11952 & n12002;
  assign n12004 = ~n11952 & ~n12002;
  assign n12005 = ~n12003 & ~n12004;
  assign n12006_1 = n11951_1 & n12005;
  assign n12007 = ~n11951_1 & ~n12005;
  assign n12008 = ~n12006_1 & ~n12007;
  assign n12009 = ~n10267 & ~n10472;
  assign n12010 = ~n12008 & ~n12009;
  assign n12011_1 = n12008 & n12009;
  assign n12012 = ~n12010 & ~n12011_1;
  assign n12013 = ~n11389 & ~n11392;
  assign n12014 = ~n11393 & ~n11399;
  assign n12015 = ~n12013 & n12014;
  assign n12016_1 = ~n12012 & ~n12015;
  assign n12017 = n12012 & n12015;
  assign n12018 = ~n12016_1 & ~n12017;
  assign n12019 = n11949 & n12018;
  assign n12020 = ~n11949 & ~n12018;
  assign n12021_1 = ~n12019 & ~n12020;
  assign n12022 = ~n11947 & n12021_1;
  assign n12023 = n11947 & ~n12021_1;
  assign n12024 = ~n12022 & ~n12023;
  assign n12025 = n11942 & n12024;
  assign n12026_1 = ~n11942 & ~n12024;
  assign n12027 = ~n12025 & ~n12026_1;
  assign n12028 = n11939 & n12027;
  assign n12029 = ~n11939 & ~n12027;
  assign n12030 = ~n12028 & ~n12029;
  assign n12031_1 = ~n10130 & ~n10190;
  assign n12032 = ~n12030 & ~n12031_1;
  assign n12033 = n12030 & n12031_1;
  assign n12034 = ~n12032 & ~n12033;
  assign n12035 = n11937 & n12034;
  assign n12036_1 = ~n11937 & ~n12034;
  assign n12037 = ~n12035 & ~n12036_1;
  assign n12038 = n11934 & n12037;
  assign n12039 = ~n11934 & ~n12037;
  assign n12040 = ~n12038 & ~n12039;
  assign n12041_1 = ~n10172 & ~n10869;
  assign n12042 = ~n10121_1 & ~n10464;
  assign n12043 = n12041_1 & ~n12042;
  assign n12044 = ~n12041_1 & n12042;
  assign n12045 = ~n12043 & ~n12044;
  assign n12046_1 = ~n12040 & n12045;
  assign n12047 = n12040 & ~n12045;
  assign n12048 = ~n12046_1 & ~n12047;
  assign n12049 = n11932 & n12048;
  assign n12050 = ~n11932 & ~n12048;
  assign n12051_1 = ~n12049 & ~n12050;
  assign n12052 = n11931_1 & n12051_1;
  assign n12053 = ~n11931_1 & ~n12051_1;
  assign n12054 = ~n12052 & ~n12053;
  assign n12055 = ~n10138 & ~n11310;
  assign n12056_1 = ~n12054 & ~n12055;
  assign n12057 = n12054 & n12055;
  assign n12058 = ~n12056_1 & ~n12057;
  assign n12059 = ~n11317 & ~n11465;
  assign n12060 = ~n11464 & ~n12059;
  assign n12061_1 = ~n12058 & ~n12060;
  assign n12062 = n12058 & n12060;
  assign n12063 = ~n12061_1 & ~n12062;
  assign n12064 = n11928 & n12063;
  assign n12065 = ~n11928 & ~n12063;
  assign n12066_1 = ~n12064 & ~n12065;
  assign n12067 = ~n11925 & n12066_1;
  assign n12068 = n11925 & ~n12066_1;
  assign n12069 = ~n12067 & ~n12068;
  assign n12070 = n11920 & n12069;
  assign n12071_1 = ~n11920 & ~n12069;
  assign n12072 = ~n12070 & ~n12071_1;
  assign n12073 = n11918 & n12072;
  assign n12074 = ~n11918 & ~n12072;
  assign n12075 = ~n12073 & ~n12074;
  assign n12076_1 = ~n11915 & n12075;
  assign n12077 = n11915 & ~n12075;
  assign n12078 = ~n12076_1 & ~n12077;
  assign n12079 = n11885 & n12078;
  assign n12080 = ~n11885 & ~n12078;
  assign n12081_1 = ~n12079 & ~n12080;
  assign n12082 = ~n11893 & ~n11911_1;
  assign n12083 = ~n11697 & ~n11911_1;
  assign n12084 = ~n11495 & ~n11911_1;
  assign n12085 = ~n11860 & ~n11869;
  assign n12086_1 = ~n11868 & n12085;
  assign n12087 = n11868 & ~n12085;
  assign n12088 = ~n12086_1 & ~n12087;
  assign n12089 = n12084 & ~n12088;
  assign n12090 = ~n12084 & n12088;
  assign n12091_1 = ~n11310 & ~n11911_1;
  assign n12092 = ~n10066_1 & ~n11911_1;
  assign n12093 = ~n11728 & n11729;
  assign n12094 = n11728 & ~n11729;
  assign n12095 = ~n12093 & ~n12094;
  assign n12096_1 = n11853 & ~n12095;
  assign n12097 = ~n11730 & ~n11731_1;
  assign n12098 = ~n11853 & ~n12097;
  assign n12099 = ~n12096_1 & ~n12098;
  assign n12100 = n12092 & ~n12099;
  assign n12101_1 = ~n12092 & n12099;
  assign n12102 = ~n11732 & n11849;
  assign n12103 = ~n11850 & ~n12102;
  assign n12104 = n11844 & ~n12103;
  assign n12105 = ~n11732 & ~n11849;
  assign n12106_1 = ~n11844 & n12105;
  assign n12107 = n11845 & n11849;
  assign n12108 = ~n12104 & ~n12106_1;
  assign n12109 = ~n12107 & n12108;
  assign n12110 = ~n10121_1 & ~n11911_1;
  assign n12111_1 = n12109 & n12110;
  assign n12112 = ~n12109 & ~n12110;
  assign n12113 = ~n10869 & ~n11911_1;
  assign n12114 = ~n11833 & ~n11842;
  assign n12115 = ~n11841_1 & n12114;
  assign n12116_1 = n11841_1 & ~n12114;
  assign n12117 = ~n12115 & ~n12116_1;
  assign n12118 = n12113 & ~n12117;
  assign n12119 = ~n12113 & n12117;
  assign n12120 = ~n10130 & ~n11911_1;
  assign n12121_1 = ~n10642 & ~n11911_1;
  assign n12122 = ~n10147 & ~n11911_1;
  assign n12123 = ~n10472 & ~n11911_1;
  assign n12124 = ~n11744 & n11745;
  assign n12125 = n11744 & ~n11745;
  assign n12126_1 = ~n12124 & ~n12125;
  assign n12127 = n11797 & ~n12126_1;
  assign n12128 = ~n11746_1 & ~n11747;
  assign n12129 = ~n11797 & ~n12128;
  assign n12130 = ~n12127 & ~n12129;
  assign n12131_1 = n12123 & ~n12130;
  assign n12132 = ~n12123 & n12130;
  assign n12133 = ~n11748 & n11793;
  assign n12134 = ~n11794 & ~n12133;
  assign n12135 = n11785 & ~n12134;
  assign n12136_1 = ~n11748 & ~n11793;
  assign n12137 = ~n11785 & n12136_1;
  assign n12138 = n11786_1 & n11793;
  assign n12139 = ~n12135 & ~n12137;
  assign n12140 = ~n12138 & n12139;
  assign n12141_1 = ~n10383 & ~n11911_1;
  assign n12142 = n12140 & n12141_1;
  assign n12143 = ~n12140 & ~n12141_1;
  assign n12144 = ~n10164 & ~n11911_1;
  assign n12145 = ~n10181_1 & ~n11911_1;
  assign n12146_1 = ~n10257 & ~n11911_1;
  assign n12147 = ~n11769 & ~n11772;
  assign n12148 = ~n11771_1 & n12147;
  assign n12149 = n11771_1 & ~n12147;
  assign n12150 = ~n12148 & ~n12149;
  assign n12151_1 = n12146_1 & ~n12150;
  assign n12152 = ~n12146_1 & n12150;
  assign MUL_1411_U5 = ~n10225 & ~n11911_1;
  assign n12154 = ~n10216_1 & ~n11706_1;
  assign n12155 = MUL_1411_U5 & n12154;
  assign n12156_1 = ~n10198 & ~n11911_1;
  assign n12157 = n12155 & n12156_1;
  assign n12158 = ~n12155 & ~n12156_1;
  assign n12159 = ~n10216_1 & n11503;
  assign n12160 = ~n10226_1 & ~n12159;
  assign n12161_1 = ~n11706_1 & ~n12160;
  assign n12162 = ~n10225 & n11706_1;
  assign n12163 = ~n10238 & ~n12162;
  assign n12164 = ~n11503 & ~n12163;
  assign n12165 = ~n12161_1 & ~n12164;
  assign n12166_1 = ~n12158 & ~n12165;
  assign n12167 = ~n12157 & ~n12166_1;
  assign n12168 = ~n12152 & ~n12167;
  assign n12169 = ~n12151_1 & ~n12168;
  assign n12170 = n12145 & ~n12169;
  assign n12171_1 = ~n11760 & n11779;
  assign n12172 = ~n11780 & ~n12171_1;
  assign n12173 = n11774 & ~n12172;
  assign n12174 = ~n11760 & ~n11779;
  assign n12175 = ~n11774 & n12174;
  assign n12176_1 = n11775 & n11779;
  assign n12177 = ~n12173 & ~n12175;
  assign n12178 = ~n12176_1 & n12177;
  assign n12179 = ~n12145 & n12169;
  assign n12180 = n12178 & ~n12179;
  assign n12181_1 = ~n12170 & ~n12180;
  assign n12182 = n12144 & ~n12181_1;
  assign n12183 = ~n11756_1 & n11757;
  assign n12184 = n11756_1 & ~n11757;
  assign n12185 = ~n12183 & ~n12184;
  assign n12186_1 = n11783 & ~n12185;
  assign n12187 = ~n11758 & ~n11759;
  assign n12188 = ~n11783 & ~n12187;
  assign n12189 = ~n12186_1 & ~n12188;
  assign n12190 = ~n12144 & n12181_1;
  assign n12191_1 = ~n12189 & ~n12190;
  assign n12192 = ~n12182 & ~n12191_1;
  assign n12193 = ~n12143 & ~n12192;
  assign n12194 = ~n12142 & ~n12193;
  assign n12195 = ~n12132 & ~n12194;
  assign n12196_1 = ~n12131_1 & ~n12195;
  assign n12197 = n12122 & ~n12196_1;
  assign n12198 = ~n11736_1 & n11804;
  assign n12199 = ~n11805 & ~n12198;
  assign n12200 = n11799 & ~n12199;
  assign n12201_1 = ~n11736_1 & ~n11804;
  assign n12202 = ~n11799 & n12201_1;
  assign n12203 = n11800 & n11804;
  assign n12204 = ~n12200 & ~n12202;
  assign n12205 = ~n12203 & n12204;
  assign n12206_1 = ~n12122 & n12196_1;
  assign n12207 = n12205 & ~n12206_1;
  assign n12208 = ~n12197 & ~n12207;
  assign n12209 = n12121_1 & ~n12208;
  assign n12210 = ~n12121_1 & n12208;
  assign n12211_1 = n11735 & ~n11817;
  assign n12212 = ~n11735 & n11817;
  assign n12213 = ~n12211_1 & ~n12212;
  assign n12214 = n11808 & ~n12213;
  assign n12215 = ~n11735 & ~n11817;
  assign n12216_1 = ~n11808 & n12215;
  assign n12217 = n11809 & n11817;
  assign n12218 = ~n12214 & ~n12216_1;
  assign n12219 = ~n12217 & n12218;
  assign n12220 = ~n12210 & ~n12219;
  assign n12221_1 = ~n12209 & ~n12220;
  assign n12222 = n12120 & ~n12221_1;
  assign n12223 = ~n11734 & n11828;
  assign n12224 = ~n11829 & ~n12223;
  assign n12225 = n11820 & ~n12224;
  assign n12226_1 = ~n11734 & ~n11828;
  assign n12227 = ~n11820 & n12226_1;
  assign n12228 = n11821_1 & n11828;
  assign n12229 = ~n12225 & ~n12227;
  assign n12230 = ~n12228 & n12229;
  assign n12231_1 = ~n12120 & n12221_1;
  assign n12232 = n12230 & ~n12231_1;
  assign n12233 = ~n12222 & ~n12232;
  assign n12234 = ~n12119 & ~n12233;
  assign n12235 = ~n12118 & ~n12234;
  assign n12236_1 = ~n12112 & ~n12235;
  assign n12237 = ~n12111_1 & ~n12236_1;
  assign n12238 = ~n12101_1 & ~n12237;
  assign n12239 = ~n12100 & ~n12238;
  assign n12240 = n12091_1 & ~n12239;
  assign n12241_1 = ~n11712 & n11855;
  assign n12242 = ~n11856_1 & ~n12241_1;
  assign n12243 = n11719 & ~n12242;
  assign n12244 = ~n11712 & ~n11855;
  assign n12245 = ~n11719 & n12244;
  assign n12246_1 = n11720 & n11855;
  assign n12247 = ~n12243 & ~n12245;
  assign n12248 = ~n12246_1 & n12247;
  assign n12249 = ~n12091_1 & n12239;
  assign n12250 = n12248 & ~n12249;
  assign n12251_1 = ~n12240 & ~n12250;
  assign n12252 = ~n12090 & ~n12251_1;
  assign n12253 = ~n12089 & ~n12252;
  assign n12254 = n12083 & ~n12253;
  assign n12255 = ~n11710 & n11879;
  assign n12256_1 = ~n11880 & ~n12255;
  assign n12257 = n11871_1 & ~n12256_1;
  assign n12258 = ~n11710 & ~n11879;
  assign n12259 = ~n11871_1 & n12258;
  assign n12260 = n11872 & n11879;
  assign n12261_1 = ~n12257 & ~n12259;
  assign n12262 = ~n12260 & n12261_1;
  assign n12263 = ~n12083 & n12253;
  assign n12264 = n12262 & ~n12263;
  assign n12265 = ~n12254 & ~n12264;
  assign n12266_1 = n12082 & ~n12265;
  assign n12267 = ~n11689 & n11707;
  assign n12268 = n11689 & ~n11707;
  assign n12269 = ~n12267 & ~n12268;
  assign n12270 = n11883 & ~n12269;
  assign n12271_1 = ~n11708 & ~n11709;
  assign n12272 = ~n11883 & ~n12271_1;
  assign n12273 = ~n12270 & ~n12272;
  assign n12274 = ~n12082 & n12265;
  assign n12275 = ~n12273 & ~n12274;
  assign n12276_1 = ~n12266_1 & ~n12275;
  assign n12277 = ~n12081_1 & ~n12276_1;
  assign n12278 = n12081_1 & n12276_1;
  assign MUL_1411_U378 = n12277 | n12278;
  assign n12280 = ~n12266_1 & ~n12274;
  assign n12281_1 = n12273 & n12280;
  assign n12282 = ~n12273 & ~n12280;
  assign MUL_1411_U438 = n12281_1 | n12282;
  assign n12284 = n12083 & ~n12262;
  assign n12285 = ~n12083 & n12262;
  assign n12286_1 = ~n12284 & ~n12285;
  assign n12287 = n12253 & ~n12286_1;
  assign n12288 = ~n12083 & ~n12262;
  assign n12289 = ~n12253 & n12288;
  assign n12290 = n12254 & n12262;
  assign n12291_1 = ~n12287 & ~n12289;
  assign MUL_1411_U10 = n12290 | ~n12291_1;
  assign n12293 = ~n12084 & ~n12088;
  assign n12294 = n12084 & n12088;
  assign n12295 = ~n12293 & ~n12294;
  assign n12296_1 = n12251_1 & ~n12295;
  assign n12297 = ~n12089 & ~n12090;
  assign n12298 = ~n12251_1 & ~n12297;
  assign MUL_1411_U439 = n12296_1 | n12298;
  assign n12300 = n12091_1 & ~n12248;
  assign n12301_1 = ~n12091_1 & n12248;
  assign n12302 = ~n12300 & ~n12301_1;
  assign n12303 = n12239 & ~n12302;
  assign n12304 = ~n12091_1 & ~n12248;
  assign n12305 = ~n12239 & n12304;
  assign n12306_1 = n12240 & n12248;
  assign n12307 = ~n12303 & ~n12305;
  assign MUL_1411_U9 = n12306_1 | ~n12307;
  assign n12309 = ~n12092 & ~n12099;
  assign n12310 = n12092 & n12099;
  assign n12311_1 = ~n12309 & ~n12310;
  assign n12312 = n12237 & ~n12311_1;
  assign n12313 = ~n12100 & ~n12101_1;
  assign n12314 = ~n12237 & ~n12313;
  assign MUL_1411_U440 = n12312 | n12314;
  assign n12316_1 = n12110 & ~n12235;
  assign n12317 = ~n12110 & n12235;
  assign n12318 = ~n12316_1 & ~n12317;
  assign n12319 = ~n12109 & n12318;
  assign n12320 = n12109 & n12317;
  assign n12321_1 = n12111_1 & ~n12235;
  assign n12322 = ~n12319 & ~n12320;
  assign MUL_1411_U8 = n12321_1 | ~n12322;
  assign n12324 = ~n12113 & ~n12117;
  assign n12325 = n12113 & n12117;
  assign n12326_1 = ~n12324 & ~n12325;
  assign n12327 = n12233 & ~n12326_1;
  assign n12328 = ~n12118 & ~n12119;
  assign n12329 = ~n12233 & ~n12328;
  assign MUL_1411_U441 = n12327 | n12329;
  assign n12331_1 = n12120 & ~n12230;
  assign n12332 = ~n12120 & n12230;
  assign n12333 = ~n12331_1 & ~n12332;
  assign n12334 = n12221_1 & ~n12333;
  assign n12335 = ~n12120 & ~n12230;
  assign n12336_1 = ~n12221_1 & n12335;
  assign n12337 = n12222 & n12230;
  assign n12338 = ~n12334 & ~n12336_1;
  assign MUL_1411_U7 = n12337 | ~n12338;
  assign n12340 = ~n12209 & ~n12210;
  assign n12341_1 = n12219 & n12340;
  assign n12342 = ~n12219 & ~n12340;
  assign MUL_1411_U385 = n12341_1 | n12342;
  assign n12344 = n12122 & ~n12205;
  assign n12345 = ~n12122 & n12205;
  assign n12346_1 = ~n12344 & ~n12345;
  assign n12347 = n12196_1 & ~n12346_1;
  assign n12348 = ~n12122 & ~n12205;
  assign n12349 = ~n12196_1 & n12348;
  assign n12350 = n12197 & n12205;
  assign n12351_1 = ~n12347 & ~n12349;
  assign MUL_1411_U14 = n12350 | ~n12351_1;
  assign n12353 = ~n12123 & ~n12130;
  assign n12354 = n12123 & n12130;
  assign n12355 = ~n12353 & ~n12354;
  assign n12356_1 = n12194 & ~n12355;
  assign n12357 = ~n12131_1 & ~n12132;
  assign n12358 = ~n12194 & ~n12357;
  assign MUL_1411_U386 = n12356_1 | n12358;
  assign n12360 = n12141_1 & ~n12192;
  assign n12361_1 = ~n12141_1 & n12192;
  assign n12362 = ~n12360 & ~n12361_1;
  assign n12363 = ~n12140 & n12362;
  assign n12364 = n12140 & n12361_1;
  assign n12365 = n12142 & ~n12192;
  assign n12366_1 = ~n12363 & ~n12364;
  assign MUL_1411_U13 = n12365 | ~n12366_1;
  assign n12368 = ~n12182 & ~n12190;
  assign n12369 = n12189 & n12368;
  assign n12370 = ~n12189 & ~n12368;
  assign MUL_1411_U387 = n12369 | n12370;
  assign n12372 = n12145 & ~n12178;
  assign n12373 = ~n12145 & n12178;
  assign n12374 = ~n12372 & ~n12373;
  assign n12375 = n12169 & ~n12374;
  assign n12376_1 = ~n12145 & ~n12178;
  assign n12377 = ~n12169 & n12376_1;
  assign n12378 = n12170 & n12178;
  assign n12379 = ~n12375 & ~n12377;
  assign MUL_1411_U12 = n12378 | ~n12379;
  assign n12381_1 = ~n12146_1 & ~n12150;
  assign n12382 = n12146_1 & n12150;
  assign n12383 = ~n12381_1 & ~n12382;
  assign n12384 = n12167 & ~n12383;
  assign n12385 = ~n12151_1 & ~n12152;
  assign n12386_1 = ~n12167 & ~n12385;
  assign MUL_1411_U388 = n12384 | n12386_1;
  assign n12388 = n12156_1 & ~n12165;
  assign n12389 = ~n12156_1 & n12165;
  assign n12390 = ~n12388 & ~n12389;
  assign n12391_1 = ~n12155 & n12390;
  assign n12392 = n12155 & n12389;
  assign n12393 = n12157 & ~n12165;
  assign n12394 = ~n12391_1 & ~n12392;
  assign MUL_1411_U11 = n12393 | ~n12394;
  assign n12396_1 = ~n10225 & n11911_1;
  assign n12397 = ~n10238 & ~n12396_1;
  assign n12398 = ~n11706_1 & ~n12397;
  assign n12399 = ~n10216_1 & n11706_1;
  assign n12400 = ~n10226_1 & ~n12399;
  assign n12401_1 = ~n11911_1 & ~n12400;
  assign MUL_1411_U15 = n12398 | n12401_1;
  assign U39 = ~n10223 & ~n11909;
  assign n12404 = ~n10214 & ~n11704;
  assign n12405 = U39 & n12404;
  assign n12406_1 = ~n10060 & n10194;
  assign n12407 = ~P2_P1_ADDRESS_REG_2_ & n10060;
  assign n12408 = ~n12406_1 & ~n12407;
  assign n12409 = ~n11909 & n12408;
  assign n12410 = ~n12404 & n12409;
  assign n12411_1 = n12404 & ~n12409;
  assign n12412 = ~n12410 & ~n12411_1;
  assign n12413 = ~n10106_1 & n11499;
  assign n12414 = ~P1_P1_ADDRESS_REG_2_ & n10106_1;
  assign n12415 = ~n12413 & ~n12414;
  assign n12416_1 = ~n10223 & n12415;
  assign n12417 = ~n12412 & ~n12416_1;
  assign n12418 = n12412 & n12416_1;
  assign n12419 = ~n12417 & ~n12418;
  assign n12420 = n12405 & n12419;
  assign n12421_1 = ~n12405 & ~n12419;
  assign MUL_1421_A1_U5 = n12420 | n12421_1;
  assign n12423 = ~n10214 & ~n11909;
  assign n12424 = ~n10223 & ~n11704;
  assign n12425 = n12423 & ~n12424;
  assign n12426_1 = ~n12423 & n12424;
  assign U154 = n12425 | n12426_1;
  assign n12428 = ~P1_P1_BE_N_REG_3_ & ~P1_P1_BE_N_REG_1_;
  assign n12429 = ~P1_P1_D_C_N_REG & n12428;
  assign n12430 = ~P1_P1_ADS_N_REG & n12429;
  assign n12431_1 = ~P1_P1_BE_N_REG_0_ & n12430;
  assign n12432 = ~P1_P1_ADDRESS_REG_20_ & ~P1_P1_ADDRESS_REG_13_;
  assign n12433 = ~P1_P1_ADDRESS_REG_3_ & n12432;
  assign n12434 = ~P1_P1_ADDRESS_REG_27_ & n12433;
  assign n12435 = ~P1_P1_ADDRESS_REG_2_ & n12434;
  assign n12436_1 = ~P1_P1_ADDRESS_REG_5_ & n12435;
  assign n12437 = ~P1_P1_ADDRESS_REG_15_ & n12436_1;
  assign n12438 = ~P1_P1_ADDRESS_REG_26_ & ~P1_P1_ADDRESS_REG_21_;
  assign n12439 = ~P1_P1_ADDRESS_REG_28_ & n12438;
  assign n12440 = ~P1_P1_ADDRESS_REG_6_ & n12439;
  assign n12441_1 = ~P1_P1_ADDRESS_REG_12_ & n12440;
  assign n12442 = ~P1_P1_ADDRESS_REG_14_ & n12441_1;
  assign n12443 = ~P1_P1_ADDRESS_REG_4_ & n12442;
  assign n12444 = ~P1_P1_ADDRESS_REG_16_ & ~P1_P1_ADDRESS_REG_0_;
  assign n12445 = ~P1_P1_ADDRESS_REG_18_ & n12444;
  assign n12446_1 = ~P1_P1_ADDRESS_REG_8_ & n12445;
  assign n12447 = ~P1_P1_ADDRESS_REG_23_ & n12446_1;
  assign n12448 = ~P1_P1_ADDRESS_REG_1_ & n12447;
  assign n12449 = ~P1_P1_ADDRESS_REG_11_ & n12448;
  assign n12450 = ~P1_P1_ADDRESS_REG_17_ & ~P1_P1_ADDRESS_REG_9_;
  assign n12451_1 = ~P1_P1_ADDRESS_REG_7_ & n12450;
  assign n12452 = ~P1_P1_ADDRESS_REG_22_ & n12451_1;
  assign n12453 = ~P1_P1_ADDRESS_REG_10_ & n12452;
  assign n12454 = ~P1_P1_ADDRESS_REG_19_ & n12453;
  assign n12455 = ~P1_P1_ADDRESS_REG_25_ & n12454;
  assign n12456_1 = ~P1_P1_ADDRESS_REG_24_ & n12455;
  assign n12457 = n12437 & n12443;
  assign n12458 = n12449 & n12457;
  assign n12459 = n12456_1 & n12458;
  assign n12460 = P1_P1_ADDRESS_REG_29_ & ~n12459;
  assign n12461_1 = ~P1_P1_BE_N_REG_2_ & P1_P1_M_IO_N_REG;
  assign n12462 = P1_P1_W_R_N_REG & n12461_1;
  assign n12463 = n12431_1 & n12462;
  assign n456 = ~n12460 | ~n12463;
  assign n12465 = P1_P1_DATAO_REG_0_ & ~n456;
  assign n12466_1 = ~P1_P2_ADDRESS_REG_20_ & ~P1_P2_ADDRESS_REG_13_;
  assign n12467 = ~P1_P2_ADDRESS_REG_3_ & n12466_1;
  assign n12468 = ~P1_P2_ADDRESS_REG_27_ & n12467;
  assign n12469 = ~P1_P2_ADDRESS_REG_2_ & n12468;
  assign n12470 = ~P1_P2_ADDRESS_REG_5_ & n12469;
  assign n12471_1 = ~P1_P2_ADDRESS_REG_15_ & n12470;
  assign n12472 = ~P1_P2_ADDRESS_REG_26_ & ~P1_P2_ADDRESS_REG_21_;
  assign n12473 = ~P1_P2_ADDRESS_REG_28_ & n12472;
  assign n12474 = ~P1_P2_ADDRESS_REG_6_ & n12473;
  assign n12475 = ~P1_P2_ADDRESS_REG_12_ & n12474;
  assign n12476_1 = ~P1_P2_ADDRESS_REG_14_ & n12475;
  assign n12477 = ~P1_P2_ADDRESS_REG_4_ & n12476_1;
  assign n12478 = ~P1_P2_ADDRESS_REG_16_ & ~P1_P2_ADDRESS_REG_0_;
  assign n12479 = ~P1_P2_ADDRESS_REG_18_ & n12478;
  assign n12480 = ~P1_P2_ADDRESS_REG_8_ & n12479;
  assign n12481_1 = ~P1_P2_ADDRESS_REG_23_ & n12480;
  assign n12482 = ~P1_P2_ADDRESS_REG_1_ & n12481_1;
  assign n12483 = ~P1_P2_ADDRESS_REG_11_ & n12482;
  assign n12484 = ~P1_P2_ADDRESS_REG_17_ & ~P1_P2_ADDRESS_REG_9_;
  assign n12485 = ~P1_P2_ADDRESS_REG_7_ & n12484;
  assign n12486_1 = ~P1_P2_ADDRESS_REG_22_ & n12485;
  assign n12487 = ~P1_P2_ADDRESS_REG_10_ & n12486_1;
  assign n12488 = ~P1_P2_ADDRESS_REG_19_ & n12487;
  assign n12489 = ~P1_P2_ADDRESS_REG_25_ & n12488;
  assign n12490 = ~P1_P2_ADDRESS_REG_24_ & n12489;
  assign n12491_1 = n12471_1 & n12477;
  assign n12492 = n12483 & n12491_1;
  assign n12493 = n12490 & n12492;
  assign n12494 = P1_P2_ADDRESS_REG_29_ & ~n12493;
  assign n12495 = ~P1_P2_BE_N_REG_3_ & ~P1_P2_D_C_N_REG;
  assign n12496_1 = ~P1_P2_BE_N_REG_0_ & ~P1_P2_ADS_N_REG;
  assign n12497 = ~P1_P2_BE_N_REG_2_ & n12496_1;
  assign n12498 = ~P1_P2_BE_N_REG_1_ & n12497;
  assign n12499 = P1_P2_W_R_N_REG & P1_P2_M_IO_N_REG;
  assign n12500 = n12495 & n12499;
  assign n12501_1 = n12498 & n12500;
  assign n12502 = n12494 & n12501_1;
  assign n12503 = n456 & ~n12502;
  assign n12504 = P1_BUF1_REG_0_ & n12503;
  assign n12505 = n456 & ~n12503;
  assign n12506_1 = P1_P2_DATAO_REG_0_ & n12505;
  assign n12507 = ~n12465 & ~n12504;
  assign n121 = n12506_1 | ~n12507;
  assign n12509 = P1_P1_DATAO_REG_1_ & ~n456;
  assign n12510 = P1_BUF1_REG_1_ & n12503;
  assign n12511_1 = P1_P2_DATAO_REG_1_ & n12505;
  assign n12512 = ~n12509 & ~n12510;
  assign n126 = n12511_1 | ~n12512;
  assign n12514 = P1_P1_DATAO_REG_2_ & ~n456;
  assign n12515 = P1_BUF1_REG_2_ & n12503;
  assign n12516_1 = P1_P2_DATAO_REG_2_ & n12505;
  assign n12517 = ~n12514 & ~n12515;
  assign n131 = n12516_1 | ~n12517;
  assign n12519 = P1_P1_DATAO_REG_3_ & ~n456;
  assign n12520 = P1_BUF1_REG_3_ & n12503;
  assign n12521_1 = P1_P2_DATAO_REG_3_ & n12505;
  assign n12522 = ~n12519 & ~n12520;
  assign n136 = n12521_1 | ~n12522;
  assign n12524 = P1_P1_DATAO_REG_4_ & ~n456;
  assign n12525 = P1_BUF1_REG_4_ & n12503;
  assign n12526_1 = P1_P2_DATAO_REG_4_ & n12505;
  assign n12527 = ~n12524 & ~n12525;
  assign n141 = n12526_1 | ~n12527;
  assign n12529 = P1_P1_DATAO_REG_5_ & ~n456;
  assign n12530 = P1_BUF1_REG_5_ & n12503;
  assign n12531_1 = P1_P2_DATAO_REG_5_ & n12505;
  assign n12532 = ~n12529 & ~n12530;
  assign n146 = n12531_1 | ~n12532;
  assign n12534 = P1_P1_DATAO_REG_6_ & ~n456;
  assign n12535 = P1_BUF1_REG_6_ & n12503;
  assign n12536_1 = P1_P2_DATAO_REG_6_ & n12505;
  assign n12537 = ~n12534 & ~n12535;
  assign n151 = n12536_1 | ~n12537;
  assign n12539 = P1_P1_DATAO_REG_7_ & ~n456;
  assign n12540 = P1_BUF1_REG_7_ & n12503;
  assign n12541_1 = P1_P2_DATAO_REG_7_ & n12505;
  assign n12542 = ~n12539 & ~n12540;
  assign n156 = n12541_1 | ~n12542;
  assign n12544 = P1_P1_DATAO_REG_8_ & ~n456;
  assign n12545 = P1_BUF1_REG_8_ & n12503;
  assign n12546_1 = P1_P2_DATAO_REG_8_ & n12505;
  assign n12547 = ~n12544 & ~n12545;
  assign n161 = n12546_1 | ~n12547;
  assign n12549 = P1_P1_DATAO_REG_9_ & ~n456;
  assign n12550 = P1_BUF1_REG_9_ & n12503;
  assign n12551_1 = P1_P2_DATAO_REG_9_ & n12505;
  assign n12552 = ~n12549 & ~n12550;
  assign n166 = n12551_1 | ~n12552;
  assign n12554 = P1_P1_DATAO_REG_10_ & ~n456;
  assign n12555 = P1_BUF1_REG_10_ & n12503;
  assign n12556_1 = P1_P2_DATAO_REG_10_ & n12505;
  assign n12557 = ~n12554 & ~n12555;
  assign n171 = n12556_1 | ~n12557;
  assign n12559 = P1_P1_DATAO_REG_11_ & ~n456;
  assign n12560 = P1_BUF1_REG_11_ & n12503;
  assign n12561_1 = P1_P2_DATAO_REG_11_ & n12505;
  assign n12562 = ~n12559 & ~n12560;
  assign n176 = n12561_1 | ~n12562;
  assign n12564 = P1_P1_DATAO_REG_12_ & ~n456;
  assign n12565 = P1_BUF1_REG_12_ & n12503;
  assign n12566_1 = P1_P2_DATAO_REG_12_ & n12505;
  assign n12567 = ~n12564 & ~n12565;
  assign n181 = n12566_1 | ~n12567;
  assign n12569 = P1_P1_DATAO_REG_13_ & ~n456;
  assign n12570 = P1_BUF1_REG_13_ & n12503;
  assign n12571_1 = P1_P2_DATAO_REG_13_ & n12505;
  assign n12572 = ~n12569 & ~n12570;
  assign n186 = n12571_1 | ~n12572;
  assign n12574 = P1_P1_DATAO_REG_14_ & ~n456;
  assign n12575 = P1_BUF1_REG_14_ & n12503;
  assign n12576_1 = P1_P2_DATAO_REG_14_ & n12505;
  assign n12577 = ~n12574 & ~n12575;
  assign n191 = n12576_1 | ~n12577;
  assign n12579 = P1_P1_DATAO_REG_15_ & ~n456;
  assign n12580 = P1_BUF1_REG_15_ & n12503;
  assign n12581_1 = P1_P2_DATAO_REG_15_ & n12505;
  assign n12582 = ~n12579 & ~n12580;
  assign n196 = n12581_1 | ~n12582;
  assign n12584 = P1_P1_DATAO_REG_16_ & ~n456;
  assign n12585 = P1_BUF1_REG_16_ & n12503;
  assign n12586_1 = P1_P2_DATAO_REG_16_ & n12505;
  assign n12587 = ~n12584 & ~n12585;
  assign n201 = n12586_1 | ~n12587;
  assign n12589 = P1_P1_DATAO_REG_17_ & ~n456;
  assign n12590 = P1_BUF1_REG_17_ & n12503;
  assign n12591_1 = P1_P2_DATAO_REG_17_ & n12505;
  assign n12592 = ~n12589 & ~n12590;
  assign n206 = n12591_1 | ~n12592;
  assign n12594 = P1_P1_DATAO_REG_18_ & ~n456;
  assign n12595 = P1_BUF1_REG_18_ & n12503;
  assign n12596_1 = P1_P2_DATAO_REG_18_ & n12505;
  assign n12597 = ~n12594 & ~n12595;
  assign n211 = n12596_1 | ~n12597;
  assign n12599 = P1_P1_DATAO_REG_19_ & ~n456;
  assign n12600 = P1_BUF1_REG_19_ & n12503;
  assign n12601_1 = P1_P2_DATAO_REG_19_ & n12505;
  assign n12602 = ~n12599 & ~n12600;
  assign n216 = n12601_1 | ~n12602;
  assign n12604 = P1_P1_DATAO_REG_20_ & ~n456;
  assign n12605 = P1_BUF1_REG_20_ & n12503;
  assign n12606_1 = P1_P2_DATAO_REG_20_ & n12505;
  assign n12607 = ~n12604 & ~n12605;
  assign n221 = n12606_1 | ~n12607;
  assign n12609 = P1_P1_DATAO_REG_21_ & ~n456;
  assign n12610 = P1_BUF1_REG_21_ & n12503;
  assign n12611_1 = P1_P2_DATAO_REG_21_ & n12505;
  assign n12612 = ~n12609 & ~n12610;
  assign n226 = n12611_1 | ~n12612;
  assign n12614 = P1_P1_DATAO_REG_22_ & ~n456;
  assign n12615 = P1_BUF1_REG_22_ & n12503;
  assign n12616_1 = P1_P2_DATAO_REG_22_ & n12505;
  assign n12617 = ~n12614 & ~n12615;
  assign n231 = n12616_1 | ~n12617;
  assign n12619 = P1_P1_DATAO_REG_23_ & ~n456;
  assign n12620 = P1_BUF1_REG_23_ & n12503;
  assign n12621_1 = P1_P2_DATAO_REG_23_ & n12505;
  assign n12622 = ~n12619 & ~n12620;
  assign n236 = n12621_1 | ~n12622;
  assign n12624 = P1_P1_DATAO_REG_24_ & ~n456;
  assign n12625 = P1_BUF1_REG_24_ & n12503;
  assign n12626_1 = P1_P2_DATAO_REG_24_ & n12505;
  assign n12627 = ~n12624 & ~n12625;
  assign n241 = n12626_1 | ~n12627;
  assign n12629 = P1_P1_DATAO_REG_25_ & ~n456;
  assign n12630 = P1_BUF1_REG_25_ & n12503;
  assign n12631_1 = P1_P2_DATAO_REG_25_ & n12505;
  assign n12632 = ~n12629 & ~n12630;
  assign n246 = n12631_1 | ~n12632;
  assign n12634 = P1_P1_DATAO_REG_26_ & ~n456;
  assign n12635 = P1_BUF1_REG_26_ & n12503;
  assign n12636_1 = P1_P2_DATAO_REG_26_ & n12505;
  assign n12637 = ~n12634 & ~n12635;
  assign n251 = n12636_1 | ~n12637;
  assign n12639 = P1_P1_DATAO_REG_27_ & ~n456;
  assign n12640 = P1_BUF1_REG_27_ & n12503;
  assign n12641_1 = P1_P2_DATAO_REG_27_ & n12505;
  assign n12642 = ~n12639 & ~n12640;
  assign n256 = n12641_1 | ~n12642;
  assign n12644 = P1_P1_DATAO_REG_28_ & ~n456;
  assign n12645 = P1_BUF1_REG_28_ & n12503;
  assign n12646_1 = P1_P2_DATAO_REG_28_ & n12505;
  assign n12647 = ~n12644 & ~n12645;
  assign n261 = n12646_1 | ~n12647;
  assign n12649 = P1_P1_DATAO_REG_29_ & ~n456;
  assign n12650 = P1_BUF1_REG_29_ & n12503;
  assign n12651_1 = P1_P2_DATAO_REG_29_ & n12505;
  assign n12652 = ~n12649 & ~n12650;
  assign n266 = n12651_1 | ~n12652;
  assign n12654 = P1_P1_DATAO_REG_30_ & ~n456;
  assign n12655 = P1_BUF1_REG_30_ & n12503;
  assign n12656_1 = P1_P2_DATAO_REG_30_ & n12505;
  assign n12657 = ~n12654 & ~n12655;
  assign n271 = n12656_1 | ~n12657;
  assign n12659 = P1_P1_DATAO_REG_31_ & ~n456;
  assign n12660 = P1_BUF1_REG_31_ & n12503;
  assign n12661_1 = P1_P2_DATAO_REG_31_ & n12505;
  assign n12662 = ~n12659 & ~n12660;
  assign n276 = n12661_1 | ~n12662;
  assign n446 = P1_P2_ADDRESS_REG_29_ | ~n12501_1;
  assign n12665 = P1_P2_DATAO_REG_0_ & ~n446;
  assign n12666_1 = P1_BUF2_REG_0_ & n446;
  assign n281 = n12665 | n12666_1;
  assign n12668 = P1_P2_DATAO_REG_1_ & ~n446;
  assign n12669 = P1_BUF2_REG_1_ & n446;
  assign n286 = n12668 | n12669;
  assign n12671_1 = P1_P2_DATAO_REG_2_ & ~n446;
  assign n12672 = P1_BUF2_REG_2_ & n446;
  assign n291 = n12671_1 | n12672;
  assign n12674 = P1_P2_DATAO_REG_3_ & ~n446;
  assign n12675 = P1_BUF2_REG_3_ & n446;
  assign n296 = n12674 | n12675;
  assign n12677 = P1_P2_DATAO_REG_4_ & ~n446;
  assign n12678 = P1_BUF2_REG_4_ & n446;
  assign n301 = n12677 | n12678;
  assign n12680 = P1_P2_DATAO_REG_5_ & ~n446;
  assign n12681_1 = P1_BUF2_REG_5_ & n446;
  assign n306 = n12680 | n12681_1;
  assign n12683 = P1_P2_DATAO_REG_6_ & ~n446;
  assign n12684 = P1_BUF2_REG_6_ & n446;
  assign n311 = n12683 | n12684;
  assign n12686_1 = P1_P2_DATAO_REG_7_ & ~n446;
  assign n12687 = P1_BUF2_REG_7_ & n446;
  assign n316 = n12686_1 | n12687;
  assign n12689 = P1_P2_DATAO_REG_8_ & ~n446;
  assign n12690 = P1_BUF2_REG_8_ & n446;
  assign n321 = n12689 | n12690;
  assign n12692 = P1_P2_DATAO_REG_9_ & ~n446;
  assign n12693 = P1_BUF2_REG_9_ & n446;
  assign n326 = n12692 | n12693;
  assign n12695 = P1_P2_DATAO_REG_10_ & ~n446;
  assign n12696_1 = P1_BUF2_REG_10_ & n446;
  assign n331 = n12695 | n12696_1;
  assign n12698 = P1_P2_DATAO_REG_11_ & ~n446;
  assign n12699 = P1_BUF2_REG_11_ & n446;
  assign n336 = n12698 | n12699;
  assign n12701_1 = P1_P2_DATAO_REG_12_ & ~n446;
  assign n12702 = P1_BUF2_REG_12_ & n446;
  assign n341 = n12701_1 | n12702;
  assign n12704 = P1_P2_DATAO_REG_13_ & ~n446;
  assign n12705 = P1_BUF2_REG_13_ & n446;
  assign n346 = n12704 | n12705;
  assign n12707 = P1_P2_DATAO_REG_14_ & ~n446;
  assign n12708 = P1_BUF2_REG_14_ & n446;
  assign n351 = n12707 | n12708;
  assign n12710 = P1_P2_DATAO_REG_15_ & ~n446;
  assign n12711_1 = P1_BUF2_REG_15_ & n446;
  assign n356 = n12710 | n12711_1;
  assign n12713 = P1_P2_DATAO_REG_16_ & ~n446;
  assign n12714 = P1_BUF2_REG_16_ & n446;
  assign n361 = n12713 | n12714;
  assign n12716_1 = P1_P2_DATAO_REG_17_ & ~n446;
  assign n12717 = P1_BUF2_REG_17_ & n446;
  assign n366 = n12716_1 | n12717;
  assign n12719 = P1_P2_DATAO_REG_18_ & ~n446;
  assign n12720 = P1_BUF2_REG_18_ & n446;
  assign n371 = n12719 | n12720;
  assign n12722 = P1_P2_DATAO_REG_19_ & ~n446;
  assign n12723 = P1_BUF2_REG_19_ & n446;
  assign n376 = n12722 | n12723;
  assign n12725 = P1_P2_DATAO_REG_20_ & ~n446;
  assign n12726_1 = P1_BUF2_REG_20_ & n446;
  assign n381 = n12725 | n12726_1;
  assign n12728 = P1_P2_DATAO_REG_21_ & ~n446;
  assign n12729 = P1_BUF2_REG_21_ & n446;
  assign n386 = n12728 | n12729;
  assign n12731_1 = P1_P2_DATAO_REG_22_ & ~n446;
  assign n12732 = P1_BUF2_REG_22_ & n446;
  assign n391 = n12731_1 | n12732;
  assign n12734 = P1_P2_DATAO_REG_23_ & ~n446;
  assign n12735 = P1_BUF2_REG_23_ & n446;
  assign n396 = n12734 | n12735;
  assign n12737 = P1_P2_DATAO_REG_24_ & ~n446;
  assign n12738 = P1_BUF2_REG_24_ & n446;
  assign n401 = n12737 | n12738;
  assign n12740 = P1_P2_DATAO_REG_25_ & ~n446;
  assign n12741_1 = P1_BUF2_REG_25_ & n446;
  assign n406 = n12740 | n12741_1;
  assign n12743 = P1_P2_DATAO_REG_26_ & ~n446;
  assign n12744 = P1_BUF2_REG_26_ & n446;
  assign n411 = n12743 | n12744;
  assign n12746_1 = P1_P2_DATAO_REG_27_ & ~n446;
  assign n12747 = P1_BUF2_REG_27_ & n446;
  assign n416 = n12746_1 | n12747;
  assign n12749 = P1_P2_DATAO_REG_28_ & ~n446;
  assign n12750 = P1_BUF2_REG_28_ & n446;
  assign n421 = n12749 | n12750;
  assign n12752 = P1_P2_DATAO_REG_29_ & ~n446;
  assign n12753 = P1_BUF2_REG_29_ & n446;
  assign n426 = n12752 | n12753;
  assign n12755 = P1_P2_DATAO_REG_30_ & ~n446;
  assign n12756_1 = P1_BUF2_REG_30_ & n446;
  assign n431 = n12755 | n12756_1;
  assign n12758 = P1_P2_DATAO_REG_31_ & ~n446;
  assign n12759 = P1_BUF2_REG_31_ & n446;
  assign n436 = n12758 | n12759;
  assign n441 = ~n456 | ~n12502;
  assign n12762 = ~P1_P3_BE_N_REG_3_ & ~P1_P3_BE_N_REG_2_;
  assign n12763 = ~P1_P3_BE_N_REG_1_ & ~P1_P3_BE_N_REG_0_;
  assign n12764 = ~P1_P3_ADS_N_REG & n12763;
  assign n12765 = ~P1_P3_D_C_N_REG & n12764;
  assign n12766_1 = ~P1_P3_W_R_N_REG & n12765;
  assign n12767 = P1_P3_M_IO_N_REG & n12762;
  assign n12768 = n12766_1 & n12767;
  assign n451 = ~n446 | ~n12768;
  assign n12770 = ~P2_P1_BE_N_REG_3_ & ~P2_P1_BE_N_REG_1_;
  assign n12771_1 = ~P2_P1_D_C_N_REG & n12770;
  assign n12772 = ~P2_P1_ADS_N_REG & n12771_1;
  assign n12773 = ~P2_P1_BE_N_REG_0_ & n12772;
  assign n12774 = ~P2_P1_ADDRESS_REG_20_ & ~P2_P1_ADDRESS_REG_13_;
  assign n12775 = ~P2_P1_ADDRESS_REG_3_ & n12774;
  assign n12776_1 = ~P2_P1_ADDRESS_REG_27_ & n12775;
  assign n12777 = ~P2_P1_ADDRESS_REG_2_ & n12776_1;
  assign n12778 = ~P2_P1_ADDRESS_REG_5_ & n12777;
  assign n12779 = ~P2_P1_ADDRESS_REG_15_ & n12778;
  assign n12780 = ~P2_P1_ADDRESS_REG_26_ & ~P2_P1_ADDRESS_REG_21_;
  assign n12781_1 = ~P2_P1_ADDRESS_REG_28_ & n12780;
  assign n12782 = ~P2_P1_ADDRESS_REG_6_ & n12781_1;
  assign n12783 = ~P2_P1_ADDRESS_REG_12_ & n12782;
  assign n12784 = ~P2_P1_ADDRESS_REG_14_ & n12783;
  assign n12785 = ~P2_P1_ADDRESS_REG_4_ & n12784;
  assign n12786_1 = ~P2_P1_ADDRESS_REG_16_ & ~P2_P1_ADDRESS_REG_0_;
  assign n12787 = ~P2_P1_ADDRESS_REG_18_ & n12786_1;
  assign n12788 = ~P2_P1_ADDRESS_REG_8_ & n12787;
  assign n12789 = ~P2_P1_ADDRESS_REG_23_ & n12788;
  assign n12790 = ~P2_P1_ADDRESS_REG_1_ & n12789;
  assign n12791_1 = ~P2_P1_ADDRESS_REG_11_ & n12790;
  assign n12792 = ~P2_P1_ADDRESS_REG_17_ & ~P2_P1_ADDRESS_REG_9_;
  assign n12793 = ~P2_P1_ADDRESS_REG_7_ & n12792;
  assign n12794 = ~P2_P1_ADDRESS_REG_22_ & n12793;
  assign n12795 = ~P2_P1_ADDRESS_REG_10_ & n12794;
  assign n12796_1 = ~P2_P1_ADDRESS_REG_19_ & n12795;
  assign n12797 = ~P2_P1_ADDRESS_REG_25_ & n12796_1;
  assign n12798 = ~P2_P1_ADDRESS_REG_24_ & n12797;
  assign n12799 = n12779 & n12785;
  assign n12800 = n12791_1 & n12799;
  assign n12801_1 = n12798 & n12800;
  assign n12802 = P2_P1_ADDRESS_REG_29_ & ~n12801_1;
  assign n12803 = ~P2_P1_BE_N_REG_2_ & P2_P1_M_IO_N_REG;
  assign n12804 = P2_P1_W_R_N_REG & n12803;
  assign n12805 = n12773 & n12804;
  assign n796 = ~n12802 | ~n12805;
  assign n12807 = P2_P1_DATAO_REG_0_ & ~n796;
  assign n12808 = ~P2_P2_ADDRESS_REG_20_ & ~P2_P2_ADDRESS_REG_13_;
  assign n12809 = ~P2_P2_ADDRESS_REG_3_ & n12808;
  assign n12810 = ~P2_P2_ADDRESS_REG_27_ & n12809;
  assign n12811_1 = ~P2_P2_ADDRESS_REG_2_ & n12810;
  assign n12812 = ~P2_P2_ADDRESS_REG_5_ & n12811_1;
  assign n12813 = ~P2_P2_ADDRESS_REG_15_ & n12812;
  assign n12814 = ~P2_P2_ADDRESS_REG_26_ & ~P2_P2_ADDRESS_REG_21_;
  assign n12815 = ~P2_P2_ADDRESS_REG_28_ & n12814;
  assign n12816_1 = ~P2_P2_ADDRESS_REG_6_ & n12815;
  assign n12817 = ~P2_P2_ADDRESS_REG_12_ & n12816_1;
  assign n12818 = ~P2_P2_ADDRESS_REG_14_ & n12817;
  assign n12819 = ~P2_P2_ADDRESS_REG_4_ & n12818;
  assign n12820 = ~P2_P2_ADDRESS_REG_16_ & ~P2_P2_ADDRESS_REG_0_;
  assign n12821_1 = ~P2_P2_ADDRESS_REG_18_ & n12820;
  assign n12822 = ~P2_P2_ADDRESS_REG_8_ & n12821_1;
  assign n12823 = ~P2_P2_ADDRESS_REG_23_ & n12822;
  assign n12824 = ~P2_P2_ADDRESS_REG_1_ & n12823;
  assign n12825 = ~P2_P2_ADDRESS_REG_11_ & n12824;
  assign n12826_1 = ~P2_P2_ADDRESS_REG_17_ & ~P2_P2_ADDRESS_REG_9_;
  assign n12827 = ~P2_P2_ADDRESS_REG_7_ & n12826_1;
  assign n12828 = ~P2_P2_ADDRESS_REG_22_ & n12827;
  assign n12829 = ~P2_P2_ADDRESS_REG_10_ & n12828;
  assign n12830 = ~P2_P2_ADDRESS_REG_19_ & n12829;
  assign n12831_1 = ~P2_P2_ADDRESS_REG_25_ & n12830;
  assign n12832 = ~P2_P2_ADDRESS_REG_24_ & n12831_1;
  assign n12833 = n12813 & n12819;
  assign n12834 = n12825 & n12833;
  assign n12835 = n12832 & n12834;
  assign n12836_1 = P2_P2_ADDRESS_REG_29_ & ~n12835;
  assign n12837 = ~P2_P2_BE_N_REG_3_ & ~P2_P2_D_C_N_REG;
  assign n12838 = ~P2_P2_BE_N_REG_0_ & ~P2_P2_ADS_N_REG;
  assign n12839 = ~P2_P2_BE_N_REG_2_ & n12838;
  assign n12840 = ~P2_P2_BE_N_REG_1_ & n12839;
  assign n12841_1 = P2_P2_W_R_N_REG & P2_P2_M_IO_N_REG;
  assign n12842 = n12837 & n12841_1;
  assign n12843 = n12840 & n12842;
  assign n12844 = n12836_1 & n12843;
  assign n12845 = n796 & ~n12844;
  assign n12846_1 = P2_BUF1_REG_0_ & n12845;
  assign n12847 = n796 & ~n12845;
  assign n12848 = P2_P2_DATAO_REG_0_ & n12847;
  assign n12849 = ~n12807 & ~n12846_1;
  assign n461 = n12848 | ~n12849;
  assign n12851_1 = P2_P1_DATAO_REG_1_ & ~n796;
  assign n12852 = P2_BUF1_REG_1_ & n12845;
  assign n12853 = P2_P2_DATAO_REG_1_ & n12847;
  assign n12854 = ~n12851_1 & ~n12852;
  assign n466 = n12853 | ~n12854;
  assign n12856_1 = P2_P1_DATAO_REG_2_ & ~n796;
  assign n12857 = P2_BUF1_REG_2_ & n12845;
  assign n12858 = P2_P2_DATAO_REG_2_ & n12847;
  assign n12859 = ~n12856_1 & ~n12857;
  assign n471 = n12858 | ~n12859;
  assign n12861_1 = P2_P1_DATAO_REG_3_ & ~n796;
  assign n12862 = P2_BUF1_REG_3_ & n12845;
  assign n12863 = P2_P2_DATAO_REG_3_ & n12847;
  assign n12864 = ~n12861_1 & ~n12862;
  assign n476 = n12863 | ~n12864;
  assign n12866_1 = P2_P1_DATAO_REG_4_ & ~n796;
  assign n12867 = P2_BUF1_REG_4_ & n12845;
  assign n12868 = P2_P2_DATAO_REG_4_ & n12847;
  assign n12869 = ~n12866_1 & ~n12867;
  assign n481 = n12868 | ~n12869;
  assign n12871_1 = P2_P1_DATAO_REG_5_ & ~n796;
  assign n12872 = P2_BUF1_REG_5_ & n12845;
  assign n12873 = P2_P2_DATAO_REG_5_ & n12847;
  assign n12874 = ~n12871_1 & ~n12872;
  assign n486 = n12873 | ~n12874;
  assign n12876_1 = P2_P1_DATAO_REG_6_ & ~n796;
  assign n12877 = P2_BUF1_REG_6_ & n12845;
  assign n12878 = P2_P2_DATAO_REG_6_ & n12847;
  assign n12879 = ~n12876_1 & ~n12877;
  assign n491 = n12878 | ~n12879;
  assign n12881_1 = P2_P1_DATAO_REG_7_ & ~n796;
  assign n12882 = P2_BUF1_REG_7_ & n12845;
  assign n12883 = P2_P2_DATAO_REG_7_ & n12847;
  assign n12884 = ~n12881_1 & ~n12882;
  assign n496 = n12883 | ~n12884;
  assign n12886_1 = P2_P1_DATAO_REG_8_ & ~n796;
  assign n12887 = P2_BUF1_REG_8_ & n12845;
  assign n12888 = P2_P2_DATAO_REG_8_ & n12847;
  assign n12889 = ~n12886_1 & ~n12887;
  assign n501 = n12888 | ~n12889;
  assign n12891_1 = P2_P1_DATAO_REG_9_ & ~n796;
  assign n12892 = P2_BUF1_REG_9_ & n12845;
  assign n12893 = P2_P2_DATAO_REG_9_ & n12847;
  assign n12894 = ~n12891_1 & ~n12892;
  assign n506 = n12893 | ~n12894;
  assign n12896_1 = P2_P1_DATAO_REG_10_ & ~n796;
  assign n12897 = P2_BUF1_REG_10_ & n12845;
  assign n12898 = P2_P2_DATAO_REG_10_ & n12847;
  assign n12899 = ~n12896_1 & ~n12897;
  assign n511 = n12898 | ~n12899;
  assign n12901_1 = P2_P1_DATAO_REG_11_ & ~n796;
  assign n12902 = P2_BUF1_REG_11_ & n12845;
  assign n12903 = P2_P2_DATAO_REG_11_ & n12847;
  assign n12904 = ~n12901_1 & ~n12902;
  assign n516 = n12903 | ~n12904;
  assign n12906_1 = P2_P1_DATAO_REG_12_ & ~n796;
  assign n12907 = P2_BUF1_REG_12_ & n12845;
  assign n12908 = P2_P2_DATAO_REG_12_ & n12847;
  assign n12909 = ~n12906_1 & ~n12907;
  assign n521 = n12908 | ~n12909;
  assign n12911_1 = P2_P1_DATAO_REG_13_ & ~n796;
  assign n12912 = P2_BUF1_REG_13_ & n12845;
  assign n12913 = P2_P2_DATAO_REG_13_ & n12847;
  assign n12914 = ~n12911_1 & ~n12912;
  assign n526 = n12913 | ~n12914;
  assign n12916_1 = P2_P1_DATAO_REG_14_ & ~n796;
  assign n12917 = P2_BUF1_REG_14_ & n12845;
  assign n12918 = P2_P2_DATAO_REG_14_ & n12847;
  assign n12919 = ~n12916_1 & ~n12917;
  assign n531 = n12918 | ~n12919;
  assign n12921_1 = P2_P1_DATAO_REG_15_ & ~n796;
  assign n12922 = P2_BUF1_REG_15_ & n12845;
  assign n12923 = P2_P2_DATAO_REG_15_ & n12847;
  assign n12924 = ~n12921_1 & ~n12922;
  assign n536 = n12923 | ~n12924;
  assign n12926_1 = P2_P1_DATAO_REG_16_ & ~n796;
  assign n12927 = P2_BUF1_REG_16_ & n12845;
  assign n12928 = P2_P2_DATAO_REG_16_ & n12847;
  assign n12929 = ~n12926_1 & ~n12927;
  assign n541 = n12928 | ~n12929;
  assign n12931_1 = P2_P1_DATAO_REG_17_ & ~n796;
  assign n12932 = P2_BUF1_REG_17_ & n12845;
  assign n12933 = P2_P2_DATAO_REG_17_ & n12847;
  assign n12934 = ~n12931_1 & ~n12932;
  assign n546 = n12933 | ~n12934;
  assign n12936_1 = P2_P1_DATAO_REG_18_ & ~n796;
  assign n12937 = P2_BUF1_REG_18_ & n12845;
  assign n12938 = P2_P2_DATAO_REG_18_ & n12847;
  assign n12939 = ~n12936_1 & ~n12937;
  assign n551 = n12938 | ~n12939;
  assign n12941_1 = P2_P1_DATAO_REG_19_ & ~n796;
  assign n12942 = P2_BUF1_REG_19_ & n12845;
  assign n12943 = P2_P2_DATAO_REG_19_ & n12847;
  assign n12944 = ~n12941_1 & ~n12942;
  assign n556 = n12943 | ~n12944;
  assign n12946_1 = P2_P1_DATAO_REG_20_ & ~n796;
  assign n12947 = P2_BUF1_REG_20_ & n12845;
  assign n12948 = P2_P2_DATAO_REG_20_ & n12847;
  assign n12949 = ~n12946_1 & ~n12947;
  assign n561 = n12948 | ~n12949;
  assign n12951_1 = P2_P1_DATAO_REG_21_ & ~n796;
  assign n12952 = P2_BUF1_REG_21_ & n12845;
  assign n12953 = P2_P2_DATAO_REG_21_ & n12847;
  assign n12954 = ~n12951_1 & ~n12952;
  assign n566 = n12953 | ~n12954;
  assign n12956_1 = P2_P1_DATAO_REG_22_ & ~n796;
  assign n12957 = P2_BUF1_REG_22_ & n12845;
  assign n12958 = P2_P2_DATAO_REG_22_ & n12847;
  assign n12959 = ~n12956_1 & ~n12957;
  assign n571 = n12958 | ~n12959;
  assign n12961_1 = P2_P1_DATAO_REG_23_ & ~n796;
  assign n12962 = P2_BUF1_REG_23_ & n12845;
  assign n12963 = P2_P2_DATAO_REG_23_ & n12847;
  assign n12964 = ~n12961_1 & ~n12962;
  assign n576 = n12963 | ~n12964;
  assign n12966_1 = P2_P1_DATAO_REG_24_ & ~n796;
  assign n12967 = P2_BUF1_REG_24_ & n12845;
  assign n12968 = P2_P2_DATAO_REG_24_ & n12847;
  assign n12969 = ~n12966_1 & ~n12967;
  assign n581 = n12968 | ~n12969;
  assign n12971_1 = P2_P1_DATAO_REG_25_ & ~n796;
  assign n12972 = P2_BUF1_REG_25_ & n12845;
  assign n12973 = P2_P2_DATAO_REG_25_ & n12847;
  assign n12974 = ~n12971_1 & ~n12972;
  assign n586 = n12973 | ~n12974;
  assign n12976_1 = P2_P1_DATAO_REG_26_ & ~n796;
  assign n12977 = P2_BUF1_REG_26_ & n12845;
  assign n12978 = P2_P2_DATAO_REG_26_ & n12847;
  assign n12979 = ~n12976_1 & ~n12977;
  assign n591 = n12978 | ~n12979;
  assign n12981_1 = P2_P1_DATAO_REG_27_ & ~n796;
  assign n12982 = P2_BUF1_REG_27_ & n12845;
  assign n12983 = P2_P2_DATAO_REG_27_ & n12847;
  assign n12984 = ~n12981_1 & ~n12982;
  assign n596 = n12983 | ~n12984;
  assign n12986_1 = P2_P1_DATAO_REG_28_ & ~n796;
  assign n12987 = P2_BUF1_REG_28_ & n12845;
  assign n12988 = P2_P2_DATAO_REG_28_ & n12847;
  assign n12989 = ~n12986_1 & ~n12987;
  assign n601 = n12988 | ~n12989;
  assign n12991_1 = P2_P1_DATAO_REG_29_ & ~n796;
  assign n12992 = P2_BUF1_REG_29_ & n12845;
  assign n12993 = P2_P2_DATAO_REG_29_ & n12847;
  assign n12994 = ~n12991_1 & ~n12992;
  assign n606 = n12993 | ~n12994;
  assign n12996_1 = P2_P1_DATAO_REG_30_ & ~n796;
  assign n12997 = P2_BUF1_REG_30_ & n12845;
  assign n12998 = P2_P2_DATAO_REG_30_ & n12847;
  assign n12999 = ~n12996_1 & ~n12997;
  assign n611 = n12998 | ~n12999;
  assign n13001_1 = P2_P1_DATAO_REG_31_ & ~n796;
  assign n13002 = P2_BUF1_REG_31_ & n12845;
  assign n13003 = P2_P2_DATAO_REG_31_ & n12847;
  assign n13004 = ~n13001_1 & ~n13002;
  assign n616 = n13003 | ~n13004;
  assign n786 = P2_P2_ADDRESS_REG_29_ | ~n12843;
  assign n13007 = P2_P2_DATAO_REG_0_ & ~n786;
  assign n13008 = P2_BUF2_REG_0_ & n786;
  assign n621 = n13007 | n13008;
  assign n13010 = P2_P2_DATAO_REG_1_ & ~n786;
  assign n13011_1 = P2_BUF2_REG_1_ & n786;
  assign n626 = n13010 | n13011_1;
  assign n13013 = P2_P2_DATAO_REG_2_ & ~n786;
  assign n13014 = P2_BUF2_REG_2_ & n786;
  assign n631 = n13013 | n13014;
  assign n13016_1 = P2_P2_DATAO_REG_3_ & ~n786;
  assign n13017 = P2_BUF2_REG_3_ & n786;
  assign n636 = n13016_1 | n13017;
  assign n13019 = P2_P2_DATAO_REG_4_ & ~n786;
  assign n13020 = P2_BUF2_REG_4_ & n786;
  assign n641 = n13019 | n13020;
  assign n13022 = P2_P2_DATAO_REG_5_ & ~n786;
  assign n13023 = P2_BUF2_REG_5_ & n786;
  assign n646 = n13022 | n13023;
  assign n13025 = P2_P2_DATAO_REG_6_ & ~n786;
  assign n13026_1 = P2_BUF2_REG_6_ & n786;
  assign n651 = n13025 | n13026_1;
  assign n13028 = P2_P2_DATAO_REG_7_ & ~n786;
  assign n13029 = P2_BUF2_REG_7_ & n786;
  assign n656 = n13028 | n13029;
  assign n13031_1 = P2_P2_DATAO_REG_8_ & ~n786;
  assign n13032 = P2_BUF2_REG_8_ & n786;
  assign n661 = n13031_1 | n13032;
  assign n13034 = P2_P2_DATAO_REG_9_ & ~n786;
  assign n13035 = P2_BUF2_REG_9_ & n786;
  assign n666 = n13034 | n13035;
  assign n13037 = P2_P2_DATAO_REG_10_ & ~n786;
  assign n13038 = P2_BUF2_REG_10_ & n786;
  assign n671 = n13037 | n13038;
  assign n13040 = P2_P2_DATAO_REG_11_ & ~n786;
  assign n13041_1 = P2_BUF2_REG_11_ & n786;
  assign n676 = n13040 | n13041_1;
  assign n13043 = P2_P2_DATAO_REG_12_ & ~n786;
  assign n13044 = P2_BUF2_REG_12_ & n786;
  assign n681 = n13043 | n13044;
  assign n13046_1 = P2_P2_DATAO_REG_13_ & ~n786;
  assign n13047 = P2_BUF2_REG_13_ & n786;
  assign n686 = n13046_1 | n13047;
  assign n13049 = P2_P2_DATAO_REG_14_ & ~n786;
  assign n13050 = P2_BUF2_REG_14_ & n786;
  assign n691 = n13049 | n13050;
  assign n13052 = P2_P2_DATAO_REG_15_ & ~n786;
  assign n13053 = P2_BUF2_REG_15_ & n786;
  assign n696 = n13052 | n13053;
  assign n13055 = P2_P2_DATAO_REG_16_ & ~n786;
  assign n13056_1 = P2_BUF2_REG_16_ & n786;
  assign n701 = n13055 | n13056_1;
  assign n13058 = P2_P2_DATAO_REG_17_ & ~n786;
  assign n13059 = P2_BUF2_REG_17_ & n786;
  assign n706 = n13058 | n13059;
  assign n13061_1 = P2_P2_DATAO_REG_18_ & ~n786;
  assign n13062 = P2_BUF2_REG_18_ & n786;
  assign n711 = n13061_1 | n13062;
  assign n13064 = P2_P2_DATAO_REG_19_ & ~n786;
  assign n13065 = P2_BUF2_REG_19_ & n786;
  assign n716 = n13064 | n13065;
  assign n13067 = P2_P2_DATAO_REG_20_ & ~n786;
  assign n13068 = P2_BUF2_REG_20_ & n786;
  assign n721 = n13067 | n13068;
  assign n13070 = P2_P2_DATAO_REG_21_ & ~n786;
  assign n13071_1 = P2_BUF2_REG_21_ & n786;
  assign n726 = n13070 | n13071_1;
  assign n13073 = P2_P2_DATAO_REG_22_ & ~n786;
  assign n13074 = P2_BUF2_REG_22_ & n786;
  assign n731 = n13073 | n13074;
  assign n13076_1 = P2_P2_DATAO_REG_23_ & ~n786;
  assign n13077 = P2_BUF2_REG_23_ & n786;
  assign n736 = n13076_1 | n13077;
  assign n13079 = P2_P2_DATAO_REG_24_ & ~n786;
  assign n13080 = P2_BUF2_REG_24_ & n786;
  assign n741 = n13079 | n13080;
  assign n13082 = P2_P2_DATAO_REG_25_ & ~n786;
  assign n13083 = P2_BUF2_REG_25_ & n786;
  assign n746 = n13082 | n13083;
  assign n13085 = P2_P2_DATAO_REG_26_ & ~n786;
  assign n13086_1 = P2_BUF2_REG_26_ & n786;
  assign n751 = n13085 | n13086_1;
  assign n13088 = P2_P2_DATAO_REG_27_ & ~n786;
  assign n13089 = P2_BUF2_REG_27_ & n786;
  assign n756 = n13088 | n13089;
  assign n13091_1 = P2_P2_DATAO_REG_28_ & ~n786;
  assign n13092 = P2_BUF2_REG_28_ & n786;
  assign n761 = n13091_1 | n13092;
  assign n13094 = P2_P2_DATAO_REG_29_ & ~n786;
  assign n13095 = P2_BUF2_REG_29_ & n786;
  assign n766 = n13094 | n13095;
  assign n13097 = P2_P2_DATAO_REG_30_ & ~n786;
  assign n13098 = P2_BUF2_REG_30_ & n786;
  assign n771 = n13097 | n13098;
  assign n13100 = P2_P2_DATAO_REG_31_ & ~n786;
  assign n13101_1 = P2_BUF2_REG_31_ & n786;
  assign n776 = n13100 | n13101_1;
  assign n781 = ~n796 | ~n12844;
  assign n13104 = ~P2_P3_BE_N_REG_3_ & ~P2_P3_BE_N_REG_2_;
  assign n13105 = ~P2_P3_BE_N_REG_1_ & ~P2_P3_BE_N_REG_0_;
  assign n13106_1 = ~P2_P3_ADS_N_REG & n13105;
  assign n13107 = ~P2_P3_D_C_N_REG & n13106_1;
  assign n13108 = ~P2_P3_W_R_N_REG & n13107;
  assign n13109 = P2_P3_M_IO_N_REG & n13104;
  assign n13110 = n13108 & n13109;
  assign n791 = ~n786 | ~n13110;
  assign n13112 = ~P3_IR_REG_31_ & P3_STATE_REG;
  assign n13113 = P3_IR_REG_0_ & n13112;
  assign n13114 = ~P3_STATE_REG & P1_P3_DATAO_REG_0_;
  assign n13115 = ~n13113 & ~n13114;
  assign n13116_1 = P3_STATE_REG & ~n13112;
  assign n13117 = P3_IR_REG_0_ & n13116_1;
  assign n801 = ~n13115 | n13117;
  assign n13119 = P3_IR_REG_1_ & n13112;
  assign n13120 = ~P3_STATE_REG & P1_P3_DATAO_REG_1_;
  assign n13121_1 = ~n13119 & ~n13120;
  assign n13122 = P3_IR_REG_0_ & ~P3_IR_REG_1_;
  assign n13123 = ~P3_IR_REG_0_ & P3_IR_REG_1_;
  assign n13124 = ~n13122 & ~n13123;
  assign n13125 = n13116_1 & ~n13124;
  assign n806 = ~n13121_1 | n13125;
  assign n13127 = P3_IR_REG_2_ & n13112;
  assign n13128 = ~P3_STATE_REG & P1_P3_DATAO_REG_2_;
  assign n13129 = ~n13127 & ~n13128;
  assign n13130 = ~P3_IR_REG_0_ & ~P3_IR_REG_1_;
  assign n13131_1 = P3_IR_REG_2_ & ~n13130;
  assign n13132 = ~P3_IR_REG_2_ & n13130;
  assign n13133 = ~n13131_1 & ~n13132;
  assign n13134 = n13116_1 & n13133;
  assign n811 = ~n13129 | n13134;
  assign n13136_1 = P3_IR_REG_3_ & n13112;
  assign n13137 = ~P3_STATE_REG & P1_P3_DATAO_REG_3_;
  assign n13138 = ~n13136_1 & ~n13137;
  assign n13139 = P3_IR_REG_3_ & ~n13132;
  assign n13140 = ~P3_IR_REG_3_ & n13132;
  assign n13141_1 = ~n13139 & ~n13140;
  assign n13142 = n13116_1 & n13141_1;
  assign n816 = ~n13138 | n13142;
  assign n13144 = P3_IR_REG_4_ & n13112;
  assign n13145 = ~P3_STATE_REG & P1_P3_DATAO_REG_4_;
  assign n13146_1 = ~n13144 & ~n13145;
  assign n13147 = P3_IR_REG_4_ & ~n13140;
  assign n13148 = ~P3_IR_REG_3_ & ~P3_IR_REG_4_;
  assign n13149 = n13132 & n13148;
  assign n13150 = ~n13147 & ~n13149;
  assign n13151_1 = n13116_1 & n13150;
  assign n821 = ~n13146_1 | n13151_1;
  assign n13153 = P3_IR_REG_5_ & n13112;
  assign n13154 = ~P3_STATE_REG & P1_P3_DATAO_REG_5_;
  assign n13155 = ~n13153 & ~n13154;
  assign n13156_1 = ~P3_IR_REG_5_ & n13149;
  assign n13157 = P3_IR_REG_5_ & ~n13149;
  assign n13158 = ~n13156_1 & ~n13157;
  assign n13159 = n13116_1 & n13158;
  assign n826 = ~n13155 | n13159;
  assign n13161_1 = P3_IR_REG_6_ & n13112;
  assign n13162 = ~P3_STATE_REG & P1_P3_DATAO_REG_6_;
  assign n13163 = ~n13161_1 & ~n13162;
  assign n13164 = P3_IR_REG_6_ & ~n13156_1;
  assign n13165 = ~P3_IR_REG_5_ & ~P3_IR_REG_6_;
  assign n13166_1 = n13149 & n13165;
  assign n13167 = ~n13164 & ~n13166_1;
  assign n13168 = n13116_1 & n13167;
  assign n831 = ~n13163 | n13168;
  assign n13170 = P3_IR_REG_7_ & n13112;
  assign n13171_1 = ~P3_STATE_REG & P1_P3_DATAO_REG_7_;
  assign n13172 = ~n13170 & ~n13171_1;
  assign n13173 = P3_IR_REG_7_ & ~n13166_1;
  assign n13174 = ~P3_IR_REG_7_ & n13166_1;
  assign n13175 = ~n13173 & ~n13174;
  assign n13176_1 = n13116_1 & n13175;
  assign n836 = ~n13172 | n13176_1;
  assign n13178 = P3_IR_REG_8_ & n13112;
  assign n13179 = ~P3_STATE_REG & P1_P3_DATAO_REG_8_;
  assign n13180 = ~n13178 & ~n13179;
  assign n13181_1 = P3_IR_REG_8_ & ~n13174;
  assign n13182 = ~P3_IR_REG_7_ & ~P3_IR_REG_8_;
  assign n13183 = ~P3_IR_REG_5_ & n13148;
  assign n13184 = ~P3_IR_REG_6_ & n13183;
  assign n13185 = n13132 & n13182;
  assign n13186_1 = n13184 & n13185;
  assign n13187 = ~n13181_1 & ~n13186_1;
  assign n13188 = n13116_1 & n13187;
  assign n841 = ~n13180 | n13188;
  assign n13190 = P3_IR_REG_9_ & n13112;
  assign n13191_1 = ~P3_STATE_REG & P1_P3_DATAO_REG_9_;
  assign n13192 = ~n13190 & ~n13191_1;
  assign n13193 = ~P3_IR_REG_9_ & n13186_1;
  assign n13194 = P3_IR_REG_9_ & ~n13186_1;
  assign n13195 = ~n13193 & ~n13194;
  assign n13196_1 = n13116_1 & n13195;
  assign n846 = ~n13192 | n13196_1;
  assign n13198 = P3_IR_REG_10_ & n13112;
  assign n13199 = ~P3_STATE_REG & P1_P3_DATAO_REG_10_;
  assign n13200 = ~n13198 & ~n13199;
  assign n13201_1 = P3_IR_REG_10_ & ~n13193;
  assign n13202 = ~P3_IR_REG_9_ & ~P3_IR_REG_10_;
  assign n13203 = n13186_1 & n13202;
  assign n13204 = ~n13201_1 & ~n13203;
  assign n13205 = n13116_1 & n13204;
  assign n851 = ~n13200 | n13205;
  assign n13207 = P3_IR_REG_11_ & n13112;
  assign n13208 = ~P3_STATE_REG & P1_P3_DATAO_REG_11_;
  assign n13209 = ~n13207 & ~n13208;
  assign n13210 = P3_IR_REG_11_ & ~n13203;
  assign n13211_1 = ~P3_IR_REG_11_ & n13203;
  assign n13212 = ~n13210 & ~n13211_1;
  assign n13213 = n13116_1 & n13212;
  assign n856 = ~n13209 | n13213;
  assign n13215 = P3_IR_REG_12_ & n13112;
  assign n13216_1 = ~P3_STATE_REG & P1_P3_DATAO_REG_12_;
  assign n13217 = ~n13215 & ~n13216_1;
  assign n13218 = P3_IR_REG_12_ & ~n13211_1;
  assign n13219 = ~P3_IR_REG_10_ & ~P3_IR_REG_11_;
  assign n13220 = ~P3_IR_REG_12_ & n13219;
  assign n13221_1 = ~P3_IR_REG_9_ & n13220;
  assign n13222 = n13186_1 & n13221_1;
  assign n13223 = ~n13218 & ~n13222;
  assign n13224 = n13116_1 & n13223;
  assign n861 = ~n13217 | n13224;
  assign n13226_1 = P3_IR_REG_13_ & n13112;
  assign n13227 = ~P3_STATE_REG & P1_P3_DATAO_REG_13_;
  assign n13228 = ~n13226_1 & ~n13227;
  assign n13229 = ~P3_IR_REG_13_ & n13222;
  assign n13230 = P3_IR_REG_13_ & ~n13222;
  assign n13231_1 = ~n13229 & ~n13230;
  assign n13232 = n13116_1 & n13231_1;
  assign n866 = ~n13228 | n13232;
  assign n13234 = P3_IR_REG_14_ & n13112;
  assign n13235 = ~P3_STATE_REG & P1_P3_DATAO_REG_14_;
  assign n13236_1 = ~n13234 & ~n13235;
  assign n13237 = P3_IR_REG_14_ & ~n13229;
  assign n13238 = ~P3_IR_REG_13_ & ~P3_IR_REG_14_;
  assign n13239 = n13222 & n13238;
  assign n13240 = ~n13237 & ~n13239;
  assign n13241_1 = n13116_1 & n13240;
  assign n871 = ~n13236_1 | n13241_1;
  assign n13243 = P3_IR_REG_15_ & n13112;
  assign n13244 = ~P3_STATE_REG & P1_P3_DATAO_REG_15_;
  assign n13245 = ~n13243 & ~n13244;
  assign n13246_1 = P3_IR_REG_15_ & ~n13239;
  assign n13247 = ~P3_IR_REG_15_ & n13239;
  assign n13248 = ~n13246_1 & ~n13247;
  assign n13249 = n13116_1 & n13248;
  assign n876 = ~n13245 | n13249;
  assign n13251_1 = P3_IR_REG_16_ & n13112;
  assign n13252 = ~P3_STATE_REG & P1_P3_DATAO_REG_16_;
  assign n13253 = ~n13251_1 & ~n13252;
  assign n13254 = P3_IR_REG_16_ & ~n13247;
  assign n13255 = ~P3_IR_REG_6_ & ~P3_IR_REG_7_;
  assign n13256_1 = ~P3_IR_REG_8_ & n13255;
  assign n13257 = ~P3_IR_REG_9_ & n13256_1;
  assign n13258 = ~P3_IR_REG_2_ & ~P3_IR_REG_3_;
  assign n13259 = ~P3_IR_REG_4_ & n13258;
  assign n13260 = ~P3_IR_REG_5_ & n13259;
  assign n13261_1 = ~P3_IR_REG_15_ & ~P3_IR_REG_16_;
  assign n13262 = ~P3_IR_REG_1_ & n13261_1;
  assign n13263 = ~P3_IR_REG_0_ & n13262;
  assign n13264 = ~P3_IR_REG_12_ & n13238;
  assign n13265 = ~P3_IR_REG_10_ & n13264;
  assign n13266_1 = ~P3_IR_REG_11_ & n13265;
  assign n13267 = n13257 & n13260;
  assign n13268 = n13263 & n13267;
  assign n13269 = n13266_1 & n13268;
  assign n13270 = ~n13254 & ~n13269;
  assign n13271_1 = n13116_1 & n13270;
  assign n881 = ~n13253 | n13271_1;
  assign n13273 = P3_IR_REG_17_ & n13112;
  assign n13274 = ~P3_STATE_REG & P1_P3_DATAO_REG_17_;
  assign n13275 = ~n13273 & ~n13274;
  assign n13276_1 = ~P3_IR_REG_17_ & n13269;
  assign n13277 = P3_IR_REG_17_ & ~n13269;
  assign n13278 = ~n13276_1 & ~n13277;
  assign n13279 = n13116_1 & n13278;
  assign n886 = ~n13275 | n13279;
  assign n13281_1 = P3_IR_REG_18_ & n13112;
  assign n13282 = ~P3_STATE_REG & P1_P3_DATAO_REG_18_;
  assign n13283 = ~n13281_1 & ~n13282;
  assign n13284 = P3_IR_REG_18_ & ~n13276_1;
  assign n13285 = ~P3_IR_REG_4_ & ~P3_IR_REG_5_;
  assign n13286_1 = ~P3_IR_REG_3_ & n13285;
  assign n13287 = ~P3_IR_REG_0_ & n13286_1;
  assign n13288 = ~P3_IR_REG_2_ & n13287;
  assign n13289 = ~P3_IR_REG_1_ & ~P3_IR_REG_18_;
  assign n13290 = ~P3_IR_REG_17_ & n13289;
  assign n13291_1 = ~P3_IR_REG_15_ & n13290;
  assign n13292 = ~P3_IR_REG_16_ & n13291_1;
  assign n13293 = n13257 & n13288;
  assign n13294 = n13292 & n13293;
  assign n13295 = n13266_1 & n13294;
  assign n13296_1 = ~n13284 & ~n13295;
  assign n13297 = n13116_1 & n13296_1;
  assign n891 = ~n13283 | n13297;
  assign n13299 = P3_IR_REG_19_ & n13112;
  assign n13300 = ~P3_STATE_REG & P1_P3_DATAO_REG_19_;
  assign n13301_1 = ~n13299 & ~n13300;
  assign n13302 = P3_IR_REG_19_ & ~n13295;
  assign n13303 = ~P3_IR_REG_8_ & ~P3_IR_REG_9_;
  assign n13304 = ~P3_IR_REG_7_ & n13303;
  assign n13305 = ~P3_IR_REG_5_ & n13304;
  assign n13306_1 = ~P3_IR_REG_6_ & n13305;
  assign n13307 = ~P3_IR_REG_2_ & n13148;
  assign n13308 = ~P3_IR_REG_1_ & n13307;
  assign n13309 = ~P3_IR_REG_0_ & n13308;
  assign n13310 = ~P3_IR_REG_18_ & ~P3_IR_REG_19_;
  assign n13311_1 = ~P3_IR_REG_17_ & n13310;
  assign n13312 = ~P3_IR_REG_15_ & n13311_1;
  assign n13313 = ~P3_IR_REG_16_ & n13312;
  assign n13314 = n13306_1 & n13309;
  assign n13315 = n13313 & n13314;
  assign n13316_1 = n13266_1 & n13315;
  assign n13317 = ~n13302 & ~n13316_1;
  assign n13318 = n13116_1 & n13317;
  assign n896 = ~n13301_1 | n13318;
  assign n13320 = P3_IR_REG_20_ & n13112;
  assign n13321_1 = LOGIC0 & ~P3_STATE_REG;
  assign n13322 = ~n13320 & ~n13321_1;
  assign n13323 = P3_IR_REG_20_ & ~n13316_1;
  assign n13324 = ~P3_IR_REG_13_ & ~P3_IR_REG_15_;
  assign n13325 = ~P3_IR_REG_14_ & n13324;
  assign n13326_1 = ~P3_IR_REG_10_ & ~P3_IR_REG_12_;
  assign n13327 = ~P3_IR_REG_11_ & n13326_1;
  assign n13328 = ~P3_IR_REG_1_ & ~P3_IR_REG_19_;
  assign n13329 = ~P3_IR_REG_18_ & n13328;
  assign n13330 = ~P3_IR_REG_16_ & n13329;
  assign n13331_1 = ~P3_IR_REG_17_ & n13330;
  assign n13332 = ~P3_IR_REG_0_ & n13307;
  assign n13333 = ~P3_IR_REG_20_ & n13332;
  assign n13334 = n13325 & n13327;
  assign n13335 = n13331_1 & n13334;
  assign n13336_1 = n13306_1 & n13335;
  assign n13337 = n13333 & n13336_1;
  assign n13338 = ~n13323 & ~n13337;
  assign n13339 = n13116_1 & n13338;
  assign n901 = ~n13322 | n13339;
  assign n13341_1 = P3_IR_REG_21_ & n13112;
  assign n13342 = ~n13321_1 & ~n13341_1;
  assign n13343 = ~P3_IR_REG_21_ & n13337;
  assign n13344 = P3_IR_REG_21_ & ~n13337;
  assign n13345 = ~n13343 & ~n13344;
  assign n13346_1 = n13116_1 & n13345;
  assign n906 = ~n13342 | n13346_1;
  assign n13348 = P3_IR_REG_22_ & n13112;
  assign n13349 = ~n13321_1 & ~n13348;
  assign n13350 = ~P3_IR_REG_2_ & ~P3_IR_REG_4_;
  assign n13351_1 = ~P3_IR_REG_3_ & n13350;
  assign n13352 = ~P3_IR_REG_0_ & ~P3_IR_REG_21_;
  assign n13353 = ~P3_IR_REG_20_ & n13352;
  assign n13354 = n13351_1 & n13353;
  assign n13355 = n13306_1 & n13354;
  assign n13356_1 = n13331_1 & n13355;
  assign n13357 = n13334 & n13356_1;
  assign n13358 = P3_IR_REG_22_ & ~n13357;
  assign n13359 = ~P3_IR_REG_19_ & ~P3_IR_REG_20_;
  assign n13360 = ~P3_IR_REG_17_ & ~P3_IR_REG_18_;
  assign n13361_1 = ~P3_IR_REG_21_ & ~P3_IR_REG_22_;
  assign n13362 = n13359 & n13360;
  assign n13363 = n13361_1 & n13362;
  assign n13364 = n13269 & n13363;
  assign n13365 = ~n13358 & ~n13364;
  assign n13366_1 = n13116_1 & n13365;
  assign n911 = ~n13349 | n13366_1;
  assign n13368 = P3_IR_REG_23_ & n13112;
  assign n13369 = ~n13321_1 & ~n13368;
  assign n13370 = P3_IR_REG_23_ & ~n13364;
  assign n13371_1 = ~P3_IR_REG_7_ & ~P3_IR_REG_9_;
  assign n13372 = ~P3_IR_REG_8_ & n13371_1;
  assign n13373 = ~P3_IR_REG_4_ & ~P3_IR_REG_6_;
  assign n13374 = ~P3_IR_REG_5_ & n13373;
  assign n13375 = ~P3_IR_REG_3_ & ~P3_IR_REG_23_;
  assign n13376_1 = ~P3_IR_REG_2_ & n13375;
  assign n13377 = ~P3_IR_REG_20_ & ~P3_IR_REG_22_;
  assign n13378 = ~P3_IR_REG_21_ & n13377;
  assign n13379 = n13372 & n13374;
  assign n13380 = n13376_1 & n13379;
  assign n13381_1 = n13378 & n13380;
  assign n13382 = ~P3_IR_REG_0_ & ~P3_IR_REG_19_;
  assign n13383 = ~P3_IR_REG_1_ & n13382;
  assign n13384 = ~P3_IR_REG_16_ & ~P3_IR_REG_18_;
  assign n13385 = ~P3_IR_REG_17_ & n13384;
  assign n13386_1 = n13383 & n13385;
  assign n13387 = n13325 & n13386_1;
  assign n13388 = n13327 & n13387;
  assign n13389 = n13381_1 & n13388;
  assign n13390 = ~n13370 & ~n13389;
  assign n13391_1 = n13116_1 & n13390;
  assign n916 = ~n13369 | n13391_1;
  assign n13393 = P3_IR_REG_24_ & n13112;
  assign n13394 = ~n13321_1 & ~n13393;
  assign n13395 = P3_IR_REG_24_ & ~n13389;
  assign n13396_1 = ~P3_IR_REG_3_ & ~P3_IR_REG_24_;
  assign n13397 = ~P3_IR_REG_2_ & n13396_1;
  assign n13398 = ~P3_IR_REG_21_ & ~P3_IR_REG_23_;
  assign n13399 = ~P3_IR_REG_22_ & n13398;
  assign n13400 = n13379 & n13397;
  assign n13401_1 = n13399 & n13400;
  assign n13402 = ~P3_IR_REG_1_ & ~P3_IR_REG_20_;
  assign n13403 = ~P3_IR_REG_0_ & n13402;
  assign n13404 = ~P3_IR_REG_17_ & ~P3_IR_REG_19_;
  assign n13405 = ~P3_IR_REG_18_ & n13404;
  assign n13406_1 = ~P3_IR_REG_14_ & ~P3_IR_REG_16_;
  assign n13407 = ~P3_IR_REG_15_ & n13406_1;
  assign n13408 = ~P3_IR_REG_13_ & n13220;
  assign n13409 = n13403 & n13405;
  assign n13410 = n13407 & n13409;
  assign n13411_1 = n13408 & n13410;
  assign n13412 = n13401_1 & n13411_1;
  assign n13413 = ~n13395 & ~n13412;
  assign n13414 = n13116_1 & n13413;
  assign n921 = ~n13394 | n13414;
  assign n13416_1 = P3_IR_REG_25_ & n13112;
  assign n13417 = ~n13321_1 & ~n13416_1;
  assign n13418 = ~P3_IR_REG_25_ & n13412;
  assign n13419 = P3_IR_REG_25_ & ~n13412;
  assign n13420 = ~n13418 & ~n13419;
  assign n13421_1 = n13116_1 & n13420;
  assign n926 = ~n13417 | n13421_1;
  assign n13423 = P3_IR_REG_26_ & n13112;
  assign n13424 = ~n13321_1 & ~n13423;
  assign n13425 = ~P3_IR_REG_3_ & ~P3_IR_REG_25_;
  assign n13426_1 = ~P3_IR_REG_2_ & n13425;
  assign n13427 = ~P3_IR_REG_23_ & n13361_1;
  assign n13428 = ~P3_IR_REG_24_ & n13427;
  assign n13429 = n13379 & n13426_1;
  assign n13430 = n13428 & n13429;
  assign n13431_1 = n13411_1 & n13430;
  assign n13432 = P3_IR_REG_26_ & ~n13431_1;
  assign n13433 = ~P3_IR_REG_3_ & ~P3_IR_REG_26_;
  assign n13434 = ~P3_IR_REG_2_ & n13433;
  assign n13435 = ~P3_IR_REG_22_ & ~P3_IR_REG_23_;
  assign n13436_1 = ~P3_IR_REG_24_ & n13435;
  assign n13437 = ~P3_IR_REG_25_ & n13436_1;
  assign n13438 = n13379 & n13434;
  assign n13439 = n13437 & n13438;
  assign n13440 = ~P3_IR_REG_19_ & n13360;
  assign n13441_1 = ~P3_IR_REG_1_ & n13440;
  assign n13442 = n13353 & n13441_1;
  assign n13443 = n13407 & n13442;
  assign n13444 = n13408 & n13443;
  assign n13445 = n13439 & n13444;
  assign n13446_1 = ~n13432 & ~n13445;
  assign n13447 = n13116_1 & n13446_1;
  assign n931 = ~n13424 | n13447;
  assign n13449 = P3_IR_REG_27_ & n13112;
  assign n13450 = ~n13321_1 & ~n13449;
  assign n13451_1 = ~P3_IR_REG_27_ & ~n13445;
  assign n13452 = P3_IR_REG_27_ & n13445;
  assign n13453 = ~n13451_1 & ~n13452;
  assign n13454 = n13116_1 & ~n13453;
  assign n936 = ~n13450 | n13454;
  assign n13456_1 = P3_IR_REG_28_ & n13112;
  assign n13457 = ~n13321_1 & ~n13456_1;
  assign n13458 = ~P3_IR_REG_2_ & ~P3_IR_REG_26_;
  assign n13459 = ~P3_IR_REG_27_ & n13458;
  assign n13460 = n13184 & n13372;
  assign n13461_1 = n13459 & n13460;
  assign n13462 = n13437 & n13461_1;
  assign n13463 = n13444 & n13462;
  assign n13464 = P3_IR_REG_28_ & ~n13463;
  assign n13465 = ~P3_IR_REG_2_ & ~P3_IR_REG_27_;
  assign n13466_1 = ~P3_IR_REG_28_ & n13465;
  assign n13467 = ~P3_IR_REG_23_ & ~P3_IR_REG_24_;
  assign n13468 = ~P3_IR_REG_25_ & n13467;
  assign n13469 = ~P3_IR_REG_26_ & n13468;
  assign n13470 = n13460 & n13466_1;
  assign n13471_1 = n13469 & n13470;
  assign n13472 = ~P3_IR_REG_1_ & n13310;
  assign n13473 = ~P3_IR_REG_0_ & n13472;
  assign n13474 = ~P3_IR_REG_14_ & ~P3_IR_REG_15_;
  assign n13475 = ~P3_IR_REG_16_ & n13474;
  assign n13476_1 = ~P3_IR_REG_17_ & n13475;
  assign n13477 = n13378 & n13473;
  assign n13478 = n13476_1 & n13477;
  assign n13479 = n13408 & n13478;
  assign n13480 = n13471_1 & n13479;
  assign n13481_1 = ~n13464 & ~n13480;
  assign n13482 = n13116_1 & n13481_1;
  assign n941 = ~n13457 | n13482;
  assign n13484 = P3_IR_REG_29_ & n13112;
  assign n13485 = ~n13321_1 & ~n13484;
  assign n13486_1 = P3_IR_REG_29_ & ~n13480;
  assign n13487 = ~P3_IR_REG_27_ & ~P3_IR_REG_28_;
  assign n13488 = ~P3_IR_REG_29_ & n13487;
  assign n13489 = ~P3_IR_REG_2_ & n13488;
  assign n13490 = n13460 & n13489;
  assign n13491_1 = n13469 & n13490;
  assign n13492 = n13479 & n13491_1;
  assign n13493 = ~n13486_1 & ~n13492;
  assign n13494 = n13116_1 & n13493;
  assign n946 = ~n13485 | n13494;
  assign n13496_1 = P3_IR_REG_30_ & n13112;
  assign n13497 = ~n13321_1 & ~n13496_1;
  assign n13498 = ~P3_IR_REG_30_ & n13492;
  assign n13499 = P3_IR_REG_30_ & ~n13492;
  assign n13500 = ~n13498 & ~n13499;
  assign n13501_1 = n13116_1 & n13500;
  assign n951 = ~n13497 | n13501_1;
  assign n13503 = P3_IR_REG_31_ & n13112;
  assign n13504 = ~n13321_1 & ~n13503;
  assign n13505 = P3_IR_REG_31_ & n13498;
  assign n13506_1 = ~P3_IR_REG_31_ & ~n13498;
  assign n13507 = ~n13505 & ~n13506_1;
  assign n13508 = n13116_1 & ~n13507;
  assign n956 = ~n13504 | n13508;
  assign n13510 = P3_IR_REG_31_ & n13390;
  assign n13511_1 = P3_IR_REG_23_ & ~P3_IR_REG_31_;
  assign n13512 = ~n13510 & ~n13511_1;
  assign n13513 = P3_IR_REG_31_ & n13413;
  assign n13514 = P3_IR_REG_24_ & ~P3_IR_REG_31_;
  assign n13515 = ~n13513 & ~n13514;
  assign n13516_1 = P3_IR_REG_31_ & n13446_1;
  assign n13517 = P3_IR_REG_26_ & ~P3_IR_REG_31_;
  assign n13518 = ~n13516_1 & ~n13517;
  assign n13519 = ~n13515 & ~n13518;
  assign n13520 = P3_IR_REG_31_ & n13420;
  assign n13521_1 = P3_IR_REG_25_ & ~P3_IR_REG_31_;
  assign n13522 = ~n13520 & ~n13521_1;
  assign n13523 = n13519 & ~n13522;
  assign n13524 = n13512 & ~n13523;
  assign n13525 = P3_STATE_REG & n13524;
  assign n13526_1 = ~n13518 & n13522;
  assign n13527 = n13515 & n13526_1;
  assign n13528 = P3_B_REG & n13527;
  assign n13529 = ~P3_B_REG & n13519;
  assign n13530 = ~n13528 & ~n13529;
  assign n13531_1 = ~n13518 & n13530;
  assign n13532 = n13525 & ~n13531_1;
  assign n13533 = n13515 & ~n13526_1;
  assign n13534 = n13532 & ~n13533;
  assign n13535 = P3_D_REG_0_ & ~n13532;
  assign n961 = n13534 | n13535;
  assign n13537 = n13522 & ~n13526_1;
  assign n13538 = n13532 & ~n13537;
  assign n13539 = P3_D_REG_1_ & ~n13532;
  assign n966 = n13538 | n13539;
  assign n971 = P3_D_REG_2_ & ~n13532;
  assign n976 = P3_D_REG_3_ & ~n13532;
  assign n981 = P3_D_REG_4_ & ~n13532;
  assign n986 = P3_D_REG_5_ & ~n13532;
  assign n991 = P3_D_REG_6_ & ~n13532;
  assign n996 = P3_D_REG_7_ & ~n13532;
  assign n1001 = P3_D_REG_8_ & ~n13532;
  assign n1006 = P3_D_REG_9_ & ~n13532;
  assign n1011 = P3_D_REG_10_ & ~n13532;
  assign n1016 = P3_D_REG_11_ & ~n13532;
  assign n1021 = P3_D_REG_12_ & ~n13532;
  assign n1026 = P3_D_REG_13_ & ~n13532;
  assign n1031 = P3_D_REG_14_ & ~n13532;
  assign n1036 = P3_D_REG_15_ & ~n13532;
  assign n1041 = P3_D_REG_16_ & ~n13532;
  assign n1046 = P3_D_REG_17_ & ~n13532;
  assign n1051 = P3_D_REG_18_ & ~n13532;
  assign n1056 = P3_D_REG_19_ & ~n13532;
  assign n1061 = P3_D_REG_20_ & ~n13532;
  assign n1066 = P3_D_REG_21_ & ~n13532;
  assign n1071 = P3_D_REG_22_ & ~n13532;
  assign n1076 = P3_D_REG_23_ & ~n13532;
  assign n1081 = P3_D_REG_24_ & ~n13532;
  assign n1086 = P3_D_REG_25_ & ~n13532;
  assign n1091 = P3_D_REG_26_ & ~n13532;
  assign n1096 = P3_D_REG_27_ & ~n13532;
  assign n1101 = P3_D_REG_28_ & ~n13532;
  assign n1106 = P3_D_REG_29_ & ~n13532;
  assign n1111 = P3_D_REG_30_ & ~n13532;
  assign n1116 = P3_D_REG_31_ & ~n13532;
  assign n13571_1 = P3_D_REG_0_ & n13531_1;
  assign n13572 = n13515 & n13518;
  assign n13573 = ~n13531_1 & ~n13572;
  assign n13574 = ~n13571_1 & ~n13573;
  assign n13575 = n13525 & n13574;
  assign n13576_1 = ~n13531_1 & ~n13537;
  assign n13577 = P3_D_REG_1_ & n13531_1;
  assign n13578 = ~n13576_1 & ~n13577;
  assign n13579 = P3_IR_REG_31_ & n13365;
  assign n13580 = P3_IR_REG_22_ & ~P3_IR_REG_31_;
  assign n13581_1 = ~n13579 & ~n13580;
  assign n13582 = P3_IR_REG_31_ & n13338;
  assign n13583 = P3_IR_REG_20_ & ~P3_IR_REG_31_;
  assign n13584 = ~n13582 & ~n13583;
  assign n13585 = P3_IR_REG_31_ & n13345;
  assign n13586_1 = P3_IR_REG_21_ & ~P3_IR_REG_31_;
  assign n13587 = ~n13585 & ~n13586_1;
  assign n13588 = n13584 & n13587;
  assign n13589 = n13581_1 & ~n13588;
  assign n13590 = ~n13581_1 & n13587;
  assign n13591_1 = P3_IR_REG_31_ & n13317;
  assign n13592 = P3_IR_REG_19_ & ~P3_IR_REG_31_;
  assign n13593 = ~n13591_1 & ~n13592;
  assign n13594 = n13584 & n13593;
  assign n13595 = ~n13589 & ~n13590;
  assign n13596_1 = ~n13594 & n13595;
  assign n13597 = n13578 & ~n13596_1;
  assign n13598 = P3_D_REG_8_ & n13531_1;
  assign n13599 = P3_D_REG_7_ & n13531_1;
  assign n13600 = P3_D_REG_9_ & n13531_1;
  assign n13601_1 = ~n13598 & ~n13599;
  assign n13602 = ~n13600 & n13601_1;
  assign n13603 = P3_D_REG_6_ & n13531_1;
  assign n13604 = P3_D_REG_5_ & n13531_1;
  assign n13605 = P3_D_REG_4_ & n13531_1;
  assign n13606_1 = P3_D_REG_3_ & n13531_1;
  assign n13607 = ~n13603 & ~n13604;
  assign n13608 = ~n13605 & n13607;
  assign n13609 = ~n13606_1 & n13608;
  assign n13610 = P3_D_REG_31_ & n13531_1;
  assign n13611_1 = P3_D_REG_30_ & n13531_1;
  assign n13612 = P3_D_REG_2_ & n13531_1;
  assign n13613 = P3_D_REG_29_ & n13531_1;
  assign n13614 = ~n13610 & ~n13611_1;
  assign n13615 = ~n13612 & n13614;
  assign n13616_1 = ~n13613 & n13615;
  assign n13617 = P3_D_REG_28_ & n13531_1;
  assign n13618 = P3_D_REG_27_ & n13531_1;
  assign n13619 = P3_D_REG_26_ & n13531_1;
  assign n13620 = P3_D_REG_25_ & n13531_1;
  assign n13621_1 = ~n13617 & ~n13618;
  assign n13622 = ~n13619 & n13621_1;
  assign n13623 = ~n13620 & n13622;
  assign n13624 = n13602 & n13609;
  assign n13625 = n13616_1 & n13624;
  assign n13626_1 = n13623 & n13625;
  assign n13627 = P3_D_REG_23_ & n13531_1;
  assign n13628 = P3_D_REG_22_ & n13531_1;
  assign n13629 = P3_D_REG_24_ & n13531_1;
  assign n13630 = ~n13627 & ~n13628;
  assign n13631_1 = ~n13629 & n13630;
  assign n13632 = P3_D_REG_21_ & n13531_1;
  assign n13633 = P3_D_REG_20_ & n13531_1;
  assign n13634 = P3_D_REG_19_ & n13531_1;
  assign n13635 = P3_D_REG_18_ & n13531_1;
  assign n13636_1 = ~n13632 & ~n13633;
  assign n13637 = ~n13634 & n13636_1;
  assign n13638 = ~n13635 & n13637;
  assign n13639 = P3_D_REG_17_ & n13531_1;
  assign n13640 = P3_D_REG_16_ & n13531_1;
  assign n13641_1 = P3_D_REG_15_ & n13531_1;
  assign n13642 = P3_D_REG_14_ & n13531_1;
  assign n13643 = ~n13639 & ~n13640;
  assign n13644 = ~n13641_1 & n13643;
  assign n13645 = ~n13642 & n13644;
  assign n13646_1 = P3_D_REG_13_ & n13531_1;
  assign n13647 = P3_D_REG_12_ & n13531_1;
  assign n13648 = P3_D_REG_11_ & n13531_1;
  assign n13649 = P3_D_REG_10_ & n13531_1;
  assign n13650 = ~n13646_1 & ~n13647;
  assign n13651_1 = ~n13648 & n13650;
  assign n13652 = ~n13649 & n13651_1;
  assign n13653 = n13631_1 & n13638;
  assign n13654 = n13645 & n13653;
  assign n13655 = n13652 & n13654;
  assign n13656_1 = n13626_1 & n13655;
  assign n13657 = n13597 & n13656_1;
  assign n13658 = n13575 & n13657;
  assign n13659 = P3_IR_REG_31_ & ~n13453;
  assign n13660 = P3_IR_REG_27_ & ~P3_IR_REG_31_;
  assign n13661_1 = ~n13659 & ~n13660;
  assign n13662 = P3_IR_REG_31_ & n13481_1;
  assign n13663 = P3_IR_REG_28_ & ~P3_IR_REG_31_;
  assign n13664 = ~n13662 & ~n13663;
  assign n13665 = n13661_1 & n13664;
  assign n13666_1 = P3_IR_REG_0_ & P3_IR_REG_31_;
  assign n13667 = P3_IR_REG_0_ & ~P3_IR_REG_31_;
  assign n13668 = ~n13666_1 & ~n13667;
  assign n13669 = n13665 & ~n13668;
  assign n13670 = P1_P3_DATAO_REG_0_ & ~n13665;
  assign n13671_1 = ~n13669 & ~n13670;
  assign n13672 = n13581_1 & n13587;
  assign n13673 = ~n13584 & n13593;
  assign n13674 = n13672 & n13673;
  assign n13675 = n13581_1 & ~n13593;
  assign n13676_1 = n13587 & n13675;
  assign n13677 = ~n13674 & ~n13676_1;
  assign n13678 = ~n13671_1 & ~n13677;
  assign n13679 = ~n13581_1 & ~n13587;
  assign n13680 = n13664 & n13679;
  assign n13681_1 = P3_IR_REG_31_ & n13500;
  assign n13682 = P3_IR_REG_30_ & ~P3_IR_REG_31_;
  assign n13683 = ~n13681_1 & ~n13682;
  assign n13684 = P3_IR_REG_31_ & n13493;
  assign n13685 = P3_IR_REG_29_ & ~P3_IR_REG_31_;
  assign n13686_1 = ~n13684 & ~n13685;
  assign n13687 = ~n13683 & ~n13686_1;
  assign n13688 = P3_REG3_REG_1_ & n13687;
  assign n13689 = n13683 & n13686_1;
  assign n13690 = P3_REG0_REG_1_ & n13689;
  assign n13691_1 = n13683 & ~n13686_1;
  assign n13692 = P3_REG1_REG_1_ & n13691_1;
  assign n13693 = ~n13683 & n13686_1;
  assign n13694 = P3_REG2_REG_1_ & n13693;
  assign n13695 = ~n13688 & ~n13690;
  assign n13696_1 = ~n13692 & n13695;
  assign n13697 = ~n13694 & n13696_1;
  assign n13698 = n13680 & ~n13697;
  assign n13699 = n13584 & n13672;
  assign n13700 = ~n13671_1 & n13699;
  assign n13701_1 = P3_REG3_REG_0_ & n13687;
  assign n13702 = P3_REG2_REG_0_ & n13693;
  assign n13703 = P3_REG1_REG_0_ & n13691_1;
  assign n13704 = P3_REG0_REG_0_ & n13689;
  assign n13705 = ~n13701_1 & ~n13702;
  assign n13706_1 = ~n13703 & n13705;
  assign n13707 = ~n13704 & n13706_1;
  assign n13708 = ~n13671_1 & n13707;
  assign n13709 = n13671_1 & ~n13707;
  assign n13710 = ~n13708 & ~n13709;
  assign n13711_1 = n13584 & n13675;
  assign n13712 = ~n13710 & n13711_1;
  assign n13713 = ~n13700 & ~n13712;
  assign n13714 = ~n13678 & ~n13698;
  assign n13715 = n13713 & n13714;
  assign n13716_1 = ~n13581_1 & n13594;
  assign n13717 = n13587 & n13716_1;
  assign n13718 = ~n13710 & n13717;
  assign n13719 = ~n13587 & n13673;
  assign n13720 = ~n13710 & n13719;
  assign n13721_1 = ~n13587 & n13594;
  assign n13722 = n13581_1 & n13721_1;
  assign n13723 = ~n13710 & n13722;
  assign n13724 = ~n13584 & ~n13593;
  assign n13725 = ~n13587 & n13724;
  assign n13726_1 = ~n13710 & n13725;
  assign n13727 = ~n13581_1 & n13673;
  assign n13728 = ~n13710 & n13727;
  assign n13729 = ~n13726_1 & ~n13728;
  assign n13730 = ~n13581_1 & n13724;
  assign n13731_1 = ~n13710 & n13730;
  assign n13732 = n13584 & ~n13593;
  assign n13733 = ~n13581_1 & n13732;
  assign n13734 = ~n13710 & n13733;
  assign n13735 = ~n13731_1 & ~n13734;
  assign n13736_1 = ~n13718 & ~n13720;
  assign n13737 = ~n13723 & n13736_1;
  assign n13738 = n13729 & n13737;
  assign n13739 = n13735 & n13738;
  assign n13740 = n13715 & n13739;
  assign n13741_1 = n13658 & ~n13740;
  assign n13742 = P3_REG0_REG_0_ & ~n13658;
  assign n1121 = n13741_1 | n13742;
  assign n13744 = P3_REG3_REG_2_ & n13687;
  assign n13745 = P3_REG0_REG_2_ & n13689;
  assign n13746_1 = P3_REG1_REG_2_ & n13691_1;
  assign n13747 = P3_REG2_REG_2_ & n13693;
  assign n13748 = ~n13744 & ~n13745;
  assign n13749 = ~n13746_1 & n13748;
  assign n13750 = ~n13747 & n13749;
  assign n13751_1 = n13680 & ~n13750;
  assign n13752 = P3_IR_REG_31_ & ~n13124;
  assign n13753 = P3_IR_REG_1_ & ~P3_IR_REG_31_;
  assign n13754 = ~n13752 & ~n13753;
  assign n13755 = n13665 & ~n13754;
  assign n13756_1 = P1_P3_DATAO_REG_1_ & ~n13665;
  assign n13757 = ~n13755 & ~n13756_1;
  assign n13758 = ~n13671_1 & n13757;
  assign n13759 = n13671_1 & ~n13757;
  assign n13760 = ~n13758 & ~n13759;
  assign n13761_1 = n13699 & ~n13760;
  assign n13762 = ~n13677 & ~n13757;
  assign n13763 = ~n13697 & ~n13757;
  assign n13764 = n13697 & n13757;
  assign n13765 = ~n13763 & ~n13764;
  assign n13766_1 = ~n13671_1 & ~n13707;
  assign n13767 = n13765 & ~n13766_1;
  assign n13768 = ~n13765 & n13766_1;
  assign n13769 = ~n13767 & ~n13768;
  assign n13770 = n13711_1 & ~n13769;
  assign n13771_1 = ~n13751_1 & ~n13761_1;
  assign n13772 = ~n13762 & n13771_1;
  assign n13773 = ~n13770 & n13772;
  assign n13774 = ~n13697 & n13757;
  assign n13775 = n13697 & ~n13757;
  assign n13776_1 = ~n13774 & ~n13775;
  assign n13777 = ~n13708 & ~n13776_1;
  assign n13778 = n13708 & n13776_1;
  assign n13779 = ~n13777 & ~n13778;
  assign n13780 = n13733 & ~n13779;
  assign n13781_1 = ~n13664 & n13679;
  assign n13782 = ~n13707 & n13781_1;
  assign n13783 = n13727 & ~n13769;
  assign n13784 = n13730 & ~n13779;
  assign n13785 = ~n13783 & ~n13784;
  assign n13786_1 = n13722 & ~n13769;
  assign n13787 = n13717 & ~n13769;
  assign n13788 = n13719 & ~n13779;
  assign n13789 = n13725 & ~n13779;
  assign n13790 = ~n13788 & ~n13789;
  assign n13791_1 = ~n13786_1 & ~n13787;
  assign n13792 = n13790 & n13791_1;
  assign n13793 = ~n13780 & ~n13782;
  assign n13794 = n13785 & n13793;
  assign n13795 = n13792 & n13794;
  assign n13796_1 = n13773 & n13795;
  assign n13797 = n13658 & ~n13796_1;
  assign n13798 = P3_REG0_REG_1_ & ~n13658;
  assign n1126 = n13797 | n13798;
  assign n13800 = ~P3_REG3_REG_3_ & n13687;
  assign n13801_1 = P3_REG0_REG_3_ & n13689;
  assign n13802 = P3_REG1_REG_3_ & n13691_1;
  assign n13803 = P3_REG2_REG_3_ & n13693;
  assign n13804 = ~n13800 & ~n13801_1;
  assign n13805 = ~n13802 & n13804;
  assign n13806_1 = ~n13803 & n13805;
  assign n13807 = n13680 & ~n13806_1;
  assign n13808 = P3_IR_REG_31_ & n13133;
  assign n13809 = P3_IR_REG_2_ & ~P3_IR_REG_31_;
  assign n13810 = ~n13808 & ~n13809;
  assign n13811_1 = n13665 & ~n13810;
  assign n13812 = P1_P3_DATAO_REG_2_ & ~n13665;
  assign n13813 = ~n13811_1 & ~n13812;
  assign n13814 = n13671_1 & n13757;
  assign n13815 = ~n13813 & ~n13814;
  assign n13816_1 = n13813 & n13814;
  assign n13817 = ~n13815 & ~n13816_1;
  assign n13818 = n13699 & n13817;
  assign n13819 = ~n13677 & ~n13813;
  assign n13820 = ~n13750 & ~n13813;
  assign n13821_1 = n13750 & n13813;
  assign n13822 = ~n13820 & ~n13821_1;
  assign n13823 = ~n13764 & n13766_1;
  assign n13824 = ~n13763 & ~n13823;
  assign n13825 = n13822 & ~n13824;
  assign n13826_1 = n13750 & ~n13813;
  assign n13827 = ~n13750 & n13813;
  assign n13828 = ~n13826_1 & ~n13827;
  assign n13829 = ~n13763 & n13828;
  assign n13830 = ~n13823 & n13829;
  assign n13831_1 = ~n13825 & ~n13830;
  assign n13832 = n13711_1 & n13831_1;
  assign n13833 = ~n13807 & ~n13818;
  assign n13834 = ~n13819 & n13833;
  assign n13835 = ~n13832 & n13834;
  assign n13836_1 = ~n13697 & ~n13708;
  assign n13837 = n13697 & n13708;
  assign n13838 = n13757 & ~n13837;
  assign n13839 = ~n13836_1 & ~n13838;
  assign n13840 = n13828 & n13839;
  assign n13841_1 = ~n13828 & ~n13839;
  assign n13842 = ~n13840 & ~n13841_1;
  assign n13843 = n13733 & ~n13842;
  assign n13844 = ~n13697 & n13781_1;
  assign n13845 = n13727 & n13831_1;
  assign n13846_1 = n13730 & ~n13842;
  assign n13847 = ~n13845 & ~n13846_1;
  assign n13848 = n13722 & n13831_1;
  assign n13849 = n13717 & n13831_1;
  assign n13850 = n13719 & ~n13842;
  assign n13851_1 = n13725 & ~n13842;
  assign n13852 = ~n13850 & ~n13851_1;
  assign n13853 = ~n13848 & ~n13849;
  assign n13854 = n13852 & n13853;
  assign n13855 = ~n13843 & ~n13844;
  assign n13856_1 = n13847 & n13855;
  assign n13857 = n13854 & n13856_1;
  assign n13858 = n13835 & n13857;
  assign n13859 = n13658 & ~n13858;
  assign n13860 = P3_REG0_REG_2_ & ~n13658;
  assign n1131 = n13859 | n13860;
  assign n13862 = ~P3_REG3_REG_4_ & P3_REG3_REG_3_;
  assign n13863 = P3_REG3_REG_4_ & ~P3_REG3_REG_3_;
  assign n13864 = ~n13862 & ~n13863;
  assign n13865 = n13687 & ~n13864;
  assign n13866_1 = P3_REG0_REG_4_ & n13689;
  assign n13867 = P3_REG1_REG_4_ & n13691_1;
  assign n13868 = P3_REG2_REG_4_ & n13693;
  assign n13869 = ~n13865 & ~n13866_1;
  assign n13870 = ~n13867 & n13869;
  assign n13871_1 = ~n13868 & n13870;
  assign n13872 = n13680 & ~n13871_1;
  assign n13873 = P3_IR_REG_31_ & n13141_1;
  assign n13874 = P3_IR_REG_3_ & ~P3_IR_REG_31_;
  assign n13875 = ~n13873 & ~n13874;
  assign n13876_1 = n13665 & ~n13875;
  assign n13877 = P1_P3_DATAO_REG_3_ & ~n13665;
  assign n13878 = ~n13876_1 & ~n13877;
  assign n13879 = ~n13816_1 & ~n13878;
  assign n13880 = n13816_1 & n13878;
  assign n13881_1 = ~n13879 & ~n13880;
  assign n13882 = n13699 & n13881_1;
  assign n13883 = ~n13677 & ~n13878;
  assign n13884 = n13763 & ~n13821_1;
  assign n13885 = ~n13820 & ~n13884;
  assign n13886_1 = ~n13821_1 & n13823;
  assign n13887 = n13885 & ~n13886_1;
  assign n13888 = n13806_1 & ~n13878;
  assign n13889 = ~n13806_1 & n13878;
  assign n13890 = ~n13888 & ~n13889;
  assign n13891_1 = n13887 & ~n13890;
  assign n13892 = ~n13806_1 & ~n13878;
  assign n13893 = n13806_1 & n13878;
  assign n13894 = ~n13892 & ~n13893;
  assign n13895 = ~n13887 & ~n13894;
  assign n13896_1 = ~n13891_1 & ~n13895;
  assign n13897 = n13711_1 & ~n13896_1;
  assign n13898 = ~n13872 & ~n13882;
  assign n13899 = ~n13883 & n13898;
  assign n13900 = ~n13897 & n13899;
  assign n13901_1 = ~n13826_1 & ~n13890;
  assign n13902 = ~n13827 & n13839;
  assign n13903 = n13901_1 & ~n13902;
  assign n13904 = ~n13827 & n13890;
  assign n13905 = ~n13826_1 & ~n13839;
  assign n13906_1 = n13904 & ~n13905;
  assign n13907 = ~n13903 & ~n13906_1;
  assign n13908 = n13733 & ~n13907;
  assign n13909 = ~n13750 & n13781_1;
  assign n13910 = n13727 & ~n13896_1;
  assign n13911_1 = n13730 & ~n13907;
  assign n13912 = ~n13910 & ~n13911_1;
  assign n13913 = n13722 & ~n13896_1;
  assign n13914 = n13717 & ~n13896_1;
  assign n13915 = n13719 & ~n13907;
  assign n13916_1 = n13725 & ~n13907;
  assign n13917 = ~n13915 & ~n13916_1;
  assign n13918 = ~n13913 & ~n13914;
  assign n13919 = n13917 & n13918;
  assign n13920 = ~n13908 & ~n13909;
  assign n13921_1 = n13912 & n13920;
  assign n13922 = n13919 & n13921_1;
  assign n13923 = n13900 & n13922;
  assign n13924 = n13658 & ~n13923;
  assign n13925 = P3_REG0_REG_3_ & ~n13658;
  assign n1136 = n13924 | n13925;
  assign n13927 = P3_REG3_REG_4_ & P3_REG3_REG_3_;
  assign n13928 = ~P3_REG3_REG_5_ & n13927;
  assign n13929 = P3_REG3_REG_5_ & ~n13927;
  assign n13930 = ~n13928 & ~n13929;
  assign n13931_1 = n13687 & ~n13930;
  assign n13932 = P3_REG0_REG_5_ & n13689;
  assign n13933 = P3_REG1_REG_5_ & n13691_1;
  assign n13934 = P3_REG2_REG_5_ & n13693;
  assign n13935 = ~n13931_1 & ~n13932;
  assign n13936_1 = ~n13933 & n13935;
  assign n13937 = ~n13934 & n13936_1;
  assign n13938 = n13680 & ~n13937;
  assign n13939 = P3_IR_REG_31_ & n13150;
  assign n13940 = P3_IR_REG_4_ & ~P3_IR_REG_31_;
  assign n13941_1 = ~n13939 & ~n13940;
  assign n13942 = n13665 & ~n13941_1;
  assign n13943 = P1_P3_DATAO_REG_4_ & ~n13665;
  assign n13944 = ~n13942 & ~n13943;
  assign n13945 = ~n13880 & ~n13944;
  assign n13946_1 = n13880 & n13944;
  assign n13947 = ~n13945 & ~n13946_1;
  assign n13948 = n13699 & n13947;
  assign n13949 = ~n13677 & ~n13944;
  assign n13950 = n13871_1 & ~n13944;
  assign n13951_1 = ~n13871_1 & n13944;
  assign n13952 = ~n13950 & ~n13951_1;
  assign n13953 = ~n13821_1 & ~n13893;
  assign n13954 = n13823 & n13953;
  assign n13955 = ~n13892 & ~n13954;
  assign n13956_1 = ~n13885 & ~n13893;
  assign n13957 = n13955 & ~n13956_1;
  assign n13958 = ~n13952 & n13957;
  assign n13959 = n13871_1 & n13944;
  assign n13960 = ~n13871_1 & ~n13944;
  assign n13961_1 = ~n13959 & ~n13960;
  assign n13962 = ~n13957 & ~n13961_1;
  assign n13963 = ~n13958 & ~n13962;
  assign n13964 = n13711_1 & ~n13963;
  assign n13965 = ~n13938 & ~n13948;
  assign n13966_1 = ~n13949 & n13965;
  assign n13967 = ~n13964 & n13966_1;
  assign n13968 = n13806_1 & ~n13827;
  assign n13969 = n13878 & ~n13968;
  assign n13970 = ~n13806_1 & n13827;
  assign n13971_1 = ~n13969 & ~n13970;
  assign n13972 = ~n13826_1 & ~n13888;
  assign n13973 = ~n13839 & n13972;
  assign n13974 = n13971_1 & ~n13973;
  assign n13975 = n13952 & n13974;
  assign n13976_1 = ~n13952 & ~n13974;
  assign n13977 = ~n13975 & ~n13976_1;
  assign n13978 = n13733 & ~n13977;
  assign n13979 = n13781_1 & ~n13806_1;
  assign n13980 = n13727 & ~n13963;
  assign n13981_1 = n13730 & ~n13977;
  assign n13982 = ~n13980 & ~n13981_1;
  assign n13983 = n13722 & ~n13963;
  assign n13984 = n13717 & ~n13963;
  assign n13985 = n13719 & ~n13977;
  assign n13986_1 = n13725 & ~n13977;
  assign n13987 = ~n13985 & ~n13986_1;
  assign n13988 = ~n13983 & ~n13984;
  assign n13989 = n13987 & n13988;
  assign n13990 = ~n13978 & ~n13979;
  assign n13991_1 = n13982 & n13990;
  assign n13992 = n13989 & n13991_1;
  assign n13993 = n13967 & n13992;
  assign n13994 = n13658 & ~n13993;
  assign n13995 = P3_REG0_REG_4_ & ~n13658;
  assign n1141 = n13994 | n13995;
  assign n13997 = P3_REG3_REG_5_ & n13927;
  assign n13998 = ~P3_REG3_REG_6_ & n13997;
  assign n13999 = P3_REG3_REG_6_ & ~n13997;
  assign n14000 = ~n13998 & ~n13999;
  assign n14001_1 = n13687 & ~n14000;
  assign n14002 = P3_REG0_REG_6_ & n13689;
  assign n14003 = P3_REG1_REG_6_ & n13691_1;
  assign n14004 = P3_REG2_REG_6_ & n13693;
  assign n14005 = ~n14001_1 & ~n14002;
  assign n14006_1 = ~n14003 & n14005;
  assign n14007 = ~n14004 & n14006_1;
  assign n14008 = n13680 & ~n14007;
  assign n14009 = P3_IR_REG_31_ & n13158;
  assign n14010 = P3_IR_REG_5_ & ~P3_IR_REG_31_;
  assign n14011_1 = ~n14009 & ~n14010;
  assign n14012 = n13665 & ~n14011_1;
  assign n14013 = P1_P3_DATAO_REG_5_ & ~n13665;
  assign n14014 = ~n14012 & ~n14013;
  assign n14015 = ~n13946_1 & ~n14014;
  assign n14016_1 = n13946_1 & n14014;
  assign n14017 = ~n14015 & ~n14016_1;
  assign n14018 = n13699 & n14017;
  assign n14019 = ~n13677 & ~n14014;
  assign n14020 = ~n13937 & ~n14014;
  assign n14021_1 = n13937 & n14014;
  assign n14022 = ~n13959 & ~n14021_1;
  assign n14023 = ~n14020 & n14022;
  assign n14024 = n13957 & ~n13960;
  assign n14025 = n14023 & ~n14024;
  assign n14026_1 = n13937 & ~n14014;
  assign n14027 = ~n13937 & n14014;
  assign n14028 = ~n14026_1 & ~n14027;
  assign n14029 = ~n13960 & n14028;
  assign n14030 = ~n13957 & ~n13959;
  assign n14031_1 = n14029 & ~n14030;
  assign n14032 = ~n14025 & ~n14031_1;
  assign n14033 = n13711_1 & n14032;
  assign n14034 = ~n14008 & ~n14018;
  assign n14035 = ~n14019 & n14034;
  assign n14036_1 = ~n14033 & n14035;
  assign n14037 = ~n13950 & ~n13974;
  assign n14038 = ~n13951_1 & ~n14037;
  assign n14039 = n14028 & n14038;
  assign n14040 = ~n14028 & ~n14038;
  assign n14041_1 = ~n14039 & ~n14040;
  assign n14042 = n13733 & ~n14041_1;
  assign n14043 = n13781_1 & ~n13871_1;
  assign n14044 = n13727 & n14032;
  assign n14045 = n13730 & ~n14041_1;
  assign n14046_1 = ~n14044 & ~n14045;
  assign n14047 = n13722 & n14032;
  assign n14048 = n13717 & n14032;
  assign n14049 = n13719 & ~n14041_1;
  assign n14050 = n13725 & ~n14041_1;
  assign n14051_1 = ~n14049 & ~n14050;
  assign n14052 = ~n14047 & ~n14048;
  assign n14053 = n14051_1 & n14052;
  assign n14054 = ~n14042 & ~n14043;
  assign n14055 = n14046_1 & n14054;
  assign n14056_1 = n14053 & n14055;
  assign n14057 = n14036_1 & n14056_1;
  assign n14058 = n13658 & ~n14057;
  assign n14059 = P3_REG0_REG_5_ & ~n13658;
  assign n1146 = n14058 | n14059;
  assign n14061_1 = P3_IR_REG_31_ & n13167;
  assign n14062 = P3_IR_REG_6_ & ~P3_IR_REG_31_;
  assign n14063 = ~n14061_1 & ~n14062;
  assign n14064 = n13665 & ~n14063;
  assign n14065 = P1_P3_DATAO_REG_6_ & ~n13665;
  assign n14066_1 = ~n14064 & ~n14065;
  assign n14067 = ~n13677 & ~n14066_1;
  assign n14068 = n14007 & ~n14066_1;
  assign n14069 = ~n14007 & n14066_1;
  assign n14070 = ~n14068 & ~n14069;
  assign n14071_1 = n13960 & ~n14014;
  assign n14072 = ~n13960 & n14014;
  assign n14073 = ~n13937 & ~n14072;
  assign n14074 = ~n14071_1 & ~n14073;
  assign n14075 = n13820 & ~n13893;
  assign n14076_1 = ~n13892 & ~n14075;
  assign n14077 = ~n13824 & n13953;
  assign n14078 = n14076_1 & ~n14077;
  assign n14079 = n14022 & ~n14078;
  assign n14080 = n14074 & ~n14079;
  assign n14081_1 = ~n14070 & n14080;
  assign n14082 = n14007 & n14066_1;
  assign n14083 = ~n14007 & ~n14066_1;
  assign n14084 = ~n14082 & ~n14083;
  assign n14085 = ~n14080 & ~n14084;
  assign n14086_1 = ~n14081_1 & ~n14085;
  assign n14087 = n13711_1 & ~n14086_1;
  assign n14088 = P3_REG3_REG_6_ & n13997;
  assign n14089 = ~P3_REG3_REG_7_ & n14088;
  assign n14090 = P3_REG3_REG_7_ & ~n14088;
  assign n14091_1 = ~n14089 & ~n14090;
  assign n14092 = n13687 & ~n14091_1;
  assign n14093 = P3_REG0_REG_7_ & n13689;
  assign n14094 = P3_REG1_REG_7_ & n13691_1;
  assign n14095 = P3_REG2_REG_7_ & n13693;
  assign n14096_1 = ~n14092 & ~n14093;
  assign n14097 = ~n14094 & n14096_1;
  assign n14098 = ~n14095 & n14097;
  assign n14099 = n13680 & ~n14098;
  assign n14100 = ~n14016_1 & ~n14066_1;
  assign n14101_1 = n14016_1 & n14066_1;
  assign n14102 = ~n14100 & ~n14101_1;
  assign n14103 = n13699 & n14102;
  assign n14104 = ~n14067 & ~n14087;
  assign n14105 = ~n14099 & n14104;
  assign n14106_1 = ~n14103 & n14105;
  assign n14107 = ~n14026_1 & ~n14070;
  assign n14108 = ~n14027 & n14038;
  assign n14109 = n14107 & ~n14108;
  assign n14110 = ~n14027 & ~n14069;
  assign n14111_1 = ~n14068 & n14110;
  assign n14112 = ~n14026_1 & ~n14038;
  assign n14113 = n14111_1 & ~n14112;
  assign n14114 = ~n14109 & ~n14113;
  assign n14115 = n13733 & ~n14114;
  assign n14116_1 = n13781_1 & ~n13937;
  assign n14117 = n13727 & ~n14086_1;
  assign n14118 = n13730 & ~n14114;
  assign n14119 = ~n14117 & ~n14118;
  assign n14120 = n13722 & ~n14086_1;
  assign n14121_1 = n13717 & ~n14086_1;
  assign n14122 = n13719 & ~n14114;
  assign n14123 = n13725 & ~n14114;
  assign n14124 = ~n14122 & ~n14123;
  assign n14125 = ~n14120 & ~n14121_1;
  assign n14126_1 = n14124 & n14125;
  assign n14127 = ~n14115 & ~n14116_1;
  assign n14128 = n14119 & n14127;
  assign n14129 = n14126_1 & n14128;
  assign n14130 = n14106_1 & n14129;
  assign n14131_1 = n13658 & ~n14130;
  assign n14132 = P3_REG0_REG_6_ & ~n13658;
  assign n1151 = n14131_1 | n14132;
  assign n14134 = P3_IR_REG_31_ & n13175;
  assign n14135 = P3_IR_REG_7_ & ~P3_IR_REG_31_;
  assign n14136_1 = ~n14134 & ~n14135;
  assign n14137 = n13665 & ~n14136_1;
  assign n14138 = P1_P3_DATAO_REG_7_ & ~n13665;
  assign n14139 = ~n14137 & ~n14138;
  assign n14140 = ~n13677 & ~n14139;
  assign n14141_1 = ~n14098 & ~n14139;
  assign n14142 = n14098 & n14139;
  assign n14143 = ~n14082 & ~n14142;
  assign n14144 = ~n14141_1 & n14143;
  assign n14145 = n14080 & ~n14083;
  assign n14146_1 = n14144 & ~n14145;
  assign n14147 = n14098 & ~n14139;
  assign n14148 = ~n14098 & n14139;
  assign n14149 = ~n14147 & ~n14148;
  assign n14150 = ~n14083 & n14149;
  assign n14151_1 = ~n14080 & ~n14082;
  assign n14152 = n14150 & ~n14151_1;
  assign n14153 = ~n14146_1 & ~n14152;
  assign n14154 = n13711_1 & n14153;
  assign n14155 = P3_REG3_REG_7_ & n14088;
  assign n14156_1 = ~P3_REG3_REG_8_ & n14155;
  assign n14157 = P3_REG3_REG_8_ & ~n14155;
  assign n14158 = ~n14156_1 & ~n14157;
  assign n14159 = n13687 & ~n14158;
  assign n14160 = P3_REG0_REG_8_ & n13689;
  assign n14161_1 = P3_REG1_REG_8_ & n13691_1;
  assign n14162 = P3_REG2_REG_8_ & n13693;
  assign n14163 = ~n14159 & ~n14160;
  assign n14164 = ~n14161_1 & n14163;
  assign n14165 = ~n14162 & n14164;
  assign n14166_1 = n13680 & ~n14165;
  assign n14167 = ~n14101_1 & ~n14139;
  assign n14168 = n14101_1 & n14139;
  assign n14169 = ~n14167 & ~n14168;
  assign n14170 = n13699 & n14169;
  assign n14171_1 = ~n14140 & ~n14154;
  assign n14172 = ~n14166_1 & n14171_1;
  assign n14173 = ~n14170 & n14172;
  assign n14174 = ~n14026_1 & ~n14068;
  assign n14175 = n13951_1 & n14174;
  assign n14176_1 = n14110 & ~n14175;
  assign n14177 = ~n14068 & ~n14176_1;
  assign n14178 = ~n13950 & n14174;
  assign n14179 = ~n13974 & n14178;
  assign n14180 = ~n14177 & ~n14179;
  assign n14181_1 = n14149 & n14180;
  assign n14182 = ~n14149 & ~n14180;
  assign n14183 = ~n14181_1 & ~n14182;
  assign n14184 = n13733 & ~n14183;
  assign n14185 = n13781_1 & ~n14007;
  assign n14186_1 = n13727 & n14153;
  assign n14187 = n13730 & ~n14183;
  assign n14188 = ~n14186_1 & ~n14187;
  assign n14189 = n13722 & n14153;
  assign n14190 = n13717 & n14153;
  assign n14191_1 = n13719 & ~n14183;
  assign n14192 = n13725 & ~n14183;
  assign n14193 = ~n14191_1 & ~n14192;
  assign n14194 = ~n14189 & ~n14190;
  assign n14195 = n14193 & n14194;
  assign n14196_1 = ~n14184 & ~n14185;
  assign n14197 = n14188 & n14196_1;
  assign n14198 = n14195 & n14197;
  assign n14199 = n14173 & n14198;
  assign n14200 = n13658 & ~n14199;
  assign n14201_1 = P3_REG0_REG_7_ & ~n13658;
  assign n1156 = n14200 | n14201_1;
  assign n14203 = P3_IR_REG_31_ & n13187;
  assign n14204 = P3_IR_REG_8_ & ~P3_IR_REG_31_;
  assign n14205 = ~n14203 & ~n14204;
  assign n14206_1 = n13665 & ~n14205;
  assign n14207 = P1_P3_DATAO_REG_8_ & ~n13665;
  assign n14208 = ~n14206_1 & ~n14207;
  assign n14209 = ~n13677 & ~n14208;
  assign n14210 = n14168 & n14208;
  assign n14211_1 = ~n14168 & ~n14208;
  assign n14212 = ~n14210 & ~n14211_1;
  assign n14213 = n13699 & n14212;
  assign n14214 = P3_REG1_REG_9_ & n13691_1;
  assign n14215 = P3_REG0_REG_9_ & n13689;
  assign n14216_1 = P3_REG2_REG_9_ & n13693;
  assign n14217 = P3_REG3_REG_8_ & n14155;
  assign n14218 = ~P3_REG3_REG_9_ & n14217;
  assign n14219 = P3_REG3_REG_9_ & ~n14217;
  assign n14220 = ~n14218 & ~n14219;
  assign n14221_1 = n13687 & ~n14220;
  assign n14222 = ~n14214 & ~n14215;
  assign n14223 = ~n14216_1 & n14222;
  assign n14224 = ~n14221_1 & n14223;
  assign n14225 = n13680 & ~n14224;
  assign n14226_1 = n14083 & ~n14139;
  assign n14227 = ~n14083 & n14139;
  assign n14228 = ~n14098 & ~n14227;
  assign n14229 = ~n14226_1 & ~n14228;
  assign n14230 = ~n14080 & n14143;
  assign n14231_1 = n14229 & ~n14230;
  assign n14232 = n14165 & ~n14208;
  assign n14233 = ~n14165 & n14208;
  assign n14234 = ~n14232 & ~n14233;
  assign n14235 = n14231_1 & ~n14234;
  assign n14236_1 = n14165 & n14208;
  assign n14237 = ~n14165 & ~n14208;
  assign n14238 = ~n14236_1 & ~n14237;
  assign n14239 = ~n14231_1 & ~n14238;
  assign n14240 = ~n14235 & ~n14239;
  assign n14241_1 = n13711_1 & ~n14240;
  assign n14242 = ~n14209 & ~n14213;
  assign n14243 = ~n14225 & n14242;
  assign n14244 = ~n14241_1 & n14243;
  assign n14245 = ~n14147 & ~n14234;
  assign n14246_1 = ~n14148 & n14180;
  assign n14247 = n14245 & ~n14246_1;
  assign n14248 = ~n14148 & n14234;
  assign n14249 = ~n14147 & ~n14180;
  assign n14250 = n14248 & ~n14249;
  assign n14251_1 = ~n14247 & ~n14250;
  assign n14252 = n13733 & ~n14251_1;
  assign n14253 = n13781_1 & ~n14098;
  assign n14254 = n13727 & ~n14240;
  assign n14255 = n13730 & ~n14251_1;
  assign n14256_1 = ~n14254 & ~n14255;
  assign n14257 = n13722 & ~n14240;
  assign n14258 = n13717 & ~n14240;
  assign n14259 = n13719 & ~n14251_1;
  assign n14260 = n13725 & ~n14251_1;
  assign n14261_1 = ~n14259 & ~n14260;
  assign n14262 = ~n14257 & ~n14258;
  assign n14263 = n14261_1 & n14262;
  assign n14264 = ~n14252 & ~n14253;
  assign n14265 = n14256_1 & n14264;
  assign n14266_1 = n14263 & n14265;
  assign n14267 = n14244 & n14266_1;
  assign n14268 = n13658 & ~n14267;
  assign n14269 = P3_REG0_REG_8_ & ~n13658;
  assign n1161 = n14268 | n14269;
  assign n14271_1 = P3_IR_REG_31_ & n13195;
  assign n14272 = P3_IR_REG_9_ & ~P3_IR_REG_31_;
  assign n14273 = ~n14271_1 & ~n14272;
  assign n14274 = n13665 & ~n14273;
  assign n14275 = P1_P3_DATAO_REG_9_ & ~n13665;
  assign n14276_1 = ~n14274 & ~n14275;
  assign n14277 = ~n13677 & ~n14276_1;
  assign n14278 = n14210 & n14276_1;
  assign n14279 = ~n14210 & ~n14276_1;
  assign n14280 = ~n14278 & ~n14279;
  assign n14281_1 = n13699 & n14280;
  assign n14282 = P3_REG1_REG_10_ & n13691_1;
  assign n14283 = P3_REG0_REG_10_ & n13689;
  assign n14284 = P3_REG2_REG_10_ & n13693;
  assign n14285 = P3_REG3_REG_9_ & n14217;
  assign n14286_1 = ~P3_REG3_REG_10_ & n14285;
  assign n14287 = P3_REG3_REG_10_ & ~n14285;
  assign n14288 = ~n14286_1 & ~n14287;
  assign n14289 = n13687 & ~n14288;
  assign n14290 = ~n14282 & ~n14283;
  assign n14291_1 = ~n14284 & n14290;
  assign n14292 = ~n14289 & n14291_1;
  assign n14293 = n13680 & ~n14292;
  assign n14294 = n14224 & ~n14276_1;
  assign n14295 = ~n14224 & n14276_1;
  assign n14296_1 = ~n14294 & ~n14295;
  assign n14297 = ~n14231_1 & ~n14236_1;
  assign n14298 = ~n14237 & ~n14297;
  assign n14299 = ~n14296_1 & n14298;
  assign n14300 = n14224 & n14276_1;
  assign n14301_1 = ~n14224 & ~n14276_1;
  assign n14302 = ~n14300 & ~n14301_1;
  assign n14303 = ~n14298 & ~n14302;
  assign n14304 = ~n14299 & ~n14303;
  assign n14305 = n13711_1 & ~n14304;
  assign n14306_1 = ~n14277 & ~n14281_1;
  assign n14307 = ~n14293 & n14306_1;
  assign n14308 = ~n14305 & n14307;
  assign n14309 = ~n14148 & n14165;
  assign n14310 = n14208 & ~n14309;
  assign n14311_1 = n14148 & ~n14165;
  assign n14312 = ~n14310 & ~n14311_1;
  assign n14313 = ~n14147 & ~n14232;
  assign n14314 = ~n14180 & n14313;
  assign n14315 = n14312 & ~n14314;
  assign n14316_1 = n14296_1 & n14315;
  assign n14317 = ~n14296_1 & ~n14315;
  assign n14318 = ~n14316_1 & ~n14317;
  assign n14319 = n13733 & ~n14318;
  assign n14320 = n13781_1 & ~n14165;
  assign n14321_1 = n13727 & ~n14304;
  assign n14322 = n13730 & ~n14318;
  assign n14323 = ~n14321_1 & ~n14322;
  assign n14324 = n13722 & ~n14304;
  assign n14325 = n13717 & ~n14304;
  assign n14326_1 = n13719 & ~n14318;
  assign n14327 = n13725 & ~n14318;
  assign n14328 = ~n14326_1 & ~n14327;
  assign n14329 = ~n14324 & ~n14325;
  assign n14330 = n14328 & n14329;
  assign n14331_1 = ~n14319 & ~n14320;
  assign n14332 = n14323 & n14331_1;
  assign n14333 = n14330 & n14332;
  assign n14334 = n14308 & n14333;
  assign n14335 = n13658 & ~n14334;
  assign n14336_1 = P3_REG0_REG_9_ & ~n13658;
  assign n1166 = n14335 | n14336_1;
  assign n14338 = P3_REG1_REG_11_ & n13691_1;
  assign n14339 = P3_REG0_REG_11_ & n13689;
  assign n14340 = P3_REG2_REG_11_ & n13693;
  assign n14341_1 = P3_REG3_REG_10_ & n14285;
  assign n14342 = ~P3_REG3_REG_11_ & n14341_1;
  assign n14343 = P3_REG3_REG_11_ & ~n14341_1;
  assign n14344 = ~n14342 & ~n14343;
  assign n14345 = n13687 & ~n14344;
  assign n14346_1 = ~n14338 & ~n14339;
  assign n14347 = ~n14340 & n14346_1;
  assign n14348 = ~n14345 & n14347;
  assign n14349 = n13680 & ~n14348;
  assign n14350 = P3_IR_REG_31_ & n13204;
  assign n14351_1 = P3_IR_REG_10_ & ~P3_IR_REG_31_;
  assign n14352 = ~n14350 & ~n14351_1;
  assign n14353 = n13665 & ~n14352;
  assign n14354 = P1_P3_DATAO_REG_10_ & ~n13665;
  assign n14355 = ~n14353 & ~n14354;
  assign n14356_1 = ~n14292 & ~n14355;
  assign n14357 = n14292 & n14355;
  assign n14358 = ~n14300 & ~n14357;
  assign n14359 = ~n14356_1 & n14358;
  assign n14360 = n14298 & ~n14301_1;
  assign n14361_1 = n14359 & ~n14360;
  assign n14362 = n14292 & ~n14355;
  assign n14363 = ~n14292 & n14355;
  assign n14364 = ~n14362 & ~n14363;
  assign n14365 = ~n14301_1 & n14364;
  assign n14366_1 = ~n14298 & ~n14300;
  assign n14367 = n14365 & ~n14366_1;
  assign n14368 = ~n14361_1 & ~n14367;
  assign n14369 = n13711_1 & n14368;
  assign n14370 = ~n13677 & ~n14355;
  assign n14371_1 = n14278 & n14355;
  assign n14372 = ~n14278 & ~n14355;
  assign n14373 = ~n14371_1 & ~n14372;
  assign n14374 = n13699 & n14373;
  assign n14375 = ~n14349 & ~n14369;
  assign n14376_1 = ~n14370 & n14375;
  assign n14377 = ~n14374 & n14376_1;
  assign n14378 = ~n14294 & ~n14315;
  assign n14379 = ~n14295 & ~n14378;
  assign n14380 = n14364 & n14379;
  assign n14381_1 = ~n14364 & ~n14379;
  assign n14382 = ~n14380 & ~n14381_1;
  assign n14383 = n13733 & ~n14382;
  assign n14384 = n13781_1 & ~n14224;
  assign n14385 = n13727 & n14368;
  assign n14386_1 = n13730 & ~n14382;
  assign n14387 = ~n14385 & ~n14386_1;
  assign n14388 = n13722 & n14368;
  assign n14389 = n13717 & n14368;
  assign n14390 = n13719 & ~n14382;
  assign n14391_1 = n13725 & ~n14382;
  assign n14392 = ~n14390 & ~n14391_1;
  assign n14393 = ~n14388 & ~n14389;
  assign n14394 = n14392 & n14393;
  assign n14395 = ~n14383 & ~n14384;
  assign n14396_1 = n14387 & n14395;
  assign n14397 = n14394 & n14396_1;
  assign n14398 = n14377 & n14397;
  assign n14399 = n13658 & ~n14398;
  assign n14400 = P3_REG0_REG_10_ & ~n13658;
  assign n1171 = n14399 | n14400;
  assign n14402 = P3_IR_REG_31_ & n13212;
  assign n14403 = P3_IR_REG_11_ & ~P3_IR_REG_31_;
  assign n14404 = ~n14402 & ~n14403;
  assign n14405 = n13665 & ~n14404;
  assign n14406_1 = P1_P3_DATAO_REG_11_ & ~n13665;
  assign n14407 = ~n14405 & ~n14406_1;
  assign n14408 = ~n14348 & n14407;
  assign n14409 = n14348 & ~n14407;
  assign n14410 = ~n14408 & ~n14409;
  assign n14411_1 = ~n14362 & ~n14410;
  assign n14412 = ~n14363 & n14379;
  assign n14413 = n14411_1 & ~n14412;
  assign n14414 = ~n14363 & ~n14408;
  assign n14415 = ~n14409 & n14414;
  assign n14416_1 = ~n14362 & ~n14379;
  assign n14417 = n14415 & ~n14416_1;
  assign n14418 = ~n14413 & ~n14417;
  assign n14419 = n13733 & ~n14418;
  assign n14420 = n13781_1 & ~n14292;
  assign n14421_1 = ~n14301_1 & ~n14356_1;
  assign n14422 = n14237 & n14358;
  assign n14423 = n14421_1 & ~n14422;
  assign n14424 = ~n14357 & ~n14423;
  assign n14425 = ~n14236_1 & n14358;
  assign n14426_1 = ~n14231_1 & n14425;
  assign n14427 = ~n14424 & ~n14426_1;
  assign n14428 = ~n14410 & n14427;
  assign n14429 = n14348 & n14407;
  assign n14430 = ~n14348 & ~n14407;
  assign n14431_1 = ~n14429 & ~n14430;
  assign n14432 = ~n14427 & ~n14431_1;
  assign n14433 = ~n14428 & ~n14432;
  assign n14434 = n13727 & ~n14433;
  assign n14435 = n13730 & ~n14418;
  assign n14436_1 = ~n14434 & ~n14435;
  assign n14437 = n13722 & ~n14433;
  assign n14438 = n13717 & ~n14433;
  assign n14439 = n13719 & ~n14418;
  assign n14440 = n13725 & ~n14418;
  assign n14441_1 = ~n14439 & ~n14440;
  assign n14442 = ~n14437 & ~n14438;
  assign n14443 = n14441_1 & n14442;
  assign n14444 = ~n14419 & ~n14420;
  assign n14445 = n14436_1 & n14444;
  assign n14446_1 = n14443 & n14445;
  assign n14447 = ~n13677 & ~n14407;
  assign n14448 = P3_REG1_REG_12_ & n13691_1;
  assign n14449 = P3_REG0_REG_12_ & n13689;
  assign n14450 = P3_REG2_REG_12_ & n13693;
  assign n14451_1 = P3_REG3_REG_11_ & n14341_1;
  assign n14452 = ~P3_REG3_REG_12_ & n14451_1;
  assign n14453 = P3_REG3_REG_12_ & ~n14451_1;
  assign n14454 = ~n14452 & ~n14453;
  assign n14455 = n13687 & ~n14454;
  assign n14456_1 = ~n14448 & ~n14449;
  assign n14457 = ~n14450 & n14456_1;
  assign n14458 = ~n14455 & n14457;
  assign n14459 = n13680 & ~n14458;
  assign n14460 = n13711_1 & ~n14433;
  assign n14461_1 = n14371_1 & n14407;
  assign n14462 = ~n14371_1 & ~n14407;
  assign n14463 = ~n14461_1 & ~n14462;
  assign n14464 = n13699 & n14463;
  assign n14465 = ~n14459 & ~n14460;
  assign n14466_1 = ~n14464 & n14465;
  assign n14467 = n14446_1 & ~n14447;
  assign n14468 = n14466_1 & n14467;
  assign n14469 = n13658 & ~n14468;
  assign n14470 = P3_REG0_REG_11_ & ~n13658;
  assign n1176 = n14469 | n14470;
  assign n14472 = P3_IR_REG_31_ & n13223;
  assign n14473 = P3_IR_REG_12_ & ~P3_IR_REG_31_;
  assign n14474 = ~n14472 & ~n14473;
  assign n14475 = n13665 & ~n14474;
  assign n14476_1 = P1_P3_DATAO_REG_12_ & ~n13665;
  assign n14477 = ~n14475 & ~n14476_1;
  assign n14478 = ~n14458 & n14477;
  assign n14479 = n14458 & ~n14477;
  assign n14480 = ~n14478 & ~n14479;
  assign n14481_1 = ~n14362 & ~n14409;
  assign n14482 = n14295 & n14481_1;
  assign n14483 = n14414 & ~n14482;
  assign n14484 = ~n14409 & ~n14483;
  assign n14485 = n14378 & n14481_1;
  assign n14486_1 = ~n14484 & ~n14485;
  assign n14487 = ~n14480 & ~n14486_1;
  assign n14488 = n14480 & n14486_1;
  assign n14489 = ~n14487 & ~n14488;
  assign n14490 = n13733 & ~n14489;
  assign n14491_1 = n13781_1 & ~n14348;
  assign n14492 = ~n14427 & ~n14429;
  assign n14493 = ~n14430 & ~n14492;
  assign n14494 = ~n14480 & n14493;
  assign n14495 = n14458 & n14477;
  assign n14496_1 = ~n14458 & ~n14477;
  assign n14497 = ~n14495 & ~n14496_1;
  assign n14498 = ~n14493 & ~n14497;
  assign n14499 = ~n14494 & ~n14498;
  assign n14500 = n13727 & ~n14499;
  assign n14501_1 = n13730 & ~n14489;
  assign n14502 = ~n14500 & ~n14501_1;
  assign n14503 = n13722 & ~n14499;
  assign n14504 = n13717 & ~n14499;
  assign n14505 = n13719 & ~n14489;
  assign n14506_1 = n13725 & ~n14489;
  assign n14507 = ~n14505 & ~n14506_1;
  assign n14508 = ~n14503 & ~n14504;
  assign n14509 = n14507 & n14508;
  assign n14510 = ~n14490 & ~n14491_1;
  assign n14511_1 = n14502 & n14510;
  assign n14512 = n14509 & n14511_1;
  assign n14513 = ~n13677 & ~n14477;
  assign n14514 = P3_REG1_REG_13_ & n13691_1;
  assign n14515 = P3_REG0_REG_13_ & n13689;
  assign n14516_1 = P3_REG2_REG_13_ & n13693;
  assign n14517 = P3_REG3_REG_12_ & n14451_1;
  assign n14518 = ~P3_REG3_REG_13_ & n14517;
  assign n14519 = P3_REG3_REG_13_ & ~n14517;
  assign n14520 = ~n14518 & ~n14519;
  assign n14521_1 = n13687 & ~n14520;
  assign n14522 = ~n14514 & ~n14515;
  assign n14523 = ~n14516_1 & n14522;
  assign n14524 = ~n14521_1 & n14523;
  assign n14525 = n13680 & ~n14524;
  assign n14526_1 = n13711_1 & ~n14499;
  assign n14527 = n14461_1 & n14477;
  assign n14528 = ~n14461_1 & ~n14477;
  assign n14529 = ~n14527 & ~n14528;
  assign n14530 = n13699 & n14529;
  assign n14531_1 = ~n14525 & ~n14526_1;
  assign n14532 = ~n14530 & n14531_1;
  assign n14533 = n14512 & ~n14513;
  assign n14534 = n14532 & n14533;
  assign n14535 = n13658 & ~n14534;
  assign n14536_1 = P3_REG0_REG_12_ & ~n13658;
  assign n1181 = n14535 | n14536_1;
  assign n14538 = P3_IR_REG_31_ & n13231_1;
  assign n14539 = P3_IR_REG_13_ & ~P3_IR_REG_31_;
  assign n14540 = ~n14538 & ~n14539;
  assign n14541_1 = n13665 & ~n14540;
  assign n14542 = P1_P3_DATAO_REG_13_ & ~n13665;
  assign n14543 = ~n14541_1 & ~n14542;
  assign n14544 = ~n14524 & n14543;
  assign n14545 = n14524 & ~n14543;
  assign n14546_1 = ~n14544 & ~n14545;
  assign n14547 = ~n14479 & ~n14486_1;
  assign n14548 = ~n14478 & ~n14547;
  assign n14549 = ~n14546_1 & ~n14548;
  assign n14550 = n14546_1 & n14548;
  assign n14551_1 = ~n14549 & ~n14550;
  assign n14552 = n13733 & ~n14551_1;
  assign n14553 = n13781_1 & ~n14458;
  assign n14554 = ~n14524 & ~n14543;
  assign n14555 = n14524 & n14543;
  assign n14556_1 = ~n14495 & ~n14555;
  assign n14557 = ~n14554 & n14556_1;
  assign n14558 = n14493 & ~n14496_1;
  assign n14559 = n14557 & ~n14558;
  assign n14560 = ~n14496_1 & n14546_1;
  assign n14561_1 = ~n14493 & ~n14495;
  assign n14562 = n14560 & ~n14561_1;
  assign n14563 = ~n14559 & ~n14562;
  assign n14564 = n13727 & n14563;
  assign n14565 = n13730 & ~n14551_1;
  assign n14566_1 = ~n14564 & ~n14565;
  assign n14567 = n13722 & n14563;
  assign n14568 = n13717 & n14563;
  assign n14569 = n13719 & ~n14551_1;
  assign n14570 = n13725 & ~n14551_1;
  assign n14571_1 = ~n14569 & ~n14570;
  assign n14572 = ~n14567 & ~n14568;
  assign n14573 = n14571_1 & n14572;
  assign n14574 = ~n14552 & ~n14553;
  assign n14575 = n14566_1 & n14574;
  assign n14576_1 = n14573 & n14575;
  assign n14577 = ~n13677 & ~n14543;
  assign n14578 = P3_REG1_REG_14_ & n13691_1;
  assign n14579 = P3_REG0_REG_14_ & n13689;
  assign n14580 = P3_REG2_REG_14_ & n13693;
  assign n14581_1 = P3_REG3_REG_13_ & n14517;
  assign n14582 = ~P3_REG3_REG_14_ & n14581_1;
  assign n14583 = P3_REG3_REG_14_ & ~n14581_1;
  assign n14584 = ~n14582 & ~n14583;
  assign n14585 = n13687 & ~n14584;
  assign n14586_1 = ~n14578 & ~n14579;
  assign n14587 = ~n14580 & n14586_1;
  assign n14588 = ~n14585 & n14587;
  assign n14589 = n13680 & ~n14588;
  assign n14590 = n13711_1 & n14563;
  assign n14591_1 = n14527 & n14543;
  assign n14592 = ~n14527 & ~n14543;
  assign n14593 = ~n14591_1 & ~n14592;
  assign n14594 = n13699 & n14593;
  assign n14595 = ~n14589 & ~n14590;
  assign n14596_1 = ~n14594 & n14595;
  assign n14597 = n14576_1 & ~n14577;
  assign n14598 = n14596_1 & n14597;
  assign n14599 = n13658 & ~n14598;
  assign n14600 = P3_REG0_REG_13_ & ~n13658;
  assign n1186 = n14599 | n14600;
  assign n14602 = ~n14545 & ~n14548;
  assign n14603 = ~n14544 & ~n14602;
  assign n14604 = P3_IR_REG_31_ & n13240;
  assign n14605 = P3_IR_REG_14_ & ~P3_IR_REG_31_;
  assign n14606_1 = ~n14604 & ~n14605;
  assign n14607 = n13665 & ~n14606_1;
  assign n14608 = P1_P3_DATAO_REG_14_ & ~n13665;
  assign n14609 = ~n14607 & ~n14608;
  assign n14610 = ~n14588 & n14609;
  assign n14611_1 = n14588 & ~n14609;
  assign n14612 = ~n14610 & ~n14611_1;
  assign n14613 = n14603 & n14612;
  assign n14614 = ~n14603 & ~n14612;
  assign n14615 = ~n14613 & ~n14614;
  assign n14616_1 = n13733 & ~n14615;
  assign n14617 = n13781_1 & ~n14524;
  assign n14618 = ~n14496_1 & ~n14554;
  assign n14619 = n14430 & n14556_1;
  assign n14620 = n14618 & ~n14619;
  assign n14621_1 = ~n14555 & ~n14620;
  assign n14622 = n14492 & n14556_1;
  assign n14623 = ~n14621_1 & ~n14622;
  assign n14624 = ~n14612 & n14623;
  assign n14625 = n14612 & ~n14623;
  assign n14626_1 = ~n14624 & ~n14625;
  assign n14627 = n13727 & ~n14626_1;
  assign n14628 = n13730 & ~n14615;
  assign n14629 = ~n14627 & ~n14628;
  assign n14630 = n13722 & ~n14626_1;
  assign n14631_1 = n13717 & ~n14626_1;
  assign n14632 = n13719 & ~n14615;
  assign n14633 = n13725 & ~n14615;
  assign n14634 = ~n14632 & ~n14633;
  assign n14635 = ~n14630 & ~n14631_1;
  assign n14636_1 = n14634 & n14635;
  assign n14637 = ~n14616_1 & ~n14617;
  assign n14638 = n14629 & n14637;
  assign n14639 = n14636_1 & n14638;
  assign n14640 = ~n13677 & ~n14609;
  assign n14641_1 = P3_REG1_REG_15_ & n13691_1;
  assign n14642 = P3_REG0_REG_15_ & n13689;
  assign n14643 = P3_REG2_REG_15_ & n13693;
  assign n14644 = P3_REG3_REG_14_ & n14581_1;
  assign n14645 = ~P3_REG3_REG_15_ & n14644;
  assign n14646_1 = P3_REG3_REG_15_ & ~n14644;
  assign n14647 = ~n14645 & ~n14646_1;
  assign n14648 = n13687 & ~n14647;
  assign n14649 = ~n14641_1 & ~n14642;
  assign n14650 = ~n14643 & n14649;
  assign n14651_1 = ~n14648 & n14650;
  assign n14652 = n13680 & ~n14651_1;
  assign n14653 = n13711_1 & ~n14626_1;
  assign n14654 = n14591_1 & n14609;
  assign n14655 = ~n14591_1 & ~n14609;
  assign n14656_1 = ~n14654 & ~n14655;
  assign n14657 = n13699 & n14656_1;
  assign n14658 = ~n14652 & ~n14653;
  assign n14659 = ~n14657 & n14658;
  assign n14660 = n14639 & ~n14640;
  assign n14661_1 = n14659 & n14660;
  assign n14662 = n13658 & ~n14661_1;
  assign n14663 = P3_REG0_REG_14_ & ~n13658;
  assign n1191 = n14662 | n14663;
  assign n14665 = P3_IR_REG_31_ & n13248;
  assign n14666_1 = P3_IR_REG_15_ & ~P3_IR_REG_31_;
  assign n14667 = ~n14665 & ~n14666_1;
  assign n14668 = n13665 & ~n14667;
  assign n14669 = P1_P3_DATAO_REG_15_ & ~n13665;
  assign n14670 = ~n14668 & ~n14669;
  assign n14671_1 = ~n14651_1 & n14670;
  assign n14672 = n14651_1 & ~n14670;
  assign n14673 = ~n14671_1 & ~n14672;
  assign n14674 = ~n14603 & ~n14611_1;
  assign n14675 = ~n14610 & ~n14674;
  assign n14676_1 = n14673 & n14675;
  assign n14677 = ~n14673 & ~n14675;
  assign n14678 = ~n14676_1 & ~n14677;
  assign n14679 = n13733 & ~n14678;
  assign n14680 = n13781_1 & ~n14588;
  assign n14681_1 = ~n14588 & ~n14609;
  assign n14682 = n14588 & n14609;
  assign n14683 = ~n14623 & ~n14682;
  assign n14684 = ~n14681_1 & ~n14683;
  assign n14685 = ~n14673 & n14684;
  assign n14686_1 = n14673 & ~n14684;
  assign n14687 = ~n14685 & ~n14686_1;
  assign n14688 = n13727 & ~n14687;
  assign n14689 = n13730 & ~n14678;
  assign n14690 = ~n14688 & ~n14689;
  assign n14691_1 = n13722 & ~n14687;
  assign n14692 = n13717 & ~n14687;
  assign n14693 = n13719 & ~n14678;
  assign n14694 = n13725 & ~n14678;
  assign n14695 = ~n14693 & ~n14694;
  assign n14696_1 = ~n14691_1 & ~n14692;
  assign n14697 = n14695 & n14696_1;
  assign n14698 = ~n14679 & ~n14680;
  assign n14699 = n14690 & n14698;
  assign n14700 = n14697 & n14699;
  assign n14701_1 = ~n13677 & ~n14670;
  assign n14702 = P3_REG1_REG_16_ & n13691_1;
  assign n14703 = P3_REG0_REG_16_ & n13689;
  assign n14704 = P3_REG2_REG_16_ & n13693;
  assign n14705 = P3_REG3_REG_15_ & n14644;
  assign n14706_1 = ~P3_REG3_REG_16_ & n14705;
  assign n14707 = P3_REG3_REG_16_ & ~n14705;
  assign n14708 = ~n14706_1 & ~n14707;
  assign n14709 = n13687 & ~n14708;
  assign n14710 = ~n14702 & ~n14703;
  assign n14711_1 = ~n14704 & n14710;
  assign n14712 = ~n14709 & n14711_1;
  assign n14713 = n13680 & ~n14712;
  assign n14714 = n13711_1 & ~n14687;
  assign n14715 = n14654 & n14670;
  assign n14716_1 = ~n14654 & ~n14670;
  assign n14717 = ~n14715 & ~n14716_1;
  assign n14718 = n13699 & n14717;
  assign n14719 = ~n14713 & ~n14714;
  assign n14720 = ~n14718 & n14719;
  assign n14721_1 = n14700 & ~n14701_1;
  assign n14722 = n14720 & n14721_1;
  assign n14723 = n13658 & ~n14722;
  assign n14724 = P3_REG0_REG_15_ & ~n13658;
  assign n1196 = n14723 | n14724;
  assign n14726_1 = P3_IR_REG_31_ & n13270;
  assign n14727 = P3_IR_REG_16_ & ~P3_IR_REG_31_;
  assign n14728 = ~n14726_1 & ~n14727;
  assign n14729 = n13665 & ~n14728;
  assign n14730 = P1_P3_DATAO_REG_16_ & ~n13665;
  assign n14731_1 = ~n14729 & ~n14730;
  assign n14732 = ~n14712 & n14731_1;
  assign n14733 = n14712 & ~n14731_1;
  assign n14734 = ~n14732 & ~n14733;
  assign n14735 = ~n14672 & ~n14734;
  assign n14736_1 = ~n14671_1 & n14675;
  assign n14737 = n14735 & ~n14736_1;
  assign n14738 = ~n14672 & ~n14675;
  assign n14739 = ~n14671_1 & ~n14732;
  assign n14740 = ~n14733 & ~n14738;
  assign n14741_1 = n14739 & n14740;
  assign n14742 = ~n14737 & ~n14741_1;
  assign n14743 = n13733 & ~n14742;
  assign n14744 = n13781_1 & ~n14651_1;
  assign n14745 = ~n14651_1 & ~n14670;
  assign n14746_1 = n14651_1 & n14670;
  assign n14747 = ~n14684 & ~n14746_1;
  assign n14748 = ~n14745 & ~n14747;
  assign n14749 = ~n14734 & n14748;
  assign n14750 = n14712 & n14731_1;
  assign n14751_1 = ~n14712 & ~n14731_1;
  assign n14752 = ~n14750 & ~n14751_1;
  assign n14753 = ~n14748 & ~n14752;
  assign n14754 = ~n14749 & ~n14753;
  assign n14755 = n13727 & ~n14754;
  assign n14756_1 = n13730 & ~n14742;
  assign n14757 = ~n14755 & ~n14756_1;
  assign n14758 = n13722 & ~n14754;
  assign n14759 = n13717 & ~n14754;
  assign n14760 = n13719 & ~n14742;
  assign n14761_1 = n13725 & ~n14742;
  assign n14762 = ~n14760 & ~n14761_1;
  assign n14763 = ~n14758 & ~n14759;
  assign n14764 = n14762 & n14763;
  assign n14765 = ~n14743 & ~n14744;
  assign n14766_1 = n14757 & n14765;
  assign n14767 = n14764 & n14766_1;
  assign n14768 = ~n13677 & ~n14731_1;
  assign n14769 = P3_REG1_REG_17_ & n13691_1;
  assign n14770 = P3_REG0_REG_17_ & n13689;
  assign n14771_1 = P3_REG2_REG_17_ & n13693;
  assign n14772 = P3_REG3_REG_16_ & n14705;
  assign n14773 = ~P3_REG3_REG_17_ & n14772;
  assign n14774 = P3_REG3_REG_17_ & ~n14772;
  assign n14775 = ~n14773 & ~n14774;
  assign n14776_1 = n13687 & ~n14775;
  assign n14777 = ~n14769 & ~n14770;
  assign n14778 = ~n14771_1 & n14777;
  assign n14779 = ~n14776_1 & n14778;
  assign n14780 = n13680 & ~n14779;
  assign n14781_1 = n13711_1 & ~n14754;
  assign n14782 = n14715 & n14731_1;
  assign n14783 = ~n14715 & ~n14731_1;
  assign n14784 = ~n14782 & ~n14783;
  assign n14785 = n13699 & n14784;
  assign n14786_1 = ~n14780 & ~n14781_1;
  assign n14787 = ~n14785 & n14786_1;
  assign n14788 = n14767 & ~n14768;
  assign n14789 = n14787 & n14788;
  assign n14790 = n13658 & ~n14789;
  assign n14791_1 = P3_REG0_REG_16_ & ~n13658;
  assign n1201 = n14790 | n14791_1;
  assign n14793 = P3_IR_REG_31_ & n13278;
  assign n14794 = P3_IR_REG_17_ & ~P3_IR_REG_31_;
  assign n14795 = ~n14793 & ~n14794;
  assign n14796_1 = n13665 & ~n14795;
  assign n14797 = P1_P3_DATAO_REG_17_ & ~n13665;
  assign n14798 = ~n14796_1 & ~n14797;
  assign n14799 = ~n14779 & n14798;
  assign n14800 = n14779 & ~n14798;
  assign n14801_1 = ~n14799 & ~n14800;
  assign n14802 = n14610 & ~n14672;
  assign n14803 = n14739 & ~n14802;
  assign n14804 = ~n14733 & ~n14803;
  assign n14805 = ~n14672 & n14674;
  assign n14806_1 = ~n14733 & n14805;
  assign n14807 = ~n14804 & ~n14806_1;
  assign n14808 = ~n14801_1 & ~n14807;
  assign n14809 = n14801_1 & n14807;
  assign n14810 = ~n14808 & ~n14809;
  assign n14811_1 = n13733 & ~n14810;
  assign n14812 = n13781_1 & ~n14712;
  assign n14813 = ~n14779 & ~n14798;
  assign n14814 = n14748 & ~n14751_1;
  assign n14815 = n14779 & n14798;
  assign n14816_1 = ~n14750 & ~n14815;
  assign n14817 = ~n14813 & ~n14814;
  assign n14818 = n14816_1 & n14817;
  assign n14819 = ~n14751_1 & n14801_1;
  assign n14820 = ~n14748 & ~n14750;
  assign n14821_1 = n14819 & ~n14820;
  assign n14822 = ~n14818 & ~n14821_1;
  assign n14823 = n13727 & n14822;
  assign n14824 = n13730 & ~n14810;
  assign n14825 = ~n14823 & ~n14824;
  assign n14826_1 = n13722 & n14822;
  assign n14827 = n13717 & n14822;
  assign n14828 = n13719 & ~n14810;
  assign n14829 = n13725 & ~n14810;
  assign n14830 = ~n14828 & ~n14829;
  assign n14831_1 = ~n14826_1 & ~n14827;
  assign n14832 = n14830 & n14831_1;
  assign n14833 = ~n14811_1 & ~n14812;
  assign n14834 = n14825 & n14833;
  assign n14835 = n14832 & n14834;
  assign n14836_1 = P3_REG1_REG_18_ & n13691_1;
  assign n14837 = P3_REG0_REG_18_ & n13689;
  assign n14838 = P3_REG2_REG_18_ & n13693;
  assign n14839 = P3_REG3_REG_17_ & n14772;
  assign n14840 = ~P3_REG3_REG_18_ & n14839;
  assign n14841_1 = P3_REG3_REG_18_ & ~n14839;
  assign n14842 = ~n14840 & ~n14841_1;
  assign n14843 = n13687 & ~n14842;
  assign n14844 = ~n14836_1 & ~n14837;
  assign n14845 = ~n14838 & n14844;
  assign n14846_1 = ~n14843 & n14845;
  assign n14847 = n13680 & ~n14846_1;
  assign n14848 = n13711_1 & n14822;
  assign n14849 = ~n13677 & ~n14798;
  assign n14850 = ~n14847 & ~n14848;
  assign n14851_1 = ~n14849 & n14850;
  assign n14852 = n14782 & n14798;
  assign n14853 = ~n14782 & ~n14798;
  assign n14854 = ~n14852 & ~n14853;
  assign n14855 = n13699 & n14854;
  assign n14856_1 = n14835 & n14851_1;
  assign n14857 = ~n14855 & n14856_1;
  assign n14858 = n13658 & ~n14857;
  assign n14859 = P3_REG0_REG_17_ & ~n13658;
  assign n1206 = n14858 | n14859;
  assign n14861_1 = P3_IR_REG_31_ & n13296_1;
  assign n14862 = P3_IR_REG_18_ & ~P3_IR_REG_31_;
  assign n14863 = ~n14861_1 & ~n14862;
  assign n14864 = n13665 & ~n14863;
  assign n14865 = P1_P3_DATAO_REG_18_ & ~n13665;
  assign n14866_1 = ~n14864 & ~n14865;
  assign n14867 = ~n14846_1 & n14866_1;
  assign n14868 = n14846_1 & ~n14866_1;
  assign n14869 = ~n14867 & ~n14868;
  assign n14870 = ~n14800 & ~n14807;
  assign n14871_1 = ~n14799 & ~n14870;
  assign n14872 = ~n14869 & ~n14871_1;
  assign n14873 = n14869 & n14871_1;
  assign n14874 = ~n14872 & ~n14873;
  assign n14875 = n13733 & ~n14874;
  assign n14876_1 = n13781_1 & ~n14779;
  assign n14877 = n14751_1 & ~n14798;
  assign n14878 = ~n14751_1 & n14798;
  assign n14879 = ~n14779 & ~n14878;
  assign n14880 = ~n14877 & ~n14879;
  assign n14881_1 = ~n14748 & n14816_1;
  assign n14882 = n14880 & ~n14881_1;
  assign n14883 = ~n14869 & n14882;
  assign n14884 = n14846_1 & n14866_1;
  assign n14885 = ~n14846_1 & ~n14866_1;
  assign n14886_1 = ~n14884 & ~n14885;
  assign n14887 = ~n14882 & ~n14886_1;
  assign n14888 = ~n14883 & ~n14887;
  assign n14889 = n13727 & ~n14888;
  assign n14890 = n13730 & ~n14874;
  assign n14891_1 = ~n14889 & ~n14890;
  assign n14892 = n13722 & ~n14888;
  assign n14893 = n13717 & ~n14888;
  assign n14894 = n13719 & ~n14874;
  assign n14895 = n13725 & ~n14874;
  assign n14896_1 = ~n14894 & ~n14895;
  assign n14897 = ~n14892 & ~n14893;
  assign n14898 = n14896_1 & n14897;
  assign n14899 = ~n14875 & ~n14876_1;
  assign n14900 = n14891_1 & n14899;
  assign n14901_1 = n14898 & n14900;
  assign n14902 = P3_REG1_REG_19_ & n13691_1;
  assign n14903 = P3_REG0_REG_19_ & n13689;
  assign n14904 = P3_REG2_REG_19_ & n13693;
  assign n14905 = P3_REG3_REG_18_ & n14839;
  assign n14906_1 = ~P3_REG3_REG_19_ & n14905;
  assign n14907 = P3_REG3_REG_19_ & ~n14905;
  assign n14908 = ~n14906_1 & ~n14907;
  assign n14909 = n13687 & ~n14908;
  assign n14910 = ~n14902 & ~n14903;
  assign n14911_1 = ~n14904 & n14910;
  assign n14912 = ~n14909 & n14911_1;
  assign n14913 = n13680 & ~n14912;
  assign n14914 = n13711_1 & ~n14888;
  assign n14915 = ~n13677 & ~n14866_1;
  assign n14916_1 = ~n14913 & ~n14914;
  assign n14917 = ~n14915 & n14916_1;
  assign n14918 = n14852 & n14866_1;
  assign n14919 = ~n14852 & ~n14866_1;
  assign n14920 = ~n14918 & ~n14919;
  assign n14921_1 = n13699 & n14920;
  assign n14922 = n14901_1 & n14917;
  assign n14923 = ~n14921_1 & n14922;
  assign n14924 = n13658 & ~n14923;
  assign n14925 = P3_REG0_REG_18_ & ~n13658;
  assign n1211 = n14924 | n14925;
  assign n14927 = ~n13593 & n13665;
  assign n14928 = P1_P3_DATAO_REG_19_ & ~n13665;
  assign n14929 = ~n14927 & ~n14928;
  assign n14930 = ~n14912 & n14929;
  assign n14931_1 = n14912 & ~n14929;
  assign n14932 = ~n14930 & ~n14931_1;
  assign n14933 = ~n14846_1 & ~n14871_1;
  assign n14934 = n14846_1 & n14871_1;
  assign n14935 = n14866_1 & ~n14934;
  assign n14936_1 = ~n14933 & ~n14935;
  assign n14937 = ~n14932 & ~n14936_1;
  assign n14938 = n14932 & n14936_1;
  assign n14939 = ~n14937 & ~n14938;
  assign n14940 = n13733 & ~n14939;
  assign n14941_1 = n13781_1 & ~n14846_1;
  assign n14942 = ~n14882 & ~n14884;
  assign n14943 = ~n14885 & ~n14942;
  assign n14944 = ~n14932 & n14943;
  assign n14945 = n14912 & n14929;
  assign n14946_1 = ~n14912 & ~n14929;
  assign n14947 = ~n14945 & ~n14946_1;
  assign n14948 = ~n14943 & ~n14947;
  assign n14949 = ~n14944 & ~n14948;
  assign n14950 = n13727 & ~n14949;
  assign n14951_1 = n13730 & ~n14939;
  assign n14952 = ~n14950 & ~n14951_1;
  assign n14953 = n13722 & ~n14949;
  assign n14954 = n13717 & ~n14949;
  assign n14955 = n13719 & ~n14939;
  assign n14956_1 = n13725 & ~n14939;
  assign n14957 = ~n14955 & ~n14956_1;
  assign n14958 = ~n14953 & ~n14954;
  assign n14959 = n14957 & n14958;
  assign n14960 = ~n14940 & ~n14941_1;
  assign n14961_1 = n14952 & n14960;
  assign n14962 = n14959 & n14961_1;
  assign n14963 = ~n13677 & ~n14929;
  assign n14964 = P3_REG1_REG_20_ & n13691_1;
  assign n14965 = P3_REG0_REG_20_ & n13689;
  assign n14966_1 = P3_REG2_REG_20_ & n13693;
  assign n14967 = P3_REG3_REG_19_ & n14905;
  assign n14968 = ~P3_REG3_REG_20_ & n14967;
  assign n14969 = P3_REG3_REG_20_ & ~n14967;
  assign n14970 = ~n14968 & ~n14969;
  assign n14971_1 = n13687 & ~n14970;
  assign n14972 = ~n14964 & ~n14965;
  assign n14973 = ~n14966_1 & n14972;
  assign n14974 = ~n14971_1 & n14973;
  assign n14975 = n13680 & ~n14974;
  assign n14976_1 = n13711_1 & ~n14949;
  assign n14977 = n14918 & n14929;
  assign n14978 = ~n14918 & ~n14929;
  assign n14979 = ~n14977 & ~n14978;
  assign n14980 = n13699 & n14979;
  assign n14981_1 = ~n14975 & ~n14976_1;
  assign n14982 = ~n14980 & n14981_1;
  assign n14983 = n14962 & ~n14963;
  assign n14984 = n14982 & n14983;
  assign n14985 = n13658 & ~n14984;
  assign n14986_1 = P3_REG0_REG_19_ & ~n13658;
  assign n1216 = n14985 | n14986_1;
  assign n14988 = LOGIC0 & ~n13665;
  assign n14989 = ~n14974 & ~n14988;
  assign n14990 = n14974 & n14988;
  assign n14991_1 = ~n14989 & ~n14990;
  assign n14992 = ~n14931_1 & ~n14936_1;
  assign n14993 = ~n14930 & ~n14992;
  assign n14994 = ~n14991_1 & ~n14993;
  assign n14995 = n14991_1 & n14993;
  assign n14996_1 = ~n14994 & ~n14995;
  assign n14997 = n13733 & ~n14996_1;
  assign n14998 = n13781_1 & ~n14912;
  assign n14999 = ~n14974 & n14988;
  assign n15000 = n14943 & ~n14946_1;
  assign n15001_1 = n14974 & ~n14988;
  assign n15002 = ~n14945 & ~n15001_1;
  assign n15003 = ~n14999 & ~n15000;
  assign n15004 = n15002 & n15003;
  assign n15005 = ~n14943 & ~n14945;
  assign n15006_1 = ~n14946_1 & ~n15005;
  assign n15007 = n14991_1 & n15006_1;
  assign n15008 = ~n15004 & ~n15007;
  assign n15009 = n13727 & n15008;
  assign n15010 = n13730 & ~n14996_1;
  assign n15011_1 = ~n15009 & ~n15010;
  assign n15012 = n13722 & n15008;
  assign n15013 = n13717 & n15008;
  assign n15014 = n13719 & ~n14996_1;
  assign n15015 = n13725 & ~n14996_1;
  assign n15016_1 = ~n15014 & ~n15015;
  assign n15017 = ~n15012 & ~n15013;
  assign n15018 = n15016_1 & n15017;
  assign n15019 = ~n14997 & ~n14998;
  assign n15020 = n15011_1 & n15019;
  assign n15021_1 = n15018 & n15020;
  assign n15022 = ~n13677 & n14988;
  assign n15023 = P3_REG1_REG_21_ & n13691_1;
  assign n15024 = P3_REG0_REG_21_ & n13689;
  assign n15025 = P3_REG2_REG_21_ & n13693;
  assign n15026_1 = P3_REG3_REG_20_ & n14967;
  assign n15027 = ~P3_REG3_REG_21_ & n15026_1;
  assign n15028 = P3_REG3_REG_21_ & ~n15026_1;
  assign n15029 = ~n15027 & ~n15028;
  assign n15030 = n13687 & ~n15029;
  assign n15031_1 = ~n15023 & ~n15024;
  assign n15032 = ~n15025 & n15031_1;
  assign n15033 = ~n15030 & n15032;
  assign n15034 = n13680 & ~n15033;
  assign n15035 = n13711_1 & n15008;
  assign n15036_1 = n14977 & ~n14988;
  assign n15037 = ~n14977 & n14988;
  assign n15038 = ~n15036_1 & ~n15037;
  assign n15039 = n13699 & n15038;
  assign n15040 = ~n15034 & ~n15035;
  assign n15041_1 = ~n15039 & n15040;
  assign n15042 = n15021_1 & ~n15022;
  assign n15043 = n15041_1 & n15042;
  assign n15044 = n13658 & ~n15043;
  assign n15045 = P3_REG0_REG_20_ & ~n13658;
  assign n1221 = n15044 | n15045;
  assign n15047 = ~n14990 & ~n14993;
  assign n15048 = ~n14989 & ~n15047;
  assign n15049 = ~n14988 & ~n15033;
  assign n15050 = n14988 & n15033;
  assign n15051_1 = ~n15049 & ~n15050;
  assign n15052 = n15048 & n15051_1;
  assign n15053 = ~n15048 & ~n15051_1;
  assign n15054 = ~n15052 & ~n15053;
  assign n15055 = n13733 & ~n15054;
  assign n15056_1 = n13781_1 & ~n14974;
  assign n15057 = ~n14943 & n15002;
  assign n15058 = ~n14946_1 & ~n14988;
  assign n15059 = n14946_1 & n14988;
  assign n15060 = n14974 & ~n15059;
  assign n15061_1 = ~n15058 & ~n15060;
  assign n15062 = ~n15057 & ~n15061_1;
  assign n15063 = ~n15051_1 & ~n15062;
  assign n15064 = n15051_1 & ~n15061_1;
  assign n15065 = ~n15057 & n15064;
  assign n15066_1 = ~n15063 & ~n15065;
  assign n15067 = n13727 & n15066_1;
  assign n15068 = n13730 & ~n15054;
  assign n15069 = ~n15067 & ~n15068;
  assign n15070 = n13722 & n15066_1;
  assign n15071_1 = n13717 & n15066_1;
  assign n15072 = n13719 & ~n15054;
  assign n15073 = n13725 & ~n15054;
  assign n15074 = ~n15072 & ~n15073;
  assign n15075 = ~n15070 & ~n15071_1;
  assign n15076_1 = n15074 & n15075;
  assign n15077 = ~n15055 & ~n15056_1;
  assign n15078 = n15069 & n15077;
  assign n15079 = n15076_1 & n15078;
  assign n15080 = P3_REG1_REG_22_ & n13691_1;
  assign n15081_1 = P3_REG0_REG_22_ & n13689;
  assign n15082 = P3_REG2_REG_22_ & n13693;
  assign n15083 = P3_REG3_REG_21_ & n15026_1;
  assign n15084 = ~P3_REG3_REG_22_ & n15083;
  assign n15085 = P3_REG3_REG_22_ & ~n15083;
  assign n15086_1 = ~n15084 & ~n15085;
  assign n15087 = n13687 & ~n15086_1;
  assign n15088 = ~n15080 & ~n15081_1;
  assign n15089 = ~n15082 & n15088;
  assign n15090 = ~n15087 & n15089;
  assign n15091_1 = n13680 & ~n15090;
  assign n15092 = n13711_1 & n15066_1;
  assign n15093 = ~n14988 & n15036_1;
  assign n15094 = n14988 & ~n15036_1;
  assign n15095 = ~n15093 & ~n15094;
  assign n15096_1 = n13699 & n15095;
  assign n15097 = ~n15091_1 & ~n15092;
  assign n15098 = ~n15096_1 & n15097;
  assign n15099 = ~n15022 & n15079;
  assign n15100 = n15098 & n15099;
  assign n15101_1 = n13658 & ~n15100;
  assign n15102 = P3_REG0_REG_21_ & ~n13658;
  assign n1226 = n15101_1 | n15102;
  assign n15104 = ~n14988 & ~n15090;
  assign n15105 = n14988 & n15090;
  assign n15106_1 = ~n15104 & ~n15105;
  assign n15107 = ~n15048 & ~n15050;
  assign n15108 = ~n15049 & ~n15107;
  assign n15109 = n15106_1 & n15108;
  assign n15110 = ~n15106_1 & ~n15108;
  assign n15111_1 = ~n15109 & ~n15110;
  assign n15112 = n13733 & ~n15111_1;
  assign n15113 = n13781_1 & ~n15033;
  assign n15114 = ~n14988 & n15033;
  assign n15115 = n14885 & n15002;
  assign n15116_1 = ~n15061_1 & ~n15115;
  assign n15117 = ~n15114 & ~n15116_1;
  assign n15118 = n14988 & ~n15033;
  assign n15119 = ~n15117 & ~n15118;
  assign n15120 = ~n14884 & n15002;
  assign n15121_1 = ~n14882 & ~n15114;
  assign n15122 = n15120 & n15121_1;
  assign n15123 = n15119 & ~n15122;
  assign n15124 = ~n15106_1 & n15123;
  assign n15125 = n15106_1 & ~n15123;
  assign n15126_1 = ~n15124 & ~n15125;
  assign n15127 = n13727 & ~n15126_1;
  assign n15128 = n13730 & ~n15111_1;
  assign n15129 = ~n15127 & ~n15128;
  assign n15130 = n13722 & ~n15126_1;
  assign n15131_1 = n13717 & ~n15126_1;
  assign n15132 = n13719 & ~n15111_1;
  assign n15133 = n13725 & ~n15111_1;
  assign n15134 = ~n15132 & ~n15133;
  assign n15135 = ~n15130 & ~n15131_1;
  assign n15136_1 = n15134 & n15135;
  assign n15137 = ~n15112 & ~n15113;
  assign n15138 = n15129 & n15137;
  assign n15139 = n15136_1 & n15138;
  assign n15140 = P3_REG1_REG_23_ & n13691_1;
  assign n15141_1 = P3_REG0_REG_23_ & n13689;
  assign n15142 = P3_REG2_REG_23_ & n13693;
  assign n15143 = P3_REG3_REG_22_ & n15083;
  assign n15144 = ~P3_REG3_REG_23_ & n15143;
  assign n15145 = P3_REG3_REG_23_ & ~n15143;
  assign n15146_1 = ~n15144 & ~n15145;
  assign n15147 = n13687 & ~n15146_1;
  assign n15148 = ~n15140 & ~n15141_1;
  assign n15149 = ~n15142 & n15148;
  assign n15150 = ~n15147 & n15149;
  assign n15151_1 = n13680 & ~n15150;
  assign n15152 = n13711_1 & ~n15126_1;
  assign n15153 = ~n14988 & n15093;
  assign n15154 = n14988 & ~n15093;
  assign n15155 = ~n15153 & ~n15154;
  assign n15156_1 = n13699 & n15155;
  assign n15157 = ~n15151_1 & ~n15152;
  assign n15158 = ~n15156_1 & n15157;
  assign n15159 = ~n15022 & n15139;
  assign n15160 = n15158 & n15159;
  assign n15161_1 = n13658 & ~n15160;
  assign n15162 = P3_REG0_REG_22_ & ~n13658;
  assign n1231 = n15161_1 | n15162;
  assign n15164 = ~n14988 & ~n15150;
  assign n15165 = n14988 & n15150;
  assign n15166_1 = ~n15164 & ~n15165;
  assign n15167 = ~n15105 & ~n15166_1;
  assign n15168 = ~n15104 & n15108;
  assign n15169 = n15167 & ~n15168;
  assign n15170 = ~n15105 & ~n15108;
  assign n15171_1 = ~n15104 & ~n15164;
  assign n15172 = ~n15165 & ~n15170;
  assign n15173 = n15171_1 & n15172;
  assign n15174 = ~n15169 & ~n15173;
  assign n15175 = n13733 & ~n15174;
  assign n15176_1 = n13781_1 & ~n15090;
  assign n15177 = n14988 & ~n15090;
  assign n15178 = ~n14988 & n15090;
  assign n15179 = ~n15123 & ~n15178;
  assign n15180 = ~n15177 & ~n15179;
  assign n15181_1 = ~n15166_1 & n15180;
  assign n15182 = n15166_1 & ~n15180;
  assign n15183 = ~n15181_1 & ~n15182;
  assign n15184 = n13727 & ~n15183;
  assign n15185 = n13730 & ~n15174;
  assign n15186_1 = ~n15184 & ~n15185;
  assign n15187 = n13722 & ~n15183;
  assign n15188 = n13717 & ~n15183;
  assign n15189 = n13719 & ~n15174;
  assign n15190 = n13725 & ~n15174;
  assign n15191_1 = ~n15189 & ~n15190;
  assign n15192 = ~n15187 & ~n15188;
  assign n15193 = n15191_1 & n15192;
  assign n15194 = ~n15175 & ~n15176_1;
  assign n15195 = n15186_1 & n15194;
  assign n15196_1 = n15193 & n15195;
  assign n15197 = P3_REG1_REG_24_ & n13691_1;
  assign n15198 = P3_REG0_REG_24_ & n13689;
  assign n15199 = P3_REG2_REG_24_ & n13693;
  assign n15200 = P3_REG3_REG_23_ & n15143;
  assign n15201_1 = ~P3_REG3_REG_24_ & n15200;
  assign n15202 = P3_REG3_REG_24_ & ~n15200;
  assign n15203 = ~n15201_1 & ~n15202;
  assign n15204 = n13687 & ~n15203;
  assign n15205 = ~n15197 & ~n15198;
  assign n15206_1 = ~n15199 & n15205;
  assign n15207 = ~n15204 & n15206_1;
  assign n15208 = n13680 & ~n15207;
  assign n15209 = n13711_1 & ~n15183;
  assign n15210 = ~n14988 & n15153;
  assign n15211_1 = n14988 & ~n15153;
  assign n15212 = ~n15210 & ~n15211_1;
  assign n15213 = n13699 & n15212;
  assign n15214 = ~n15208 & ~n15209;
  assign n15215 = ~n15213 & n15214;
  assign n15216_1 = ~n15022 & n15196_1;
  assign n15217 = n15215 & n15216_1;
  assign n15218 = n13658 & ~n15217;
  assign n15219 = P3_REG0_REG_23_ & ~n13658;
  assign n1236 = n15218 | n15219;
  assign n15221_1 = ~n14988 & ~n15207;
  assign n15222 = n14988 & n15207;
  assign n15223 = ~n15221_1 & ~n15222;
  assign n15224 = n15049 & ~n15105;
  assign n15225 = n15171_1 & ~n15224;
  assign n15226_1 = ~n15165 & ~n15225;
  assign n15227 = ~n15050 & ~n15105;
  assign n15228 = ~n15048 & n15227;
  assign n15229 = ~n15165 & n15228;
  assign n15230 = ~n15226_1 & ~n15229;
  assign n15231_1 = ~n15223 & ~n15230;
  assign n15232 = n15223 & n15230;
  assign n15233 = ~n15231_1 & ~n15232;
  assign n15234 = n13733 & ~n15233;
  assign n15235 = n13781_1 & ~n15150;
  assign n15236_1 = n14988 & ~n15150;
  assign n15237 = ~n14988 & n15150;
  assign n15238 = ~n15180 & ~n15237;
  assign n15239 = ~n15236_1 & ~n15238;
  assign n15240 = ~n15223 & n15239;
  assign n15241_1 = ~n14988 & n15207;
  assign n15242 = n14988 & ~n15207;
  assign n15243 = ~n15241_1 & ~n15242;
  assign n15244 = ~n15239 & ~n15243;
  assign n15245 = ~n15240 & ~n15244;
  assign n15246_1 = n13727 & ~n15245;
  assign n15247 = n13730 & ~n15233;
  assign n15248 = ~n15246_1 & ~n15247;
  assign n15249 = n13722 & ~n15245;
  assign n15250 = n13717 & ~n15245;
  assign n15251_1 = n13719 & ~n15233;
  assign n15252 = n13725 & ~n15233;
  assign n15253 = ~n15251_1 & ~n15252;
  assign n15254 = ~n15249 & ~n15250;
  assign n15255 = n15253 & n15254;
  assign n15256_1 = ~n15234 & ~n15235;
  assign n15257 = n15248 & n15256_1;
  assign n15258 = n15255 & n15257;
  assign n15259 = P3_REG1_REG_25_ & n13691_1;
  assign n15260 = P3_REG0_REG_25_ & n13689;
  assign n15261_1 = P3_REG2_REG_25_ & n13693;
  assign n15262 = P3_REG3_REG_24_ & n15200;
  assign n15263 = ~P3_REG3_REG_25_ & n15262;
  assign n15264 = P3_REG3_REG_25_ & ~n15262;
  assign n15265 = ~n15263 & ~n15264;
  assign n15266_1 = n13687 & ~n15265;
  assign n15267 = ~n15259 & ~n15260;
  assign n15268 = ~n15261_1 & n15267;
  assign n15269 = ~n15266_1 & n15268;
  assign n15270 = n13680 & ~n15269;
  assign n15271_1 = n13711_1 & ~n15245;
  assign n15272 = ~n15270 & ~n15271_1;
  assign n15273 = ~n15022 & n15272;
  assign n15274 = ~n14988 & n15210;
  assign n15275 = n14988 & ~n15210;
  assign n15276_1 = ~n15274 & ~n15275;
  assign n15277 = n13699 & n15276_1;
  assign n15278 = n15258 & n15273;
  assign n15279 = ~n15277 & n15278;
  assign n15280 = n13658 & ~n15279;
  assign n15281_1 = P3_REG0_REG_24_ & ~n13658;
  assign n1241 = n15280 | n15281_1;
  assign n15283 = ~n14988 & ~n15269;
  assign n15284 = n14988 & n15269;
  assign n15285 = ~n15283 & ~n15284;
  assign n15286_1 = ~n15222 & ~n15230;
  assign n15287 = ~n15221_1 & ~n15286_1;
  assign n15288 = ~n15285 & ~n15287;
  assign n15289 = n15285 & n15287;
  assign n15290 = ~n15288 & ~n15289;
  assign n15291_1 = n13733 & ~n15290;
  assign n15292 = n13781_1 & ~n15207;
  assign n15293 = ~n15239 & ~n15241_1;
  assign n15294 = ~n15242 & ~n15293;
  assign n15295 = ~n15285 & n15294;
  assign n15296_1 = ~n14988 & n15269;
  assign n15297 = n14988 & ~n15269;
  assign n15298 = ~n15296_1 & ~n15297;
  assign n15299 = ~n15294 & ~n15298;
  assign n15300 = ~n15295 & ~n15299;
  assign n15301_1 = n13727 & ~n15300;
  assign n15302 = n13730 & ~n15290;
  assign n15303 = ~n15301_1 & ~n15302;
  assign n15304 = n13722 & ~n15300;
  assign n15305 = n13717 & ~n15300;
  assign n15306_1 = n13719 & ~n15290;
  assign n15307 = n13725 & ~n15290;
  assign n15308 = ~n15306_1 & ~n15307;
  assign n15309 = ~n15304 & ~n15305;
  assign n15310 = n15308 & n15309;
  assign n15311_1 = ~n15291_1 & ~n15292;
  assign n15312 = n15303 & n15311_1;
  assign n15313 = n15310 & n15312;
  assign n15314 = P3_REG1_REG_26_ & n13691_1;
  assign n15315 = P3_REG0_REG_26_ & n13689;
  assign n15316_1 = P3_REG2_REG_26_ & n13693;
  assign n15317 = P3_REG3_REG_25_ & n15262;
  assign n15318 = ~P3_REG3_REG_26_ & n15317;
  assign n15319 = P3_REG3_REG_26_ & ~n15317;
  assign n15320 = ~n15318 & ~n15319;
  assign n15321_1 = n13687 & ~n15320;
  assign n15322 = ~n15314 & ~n15315;
  assign n15323 = ~n15316_1 & n15322;
  assign n15324 = ~n15321_1 & n15323;
  assign n15325 = n13680 & ~n15324;
  assign n15326_1 = n13711_1 & ~n15300;
  assign n15327 = ~n15325 & ~n15326_1;
  assign n15328 = ~n15022 & n15327;
  assign n15329 = ~n14988 & n15274;
  assign n15330 = n14988 & ~n15274;
  assign n15331_1 = ~n15329 & ~n15330;
  assign n15332 = n13699 & n15331_1;
  assign n15333 = n15313 & n15328;
  assign n15334 = ~n15332 & n15333;
  assign n15335 = n13658 & ~n15334;
  assign n15336_1 = P3_REG0_REG_25_ & ~n13658;
  assign n1246 = n15335 | n15336_1;
  assign n15338 = ~n14988 & ~n15324;
  assign n15339 = n14988 & n15324;
  assign n15340 = ~n15338 & ~n15339;
  assign n15341_1 = ~n15284 & ~n15287;
  assign n15342 = ~n15283 & ~n15341_1;
  assign n15343 = n15340 & n15342;
  assign n15344 = ~n15340 & ~n15342;
  assign n15345 = ~n15343 & ~n15344;
  assign n15346_1 = n13733 & ~n15345;
  assign n15347 = n13781_1 & ~n15269;
  assign n15348 = n15294 & ~n15297;
  assign n15349 = n14988 & ~n15324;
  assign n15350 = n14988 & ~n15296_1;
  assign n15351_1 = ~n15296_1 & ~n15324;
  assign n15352 = ~n15350 & ~n15351_1;
  assign n15353 = ~n15348 & ~n15349;
  assign n15354 = ~n15352 & n15353;
  assign n15355 = ~n15294 & ~n15296_1;
  assign n15356_1 = ~n15297 & ~n15355;
  assign n15357 = n15340 & n15356_1;
  assign n15358 = ~n15354 & ~n15357;
  assign n15359 = n13727 & n15358;
  assign n15360 = n13730 & ~n15345;
  assign n15361_1 = ~n15359 & ~n15360;
  assign n15362 = n13722 & n15358;
  assign n15363 = n13717 & n15358;
  assign n15364 = n13719 & ~n15345;
  assign n15365 = n13725 & ~n15345;
  assign n15366_1 = ~n15364 & ~n15365;
  assign n15367 = ~n15362 & ~n15363;
  assign n15368 = n15366_1 & n15367;
  assign n15369 = ~n15346_1 & ~n15347;
  assign n15370 = n15361_1 & n15369;
  assign n15371_1 = n15368 & n15370;
  assign n15372 = P3_REG1_REG_27_ & n13691_1;
  assign n15373 = P3_REG0_REG_27_ & n13689;
  assign n15374 = P3_REG2_REG_27_ & n13693;
  assign n15375 = P3_REG3_REG_26_ & n15317;
  assign n15376_1 = ~P3_REG3_REG_27_ & n15375;
  assign n15377 = P3_REG3_REG_27_ & ~n15375;
  assign n15378 = ~n15376_1 & ~n15377;
  assign n15379 = n13687 & ~n15378;
  assign n15380 = ~n15372 & ~n15373;
  assign n15381_1 = ~n15374 & n15380;
  assign n15382 = ~n15379 & n15381_1;
  assign n15383 = n13680 & ~n15382;
  assign n15384 = n13711_1 & n15358;
  assign n15385 = ~n15383 & ~n15384;
  assign n15386_1 = ~n15022 & n15385;
  assign n15387 = ~n14988 & n15329;
  assign n15388 = n14988 & ~n15329;
  assign n15389 = ~n15387 & ~n15388;
  assign n15390 = n13699 & n15389;
  assign n15391_1 = n15371_1 & n15386_1;
  assign n15392 = ~n15390 & n15391_1;
  assign n15393 = n13658 & ~n15392;
  assign n15394 = P3_REG0_REG_26_ & ~n13658;
  assign n1251 = n15393 | n15394;
  assign n15396_1 = ~n14988 & ~n15382;
  assign n15397 = n14988 & n15382;
  assign n15398 = ~n15396_1 & ~n15397;
  assign n15399 = ~n15339 & ~n15398;
  assign n15400 = ~n15338 & n15342;
  assign n15401_1 = n15399 & ~n15400;
  assign n15402 = ~n15338 & n15398;
  assign n15403 = ~n15339 & ~n15342;
  assign n15404 = n15402 & ~n15403;
  assign n15405 = ~n15401_1 & ~n15404;
  assign n15406_1 = n13733 & ~n15405;
  assign n15407 = n13781_1 & ~n15324;
  assign n15408 = ~n15242 & ~n15297;
  assign n15409 = ~n15352 & ~n15408;
  assign n15410 = n15293 & ~n15352;
  assign n15411_1 = ~n15409 & ~n15410;
  assign n15412 = ~n15349 & n15411_1;
  assign n15413 = ~n15398 & n15412;
  assign n15414 = n15398 & ~n15412;
  assign n15415 = ~n15413 & ~n15414;
  assign n15416_1 = n13727 & ~n15415;
  assign n15417 = n13730 & ~n15405;
  assign n15418 = ~n15416_1 & ~n15417;
  assign n15419 = n13722 & ~n15415;
  assign n15420 = n13717 & ~n15415;
  assign n15421_1 = n13719 & ~n15405;
  assign n15422 = n13725 & ~n15405;
  assign n15423 = ~n15421_1 & ~n15422;
  assign n15424 = ~n15419 & ~n15420;
  assign n15425 = n15423 & n15424;
  assign n15426_1 = ~n15406_1 & ~n15407;
  assign n15427 = n15418 & n15426_1;
  assign n15428 = n15425 & n15427;
  assign n15429 = P3_REG1_REG_28_ & n13691_1;
  assign n15430 = P3_REG0_REG_28_ & n13689;
  assign n15431_1 = P3_REG2_REG_28_ & n13693;
  assign n15432 = P3_REG3_REG_27_ & n15375;
  assign n15433 = ~P3_REG3_REG_28_ & n15432;
  assign n15434 = P3_REG3_REG_28_ & ~n15432;
  assign n15435 = ~n15433 & ~n15434;
  assign n15436_1 = n13687 & ~n15435;
  assign n15437 = ~n15429 & ~n15430;
  assign n15438 = ~n15431_1 & n15437;
  assign n15439 = ~n15436_1 & n15438;
  assign n15440 = n13680 & ~n15439;
  assign n15441_1 = n13711_1 & ~n15415;
  assign n15442 = ~n15440 & ~n15441_1;
  assign n15443 = ~n15022 & n15442;
  assign n15444 = ~n14988 & n15387;
  assign n15445 = n14988 & ~n15387;
  assign n15446_1 = ~n15444 & ~n15445;
  assign n15447 = n13699 & n15446_1;
  assign n15448 = n15428 & n15443;
  assign n15449 = ~n15447 & n15448;
  assign n15450 = n13658 & ~n15449;
  assign n15451_1 = P3_REG0_REG_27_ & ~n13658;
  assign n1256 = n15450 | n15451_1;
  assign n15453 = ~n14988 & ~n15439;
  assign n15454 = n14988 & n15439;
  assign n15455 = ~n15453 & ~n15454;
  assign n15456_1 = ~n15338 & n15382;
  assign n15457 = ~n14988 & ~n15456_1;
  assign n15458 = n15338 & ~n15382;
  assign n15459 = ~n15457 & ~n15458;
  assign n15460 = ~n15397 & n15403;
  assign n15461_1 = n15459 & ~n15460;
  assign n15462 = ~n15455 & ~n15461_1;
  assign n15463 = n15455 & n15461_1;
  assign n15464 = ~n15462 & ~n15463;
  assign n15465 = n13733 & ~n15464;
  assign n15466_1 = n13781_1 & ~n15382;
  assign n15467 = ~n14988 & n15382;
  assign n15468 = n15349 & ~n15467;
  assign n15469 = ~n15241_1 & ~n15467;
  assign n15470 = ~n15239 & ~n15352;
  assign n15471_1 = n15469 & n15470;
  assign n15472 = n15409 & ~n15467;
  assign n15473 = n14988 & ~n15382;
  assign n15474 = ~n15472 & ~n15473;
  assign n15475 = ~n15468 & ~n15471_1;
  assign n15476_1 = n15474 & n15475;
  assign n15477 = ~n15455 & n15476_1;
  assign n15478 = n15455 & ~n15476_1;
  assign n15479 = ~n15477 & ~n15478;
  assign n15480 = n13727 & ~n15479;
  assign n15481_1 = n13730 & ~n15464;
  assign n15482 = ~n15480 & ~n15481_1;
  assign n15483 = n13722 & ~n15479;
  assign n15484 = n13717 & ~n15479;
  assign n15485 = n13719 & ~n15464;
  assign n15486_1 = n13725 & ~n15464;
  assign n15487 = ~n15485 & ~n15486_1;
  assign n15488 = ~n15483 & ~n15484;
  assign n15489 = n15487 & n15488;
  assign n15490 = ~n15465 & ~n15466_1;
  assign n15491_1 = n15482 & n15490;
  assign n15492 = n15489 & n15491_1;
  assign n15493 = P3_REG0_REG_29_ & n13689;
  assign n15494 = P3_REG1_REG_29_ & n13691_1;
  assign n15495 = P3_REG2_REG_29_ & n13693;
  assign n15496_1 = P3_REG3_REG_28_ & P3_REG3_REG_27_;
  assign n15497 = n15375 & n15496_1;
  assign n15498 = n13687 & n15497;
  assign n15499 = ~n15493 & ~n15494;
  assign n15500 = ~n15495 & n15499;
  assign n15501_1 = ~n15498 & n15500;
  assign n15502 = n13680 & ~n15501_1;
  assign n15503 = n13711_1 & ~n15479;
  assign n15504 = ~n15502 & ~n15503;
  assign n15505 = ~n15022 & n15504;
  assign n15506_1 = ~n14988 & n15444;
  assign n15507 = n14988 & ~n15444;
  assign n15508 = ~n15506_1 & ~n15507;
  assign n15509 = n13699 & n15508;
  assign n15510 = n15492 & n15505;
  assign n15511_1 = ~n15509 & n15510;
  assign n15512 = n13658 & ~n15511_1;
  assign n15513 = P3_REG0_REG_28_ & ~n13658;
  assign n1261 = n15512 | n15513;
  assign n15515 = n14988 & ~n15476_1;
  assign n15516_1 = ~n15439 & ~n15476_1;
  assign n15517 = n14988 & ~n15439;
  assign n15518 = ~n15515 & ~n15516_1;
  assign n15519 = ~n15517 & n15518;
  assign n15520 = n14988 & n15501_1;
  assign n15521_1 = ~n14988 & ~n15501_1;
  assign n15522 = ~n15520 & ~n15521_1;
  assign n15523 = n15519 & ~n15522;
  assign n15524 = ~n15519 & n15522;
  assign n15525 = ~n15523 & ~n15524;
  assign n15526_1 = n13711_1 & ~n15525;
  assign n15527 = ~n15022 & ~n15526_1;
  assign n15528 = n13722 & ~n15525;
  assign n15529 = n13717 & ~n15525;
  assign n15530 = n15439 & n15522;
  assign n15531_1 = n14988 & n15530;
  assign n15532 = ~n15439 & ~n15522;
  assign n15533 = ~n14988 & n15532;
  assign n15534 = ~n15531_1 & ~n15533;
  assign n15535 = ~n15454 & ~n15522;
  assign n15536_1 = ~n15461_1 & n15535;
  assign n15537 = ~n15453 & n15459;
  assign n15538 = ~n15460 & n15522;
  assign n15539 = n15537 & n15538;
  assign n15540 = n15534 & ~n15536_1;
  assign n15541_1 = ~n15539 & n15540;
  assign n15542 = n13719 & ~n15541_1;
  assign n15543 = n13725 & ~n15541_1;
  assign n15544 = ~n15542 & ~n15543;
  assign n15545 = ~n15528 & ~n15529;
  assign n15546_1 = n15544 & n15545;
  assign n15547 = n13781_1 & ~n15439;
  assign n15548 = ~P3_B_REG & n13664;
  assign n15549 = ~n13665 & ~n15548;
  assign n15550 = n13679 & ~n15549;
  assign n15551_1 = P3_REG1_REG_30_ & n13691_1;
  assign n15552 = P3_REG0_REG_30_ & n13689;
  assign n15553 = P3_REG2_REG_30_ & n13693;
  assign n15554 = ~n15551_1 & ~n15552;
  assign n15555 = ~n15553 & n15554;
  assign n15556_1 = n15550 & ~n15555;
  assign n15557 = n13733 & ~n15541_1;
  assign n15558 = n13730 & ~n15541_1;
  assign n15559 = n13727 & ~n15525;
  assign n15560 = ~n15547 & ~n15556_1;
  assign n15561_1 = ~n15557 & n15560;
  assign n15562 = ~n15558 & n15561_1;
  assign n15563 = ~n15559 & n15562;
  assign n15564 = n15546_1 & n15563;
  assign n15565 = ~n14988 & n15506_1;
  assign n15566_1 = n14988 & ~n15506_1;
  assign n15567 = ~n15565 & ~n15566_1;
  assign n15568 = n13699 & n15567;
  assign n15569 = n15527 & n15564;
  assign n15570 = ~n15568 & n15569;
  assign n15571_1 = n13658 & ~n15570;
  assign n15572 = P3_REG0_REG_29_ & ~n13658;
  assign n1266 = n15571_1 | n15572;
  assign n15574 = P3_REG1_REG_31_ & n13691_1;
  assign n15575 = P3_REG0_REG_31_ & n13689;
  assign n15576_1 = P3_REG2_REG_31_ & n13693;
  assign n15577 = ~n15574 & ~n15575;
  assign n15578 = ~n15576_1 & n15577;
  assign n15579 = n15550 & ~n15578;
  assign n15580 = ~n14988 & n15565;
  assign n15581_1 = n14988 & ~n15565;
  assign n15582 = ~n15580 & ~n15581_1;
  assign n15583 = n13699 & n15582;
  assign n15584 = ~n15022 & ~n15579;
  assign n15585 = ~n15583 & n15584;
  assign n15586_1 = n13658 & ~n15585;
  assign n15587 = P3_REG0_REG_30_ & ~n13658;
  assign n1271 = n15586_1 | n15587;
  assign n15589 = ~n14988 & n15580;
  assign n15590 = n14988 & ~n15580;
  assign n15591_1 = ~n15589 & ~n15590;
  assign n15592 = n15584 & ~n15591_1;
  assign n15593 = ~n13699 & ~n15022;
  assign n15594 = ~n15579 & n15593;
  assign n15595 = ~n15592 & ~n15594;
  assign n15596_1 = n13658 & n15595;
  assign n15597 = P3_REG0_REG_31_ & ~n13658;
  assign n1276 = n15596_1 | n15597;
  assign n15599 = n13525 & ~n13574;
  assign n15600 = n13657 & n15599;
  assign n15601_1 = ~n13740 & n15600;
  assign n15602 = P3_REG1_REG_0_ & ~n15600;
  assign n1281 = n15601_1 | n15602;
  assign n15604 = ~n13796_1 & n15600;
  assign n15605 = P3_REG1_REG_1_ & ~n15600;
  assign n1286 = n15604 | n15605;
  assign n15607 = ~n13858 & n15600;
  assign n15608 = P3_REG1_REG_2_ & ~n15600;
  assign n1291 = n15607 | n15608;
  assign n15610 = ~n13923 & n15600;
  assign n15611_1 = P3_REG1_REG_3_ & ~n15600;
  assign n1296 = n15610 | n15611_1;
  assign n15613 = ~n13993 & n15600;
  assign n15614 = P3_REG1_REG_4_ & ~n15600;
  assign n1301 = n15613 | n15614;
  assign n15616_1 = ~n14057 & n15600;
  assign n15617 = P3_REG1_REG_5_ & ~n15600;
  assign n1306 = n15616_1 | n15617;
  assign n15619 = ~n14130 & n15600;
  assign n15620 = P3_REG1_REG_6_ & ~n15600;
  assign n1311 = n15619 | n15620;
  assign n15622 = ~n14199 & n15600;
  assign n15623 = P3_REG1_REG_7_ & ~n15600;
  assign n1316 = n15622 | n15623;
  assign n15625 = ~n14267 & n15600;
  assign n15626_1 = P3_REG1_REG_8_ & ~n15600;
  assign n1321 = n15625 | n15626_1;
  assign n15628 = ~n14334 & n15600;
  assign n15629 = P3_REG1_REG_9_ & ~n15600;
  assign n1326 = n15628 | n15629;
  assign n15631_1 = ~n14398 & n15600;
  assign n15632 = P3_REG1_REG_10_ & ~n15600;
  assign n1331 = n15631_1 | n15632;
  assign n15634 = ~n14468 & n15600;
  assign n15635 = P3_REG1_REG_11_ & ~n15600;
  assign n1336 = n15634 | n15635;
  assign n15637 = ~n14534 & n15600;
  assign n15638 = P3_REG1_REG_12_ & ~n15600;
  assign n1341 = n15637 | n15638;
  assign n15640 = ~n14598 & n15600;
  assign n15641_1 = P3_REG1_REG_13_ & ~n15600;
  assign n1346 = n15640 | n15641_1;
  assign n15643 = ~n14661_1 & n15600;
  assign n15644 = P3_REG1_REG_14_ & ~n15600;
  assign n1351 = n15643 | n15644;
  assign n15646_1 = ~n14722 & n15600;
  assign n15647 = P3_REG1_REG_15_ & ~n15600;
  assign n1356 = n15646_1 | n15647;
  assign n15649 = ~n14789 & n15600;
  assign n15650 = P3_REG1_REG_16_ & ~n15600;
  assign n1361 = n15649 | n15650;
  assign n15652 = ~n14857 & n15600;
  assign n15653 = P3_REG1_REG_17_ & ~n15600;
  assign n1366 = n15652 | n15653;
  assign n15655 = ~n14923 & n15600;
  assign n15656_1 = P3_REG1_REG_18_ & ~n15600;
  assign n1371 = n15655 | n15656_1;
  assign n15658 = ~n14984 & n15600;
  assign n15659 = P3_REG1_REG_19_ & ~n15600;
  assign n1376 = n15658 | n15659;
  assign n15661_1 = ~n15043 & n15600;
  assign n15662 = P3_REG1_REG_20_ & ~n15600;
  assign n1381 = n15661_1 | n15662;
  assign n15664 = ~n15100 & n15600;
  assign n15665 = P3_REG1_REG_21_ & ~n15600;
  assign n1386 = n15664 | n15665;
  assign n15667 = ~n15160 & n15600;
  assign n15668 = P3_REG1_REG_22_ & ~n15600;
  assign n1391 = n15667 | n15668;
  assign n15670 = ~n15217 & n15600;
  assign n15671_1 = P3_REG1_REG_23_ & ~n15600;
  assign n1396 = n15670 | n15671_1;
  assign n15673 = ~n15279 & n15600;
  assign n15674 = P3_REG1_REG_24_ & ~n15600;
  assign n1401 = n15673 | n15674;
  assign n15676_1 = ~n15334 & n15600;
  assign n15677 = P3_REG1_REG_25_ & ~n15600;
  assign n1406 = n15676_1 | n15677;
  assign n15679 = ~n15392 & n15600;
  assign n15680 = P3_REG1_REG_26_ & ~n15600;
  assign n1411 = n15679 | n15680;
  assign n15682 = ~n15449 & n15600;
  assign n15683 = P3_REG1_REG_27_ & ~n15600;
  assign n1416 = n15682 | n15683;
  assign n15685 = ~n15511_1 & n15600;
  assign n15686_1 = P3_REG1_REG_28_ & ~n15600;
  assign n1421 = n15685 | n15686_1;
  assign n15688 = ~n15570 & n15600;
  assign n15689 = P3_REG1_REG_29_ & ~n15600;
  assign n1426 = n15688 | n15689;
  assign n15691_1 = ~n15585 & n15600;
  assign n15692 = P3_REG1_REG_30_ & ~n15600;
  assign n1431 = n15691_1 | n15692;
  assign n15694 = n15595 & n15600;
  assign n15695 = P3_REG1_REG_31_ & ~n15600;
  assign n1436 = n15694 | n15695;
  assign n15697 = n13593 & n13699;
  assign n15698 = n13584 & n13676_1;
  assign n15699 = ~n13594 & n13679;
  assign n15700 = n13574 & ~n15699;
  assign n15701_1 = ~n13578 & n15700;
  assign n15702 = n13656_1 & n15701_1;
  assign n15703 = ~n15698 & ~n15702;
  assign n15704 = n13525 & ~n15703;
  assign n15705 = n15697 & n15704;
  assign n15706_1 = ~n13671_1 & n15705;
  assign n15707 = ~n13584 & n13676_1;
  assign n15708 = ~n13674 & ~n15707;
  assign n15709 = n15704 & ~n15708;
  assign n15710 = ~n13671_1 & n15709;
  assign n15711_1 = ~n13739 & n15704;
  assign n15712 = P3_REG2_REG_0_ & ~n15704;
  assign n15713 = ~n15711_1 & ~n15712;
  assign n15714 = ~n15706_1 & ~n15710;
  assign n15715 = n15713 & n15714;
  assign n15716_1 = n15698 & n15704;
  assign n15717 = P3_REG3_REG_0_ & n15716_1;
  assign n15718 = n13680 & n15704;
  assign n15719 = ~n13697 & n15718;
  assign n15720 = ~n13587 & n13732;
  assign n15721_1 = n15704 & n15720;
  assign n15722 = ~n13710 & n15721_1;
  assign n15723 = ~n15717 & ~n15719;
  assign n15724 = ~n15722 & n15723;
  assign n1441 = ~n15715 | ~n15724;
  assign n15726_1 = ~n13760 & n15705;
  assign n15727 = ~n13757 & n15709;
  assign n15728 = ~n13795 & n15704;
  assign n15729 = P3_REG2_REG_1_ & ~n15704;
  assign n15730 = ~n15728 & ~n15729;
  assign n15731_1 = ~n15726_1 & ~n15727;
  assign n15732 = n15730 & n15731_1;
  assign n15733 = P3_REG3_REG_1_ & n15716_1;
  assign n15734 = ~n13750 & n15718;
  assign n15735 = ~n13769 & n15721_1;
  assign n15736_1 = ~n15733 & ~n15734;
  assign n15737 = ~n15735 & n15736_1;
  assign n1446 = ~n15732 | ~n15737;
  assign n15739 = n13817 & n15705;
  assign n15740 = ~n13813 & n15709;
  assign n15741_1 = ~n13857 & n15704;
  assign n15742 = P3_REG2_REG_2_ & ~n15704;
  assign n15743 = ~n15741_1 & ~n15742;
  assign n15744 = ~n15739 & ~n15740;
  assign n15745 = n15743 & n15744;
  assign n15746_1 = P3_REG3_REG_2_ & n15716_1;
  assign n15747 = ~n13806_1 & n15718;
  assign n15748 = n13831_1 & n15721_1;
  assign n15749 = ~n15746_1 & ~n15747;
  assign n15750 = ~n15748 & n15749;
  assign n1451 = ~n15745 | ~n15750;
  assign n15752 = n13881_1 & n15705;
  assign n15753 = ~n13878 & n15709;
  assign n15754 = ~n13922 & n15704;
  assign n15755 = P3_REG2_REG_3_ & ~n15704;
  assign n15756_1 = ~n15754 & ~n15755;
  assign n15757 = ~n15752 & ~n15753;
  assign n15758 = n15756_1 & n15757;
  assign n15759 = ~P3_REG3_REG_3_ & n15716_1;
  assign n15760 = ~n13871_1 & n15718;
  assign n15761_1 = ~n13896_1 & n15721_1;
  assign n15762 = ~n15759 & ~n15760;
  assign n15763 = ~n15761_1 & n15762;
  assign n1456 = ~n15758 | ~n15763;
  assign n15765 = n13947 & n15705;
  assign n15766_1 = ~n13944 & n15709;
  assign n15767 = ~n13992 & n15704;
  assign n15768 = P3_REG2_REG_4_ & ~n15704;
  assign n15769 = ~n15767 & ~n15768;
  assign n15770 = ~n15765 & ~n15766_1;
  assign n15771_1 = n15769 & n15770;
  assign n15772 = ~n13864 & n15716_1;
  assign n15773 = ~n13937 & n15718;
  assign n15774 = ~n13963 & n15721_1;
  assign n15775 = ~n15772 & ~n15773;
  assign n15776_1 = ~n15774 & n15775;
  assign n1461 = ~n15771_1 | ~n15776_1;
  assign n15778 = n14017 & n15705;
  assign n15779 = ~n14014 & n15709;
  assign n15780 = ~n15778 & ~n15779;
  assign n15781_1 = ~n13930 & n15716_1;
  assign n15782 = ~n14007 & n15718;
  assign n15783 = n14032 & n15721_1;
  assign n15784 = ~n15781_1 & ~n15782;
  assign n15785 = ~n15783 & n15784;
  assign n15786_1 = ~n14056_1 & n15704;
  assign n15787 = P3_REG2_REG_5_ & ~n15704;
  assign n15788 = ~n15786_1 & ~n15787;
  assign n15789 = n15780 & n15785;
  assign n1466 = ~n15788 | ~n15789;
  assign n15791_1 = n14102 & n15705;
  assign n15792 = ~n14066_1 & n15709;
  assign n15793 = ~n15791_1 & ~n15792;
  assign n15794 = ~n14000 & n15716_1;
  assign n15795 = ~n14098 & n15718;
  assign n15796_1 = ~n14086_1 & n15721_1;
  assign n15797 = ~n15794 & ~n15795;
  assign n15798 = ~n15796_1 & n15797;
  assign n15799 = ~n14129 & n15704;
  assign n15800 = P3_REG2_REG_6_ & ~n15704;
  assign n15801_1 = ~n15799 & ~n15800;
  assign n15802 = n15793 & n15798;
  assign n1471 = ~n15801_1 | ~n15802;
  assign n15804 = n14169 & n15705;
  assign n15805 = ~n14139 & n15709;
  assign n15806_1 = ~n15804 & ~n15805;
  assign n15807 = ~n14091_1 & n15716_1;
  assign n15808 = ~n14165 & n15718;
  assign n15809 = n14153 & n15721_1;
  assign n15810 = ~n15807 & ~n15808;
  assign n15811_1 = ~n15809 & n15810;
  assign n15812 = ~n14198 & n15704;
  assign n15813 = P3_REG2_REG_7_ & ~n15704;
  assign n15814 = ~n15812 & ~n15813;
  assign n15815 = n15806_1 & n15811_1;
  assign n1476 = ~n15814 | ~n15815;
  assign n15817 = n14212 & n15705;
  assign n15818 = ~n14208 & n15709;
  assign n15819 = ~n15817 & ~n15818;
  assign n15820 = ~n14158 & n15716_1;
  assign n15821_1 = ~n14224 & n15718;
  assign n15822 = ~n14240 & n15721_1;
  assign n15823 = ~n15820 & ~n15821_1;
  assign n15824 = ~n15822 & n15823;
  assign n15825 = ~n14266_1 & n15704;
  assign n15826_1 = P3_REG2_REG_8_ & ~n15704;
  assign n15827 = ~n15825 & ~n15826_1;
  assign n15828 = n15819 & n15824;
  assign n1481 = ~n15827 | ~n15828;
  assign n15830 = n14280 & n15705;
  assign n15831_1 = ~n14276_1 & n15709;
  assign n15832 = ~n15830 & ~n15831_1;
  assign n15833 = ~n14220 & n15716_1;
  assign n15834 = ~n14292 & n15718;
  assign n15835 = ~n14304 & n15721_1;
  assign n15836_1 = ~n15833 & ~n15834;
  assign n15837 = ~n15835 & n15836_1;
  assign n15838 = ~n14333 & n15704;
  assign n15839 = P3_REG2_REG_9_ & ~n15704;
  assign n15840 = ~n15838 & ~n15839;
  assign n15841_1 = n15832 & n15837;
  assign n1486 = ~n15840 | ~n15841_1;
  assign n15843 = ~n14288 & n15716_1;
  assign n15844 = ~n14348 & n15718;
  assign n15845 = n14368 & n15721_1;
  assign n15846_1 = ~n14355 & n15709;
  assign n15847 = n14373 & n15705;
  assign n15848 = ~n15843 & ~n15844;
  assign n15849 = ~n15845 & n15848;
  assign n15850 = ~n15846_1 & n15849;
  assign n15851_1 = ~n15847 & n15850;
  assign n15852 = ~n14397 & n15704;
  assign n15853 = P3_REG2_REG_10_ & ~n15704;
  assign n15854 = ~n15852 & ~n15853;
  assign n1491 = ~n15851_1 | ~n15854;
  assign n15856_1 = ~n14344 & n15716_1;
  assign n15857 = ~n14458 & n15718;
  assign n15858 = ~n14433 & n15721_1;
  assign n15859 = ~n14407 & n15709;
  assign n15860 = n14463 & n15705;
  assign n15861_1 = ~n15856_1 & ~n15857;
  assign n15862 = ~n15858 & n15861_1;
  assign n15863 = ~n15859 & n15862;
  assign n15864 = ~n15860 & n15863;
  assign n15865 = ~n14446_1 & n15704;
  assign n15866_1 = P3_REG2_REG_11_ & ~n15704;
  assign n15867 = ~n15865 & ~n15866_1;
  assign n1496 = ~n15864 | ~n15867;
  assign n15869 = ~n14454 & n15716_1;
  assign n15870 = ~n14524 & n15718;
  assign n15871_1 = ~n14499 & n15721_1;
  assign n15872 = ~n14477 & n15709;
  assign n15873 = n14529 & n15705;
  assign n15874 = ~n15869 & ~n15870;
  assign n15875 = ~n15871_1 & n15874;
  assign n15876_1 = ~n15872 & n15875;
  assign n15877 = ~n15873 & n15876_1;
  assign n15878 = ~n14512 & n15704;
  assign n15879 = P3_REG2_REG_12_ & ~n15704;
  assign n15880 = ~n15878 & ~n15879;
  assign n1501 = ~n15877 | ~n15880;
  assign n15882 = ~n14520 & n15716_1;
  assign n15883 = ~n14588 & n15718;
  assign n15884 = n14563 & n15721_1;
  assign n15885 = ~n14543 & n15709;
  assign n15886_1 = n14593 & n15705;
  assign n15887 = ~n15882 & ~n15883;
  assign n15888 = ~n15884 & n15887;
  assign n15889 = ~n15885 & n15888;
  assign n15890 = ~n15886_1 & n15889;
  assign n15891_1 = ~n14576_1 & n15704;
  assign n15892 = P3_REG2_REG_13_ & ~n15704;
  assign n15893 = ~n15891_1 & ~n15892;
  assign n1506 = ~n15890 | ~n15893;
  assign n15895 = ~n14584 & n15716_1;
  assign n15896_1 = ~n14651_1 & n15718;
  assign n15897 = ~n14626_1 & n15721_1;
  assign n15898 = ~n14609 & n15709;
  assign n15899 = n14656_1 & n15705;
  assign n15900 = ~n15895 & ~n15896_1;
  assign n15901_1 = ~n15897 & n15900;
  assign n15902 = ~n15898 & n15901_1;
  assign n15903 = ~n15899 & n15902;
  assign n15904 = ~n14639 & n15704;
  assign n15905 = P3_REG2_REG_14_ & ~n15704;
  assign n15906_1 = ~n15904 & ~n15905;
  assign n1511 = ~n15903 | ~n15906_1;
  assign n15908 = ~n14647 & n15716_1;
  assign n15909 = ~n14712 & n15718;
  assign n15910 = ~n14687 & n15721_1;
  assign n15911_1 = ~n14670 & n15709;
  assign n15912 = n14717 & n15705;
  assign n15913 = ~n15908 & ~n15909;
  assign n15914 = ~n15910 & n15913;
  assign n15915 = ~n15911_1 & n15914;
  assign n15916_1 = ~n15912 & n15915;
  assign n15917 = ~n14700 & n15704;
  assign n15918 = P3_REG2_REG_15_ & ~n15704;
  assign n15919 = ~n15917 & ~n15918;
  assign n1516 = ~n15916_1 | ~n15919;
  assign n15921_1 = ~n14708 & n15716_1;
  assign n15922 = ~n14779 & n15718;
  assign n15923 = ~n14754 & n15721_1;
  assign n15924 = ~n14767 & n15704;
  assign n15925 = P3_REG2_REG_16_ & ~n15704;
  assign n15926_1 = ~n15924 & ~n15925;
  assign n15927 = ~n15921_1 & ~n15922;
  assign n15928 = ~n15923 & n15927;
  assign n15929 = n15926_1 & n15928;
  assign n15930 = n14784 & n15705;
  assign n15931_1 = ~n14731_1 & n15709;
  assign n15932 = ~n15930 & ~n15931_1;
  assign n1521 = ~n15929 | ~n15932;
  assign n15934 = ~n14775 & n15716_1;
  assign n15935 = ~n14846_1 & n15718;
  assign n15936_1 = n14822 & n15721_1;
  assign n15937 = n14854 & n15705;
  assign n15938 = ~n15934 & ~n15935;
  assign n15939 = ~n15936_1 & n15938;
  assign n15940 = ~n15937 & n15939;
  assign n15941_1 = ~n14835 & n15704;
  assign n15942 = P3_REG2_REG_17_ & ~n15704;
  assign n15943 = ~n15941_1 & ~n15942;
  assign n15944 = ~n14798 & n15709;
  assign n15945 = n15943 & ~n15944;
  assign n1526 = ~n15940 | ~n15945;
  assign n15947 = ~n14842 & n15716_1;
  assign n15948 = ~n14912 & n15718;
  assign n15949 = ~n14888 & n15721_1;
  assign n15950 = n14920 & n15705;
  assign n15951_1 = ~n15947 & ~n15948;
  assign n15952 = ~n15949 & n15951_1;
  assign n15953 = ~n15950 & n15952;
  assign n15954 = ~n14901_1 & n15704;
  assign n15955 = P3_REG2_REG_18_ & ~n15704;
  assign n15956_1 = ~n15954 & ~n15955;
  assign n15957 = ~n14866_1 & n15709;
  assign n15958 = n15956_1 & ~n15957;
  assign n1531 = ~n15953 | ~n15958;
  assign n15960 = ~n14908 & n15716_1;
  assign n15961_1 = ~n14974 & n15718;
  assign n15962 = ~n14949 & n15721_1;
  assign n15963 = ~n14929 & n15709;
  assign n15964 = n14979 & n15705;
  assign n15965 = ~n15960 & ~n15961_1;
  assign n15966_1 = ~n15962 & n15965;
  assign n15967 = ~n15963 & n15966_1;
  assign n15968 = ~n15964 & n15967;
  assign n15969 = ~n14962 & n15704;
  assign n15970 = P3_REG2_REG_19_ & ~n15704;
  assign n15971_1 = ~n15969 & ~n15970;
  assign n1536 = ~n15968 | ~n15971_1;
  assign n15973 = ~n14970 & n15716_1;
  assign n15974 = ~n15033 & n15718;
  assign n15975 = n15008 & n15721_1;
  assign n15976_1 = n14988 & n15709;
  assign n15977 = n15038 & n15705;
  assign n15978 = ~n15973 & ~n15974;
  assign n15979 = ~n15975 & n15978;
  assign n15980 = ~n15976_1 & n15979;
  assign n15981_1 = ~n15977 & n15980;
  assign n15982 = ~n15021_1 & n15704;
  assign n15983 = P3_REG2_REG_20_ & ~n15704;
  assign n15984 = ~n15982 & ~n15983;
  assign n1541 = ~n15981_1 | ~n15984;
  assign n15986_1 = ~n15029 & n15716_1;
  assign n15987 = ~n15090 & n15718;
  assign n15988 = n15066_1 & n15721_1;
  assign n15989 = n15095 & n15705;
  assign n15990 = ~n15986_1 & ~n15987;
  assign n15991_1 = ~n15988 & n15990;
  assign n15992 = ~n15976_1 & n15991_1;
  assign n15993 = ~n15989 & n15992;
  assign n15994 = ~n15079 & n15704;
  assign n15995 = P3_REG2_REG_21_ & ~n15704;
  assign n15996_1 = ~n15994 & ~n15995;
  assign n1546 = ~n15993 | ~n15996_1;
  assign n15998 = ~n15086_1 & n15716_1;
  assign n15999 = ~n15150 & n15718;
  assign n16000 = ~n15126_1 & n15721_1;
  assign n16001_1 = n15155 & n15705;
  assign n16002 = ~n15998 & ~n15999;
  assign n16003 = ~n16000 & n16002;
  assign n16004 = ~n15976_1 & n16003;
  assign n16005 = ~n16001_1 & n16004;
  assign n16006_1 = ~n15139 & n15704;
  assign n16007 = P3_REG2_REG_22_ & ~n15704;
  assign n16008 = ~n16006_1 & ~n16007;
  assign n1551 = ~n16005 | ~n16008;
  assign n16010 = ~n15146_1 & n15716_1;
  assign n16011_1 = ~n15207 & n15718;
  assign n16012 = ~n15183 & n15721_1;
  assign n16013 = ~n15196_1 & n15704;
  assign n16014 = P3_REG2_REG_23_ & ~n15704;
  assign n16015 = ~n16013 & ~n16014;
  assign n16016_1 = ~n16010 & ~n16011_1;
  assign n16017 = ~n16012 & n16016_1;
  assign n16018 = n16015 & n16017;
  assign n16019 = n15212 & n15705;
  assign n16020 = ~n15976_1 & ~n16019;
  assign n1556 = ~n16018 | ~n16020;
  assign n16022 = ~n15203 & n15716_1;
  assign n16023 = ~n15269 & n15718;
  assign n16024 = ~n15245 & n15721_1;
  assign n16025 = n15276_1 & n15705;
  assign n16026_1 = ~n16022 & ~n16023;
  assign n16027 = ~n16024 & n16026_1;
  assign n16028 = ~n16025 & n16027;
  assign n16029 = ~n15258 & n15704;
  assign n16030 = P3_REG2_REG_24_ & ~n15704;
  assign n16031_1 = ~n16029 & ~n16030;
  assign n16032 = ~n15976_1 & n16031_1;
  assign n1561 = ~n16028 | ~n16032;
  assign n16034 = ~n15265 & n15716_1;
  assign n16035 = ~n15324 & n15718;
  assign n16036_1 = ~n15300 & n15721_1;
  assign n16037 = n15331_1 & n15705;
  assign n16038 = ~n16034 & ~n16035;
  assign n16039 = ~n16036_1 & n16038;
  assign n16040 = ~n16037 & n16039;
  assign n16041_1 = ~n15313 & n15704;
  assign n16042 = P3_REG2_REG_25_ & ~n15704;
  assign n16043 = ~n16041_1 & ~n16042;
  assign n16044 = ~n15976_1 & n16043;
  assign n1566 = ~n16040 | ~n16044;
  assign n16046_1 = ~n15320 & n15716_1;
  assign n16047 = ~n15382 & n15718;
  assign n16048 = n15358 & n15721_1;
  assign n16049 = n15389 & n15705;
  assign n16050 = ~n16046_1 & ~n16047;
  assign n16051_1 = ~n16048 & n16050;
  assign n16052 = ~n16049 & n16051_1;
  assign n16053 = ~n15371_1 & n15704;
  assign n16054 = P3_REG2_REG_26_ & ~n15704;
  assign n16055 = ~n16053 & ~n16054;
  assign n16056_1 = ~n15976_1 & n16055;
  assign n1571 = ~n16052 | ~n16056_1;
  assign n16058 = ~n15378 & n15716_1;
  assign n16059 = ~n15439 & n15718;
  assign n16060 = ~n15415 & n15721_1;
  assign n16061_1 = ~n15428 & n15704;
  assign n16062 = P3_REG2_REG_27_ & ~n15704;
  assign n16063 = ~n16061_1 & ~n16062;
  assign n16064 = ~n16058 & ~n16059;
  assign n16065 = ~n16060 & n16064;
  assign n16066_1 = ~n15976_1 & n16065;
  assign n16067 = n16063 & n16066_1;
  assign n16068 = n15446_1 & n15705;
  assign n1576 = ~n16067 | n16068;
  assign n16070 = ~n15435 & n15716_1;
  assign n16071_1 = ~n15501_1 & n15718;
  assign n16072 = ~n15479 & n15721_1;
  assign n16073 = ~n15492 & n15704;
  assign n16074 = P3_REG2_REG_28_ & ~n15704;
  assign n16075 = ~n16073 & ~n16074;
  assign n16076_1 = ~n16070 & ~n16071_1;
  assign n16077 = ~n16072 & n16076_1;
  assign n16078 = ~n15976_1 & n16077;
  assign n16079 = n16075 & n16078;
  assign n16080 = n15508 & n15705;
  assign n1581 = ~n16079 | n16080;
  assign n16082 = n15497 & n15716_1;
  assign n16083 = ~n15525 & n15721_1;
  assign n16084 = ~n15564 & n15704;
  assign n16085 = P3_REG2_REG_29_ & ~n15704;
  assign n16086_1 = ~n16084 & ~n16085;
  assign n16087 = n15567 & n15705;
  assign n16088 = ~n15976_1 & ~n16082;
  assign n16089 = ~n16083 & n16088;
  assign n16090 = n16086_1 & n16089;
  assign n1586 = n16087 | ~n16090;
  assign n16092 = n15579 & n15704;
  assign n16093 = P3_REG2_REG_30_ & ~n15704;
  assign n16094 = ~n16092 & ~n16093;
  assign n16095 = n15582 & n15705;
  assign n16096_1 = ~n15976_1 & n16094;
  assign n1591 = n16095 | ~n16096_1;
  assign n16098 = P3_REG2_REG_31_ & ~n15704;
  assign n16099 = ~n16092 & ~n16098;
  assign n16100 = n15591_1 & n15705;
  assign n16101_1 = ~n15976_1 & n16099;
  assign n1596 = n16100 | ~n16101_1;
  assign n16103 = P3_STATE_REG & ~n13512;
  assign n16104 = n13512 & n13523;
  assign n16105 = n13524 & ~n13679;
  assign n16106_1 = n13512 & ~n16105;
  assign n16107 = ~n13665 & ~n16106_1;
  assign n2016 = ~P3_STATE_REG | n16107;
  assign n16109 = ~n16104 & ~n2016;
  assign n16110 = n16103 & ~n16109;
  assign n16111_1 = ~n13661_1 & ~n13664;
  assign n16112 = n16110 & n16111_1;
  assign n16113 = ~P3_REG2_REG_18_ & n14863;
  assign n16114 = P3_REG2_REG_19_ & n13593;
  assign n16115 = ~P3_REG2_REG_19_ & ~n13593;
  assign n16116_1 = ~n16114 & ~n16115;
  assign n16117 = P3_REG2_REG_16_ & ~n14728;
  assign n16118 = P3_REG2_REG_17_ & n16117;
  assign n16119 = ~P3_REG2_REG_17_ & ~n16117;
  assign n16120 = ~n14795 & ~n16119;
  assign n16121_1 = ~P3_REG2_REG_16_ & n14728;
  assign n16122 = ~P3_REG2_REG_17_ & n14795;
  assign n16123 = ~n16121_1 & ~n16122;
  assign n16124 = P3_REG2_REG_15_ & ~n14667;
  assign n16125 = ~P3_REG2_REG_15_ & n14667;
  assign n16126_1 = P3_REG2_REG_14_ & ~n14606_1;
  assign n16127 = ~P3_REG2_REG_14_ & n14606_1;
  assign n16128 = ~P3_REG2_REG_13_ & n14540;
  assign n16129 = P3_REG2_REG_13_ & ~n14540;
  assign n16130 = P3_REG2_REG_12_ & ~n14474;
  assign n16131_1 = P3_REG2_REG_11_ & ~n14404;
  assign n16132 = ~P3_REG2_REG_12_ & n14474;
  assign n16133 = ~n16128 & ~n16132;
  assign n16134 = n16131_1 & n16133;
  assign n16135 = ~n16129 & ~n16130;
  assign n16136_1 = ~n16134 & n16135;
  assign n16137 = ~n16128 & ~n16136_1;
  assign n16138 = ~P3_REG2_REG_11_ & n14404;
  assign n16139 = ~P3_REG2_REG_10_ & n14352;
  assign n16140 = P3_REG2_REG_10_ & ~n14352;
  assign n16141_1 = P3_REG2_REG_9_ & ~n14273;
  assign n16142 = P3_REG2_REG_8_ & ~n14205;
  assign n16143 = ~P3_REG2_REG_9_ & n14273;
  assign n16144 = ~n16139 & ~n16143;
  assign n16145 = n16142 & n16144;
  assign n16146_1 = ~n16140 & ~n16141_1;
  assign n16147 = ~n16145 & n16146_1;
  assign n16148 = ~n16139 & ~n16147;
  assign n16149 = ~P3_REG2_REG_8_ & n14205;
  assign n16150 = P3_REG2_REG_6_ & ~n14063;
  assign n16151_1 = P3_REG2_REG_7_ & n16150;
  assign n16152 = ~P3_REG2_REG_7_ & ~n16150;
  assign n16153 = ~n14136_1 & ~n16152;
  assign n16154 = ~P3_REG2_REG_6_ & n14063;
  assign n16155 = ~P3_REG2_REG_7_ & n14136_1;
  assign n16156_1 = ~n16154 & ~n16155;
  assign n16157 = P3_REG2_REG_4_ & ~n13941_1;
  assign n16158 = P3_REG2_REG_5_ & n16157;
  assign n16159 = ~P3_REG2_REG_5_ & ~n16157;
  assign n16160 = ~n14011_1 & ~n16159;
  assign n16161_1 = ~P3_REG2_REG_4_ & n13941_1;
  assign n16162 = ~P3_REG2_REG_5_ & n14011_1;
  assign n16163 = ~n16161_1 & ~n16162;
  assign n16164 = P3_REG2_REG_3_ & ~n13875;
  assign n16165 = ~P3_REG2_REG_3_ & n13875;
  assign n16166_1 = P3_REG2_REG_2_ & ~n13810;
  assign n16167 = ~n16165 & n16166_1;
  assign n16168 = ~P3_REG2_REG_2_ & n13810;
  assign n16169 = ~n16165 & ~n16168;
  assign n16170 = P3_REG2_REG_0_ & ~n13668;
  assign n16171_1 = ~P3_REG2_REG_1_ & n13754;
  assign n16172 = n16170 & ~n16171_1;
  assign n16173 = P3_REG2_REG_1_ & ~n13754;
  assign n16174 = ~n16172 & ~n16173;
  assign n16175 = n16169 & ~n16174;
  assign n16176_1 = ~n16164 & ~n16167;
  assign n16177 = ~n16175 & n16176_1;
  assign n16178 = n16163 & ~n16177;
  assign n16179 = ~n16158 & ~n16160;
  assign n16180 = ~n16178 & n16179;
  assign n16181_1 = n16156_1 & ~n16180;
  assign n16182 = ~n16151_1 & ~n16153;
  assign n16183 = ~n16181_1 & n16182;
  assign n16184 = n16144 & ~n16149;
  assign n16185 = ~n16183 & n16184;
  assign n16186_1 = ~n16148 & ~n16185;
  assign n16187 = n16133 & ~n16138;
  assign n16188 = ~n16186_1 & n16187;
  assign n16189 = ~n16137 & ~n16188;
  assign n16190 = ~n16127 & ~n16189;
  assign n16191_1 = ~n16126_1 & ~n16190;
  assign n16192 = ~n16125 & ~n16191_1;
  assign n16193 = ~n16124 & ~n16192;
  assign n16194 = n16123 & ~n16193;
  assign n16195 = ~n16118 & ~n16120;
  assign n16196_1 = ~n16194 & n16195;
  assign n16197 = P3_REG2_REG_18_ & ~n14863;
  assign n16198 = n16196_1 & ~n16197;
  assign n16199 = ~n16113 & ~n16116_1;
  assign n16200 = ~n16198 & n16199;
  assign n16201_1 = ~n16113 & ~n16196_1;
  assign n16202 = n16116_1 & ~n16197;
  assign n16203 = ~n16201_1 & n16202;
  assign n16204 = ~n16200 & ~n16203;
  assign n16205 = n16112 & n16204;
  assign n16206_1 = P3_REG3_REG_19_ & ~P3_STATE_REG;
  assign n16207 = ~n16205 & ~n16206_1;
  assign n16208 = P3_ADDR_REG_19_ & n16109;
  assign n16209 = n13664 & n16110;
  assign n16210 = ~n13593 & n16209;
  assign n16211_1 = n13661_1 & n16110;
  assign n16212 = ~P3_REG1_REG_18_ & n14863;
  assign n16213 = P3_REG1_REG_19_ & n13593;
  assign n16214 = ~P3_REG1_REG_19_ & ~n13593;
  assign n16215 = ~n16213 & ~n16214;
  assign n16216_1 = P3_REG1_REG_16_ & ~n14728;
  assign n16217 = P3_REG1_REG_17_ & n16216_1;
  assign n16218 = ~P3_REG1_REG_17_ & ~n16216_1;
  assign n16219 = ~n14795 & ~n16218;
  assign n16220 = ~P3_REG1_REG_16_ & n14728;
  assign n16221_1 = ~P3_REG1_REG_17_ & n14795;
  assign n16222 = ~n16220 & ~n16221_1;
  assign n16223 = P3_REG1_REG_15_ & ~n14667;
  assign n16224 = ~P3_REG1_REG_15_ & n14667;
  assign n16225 = P3_REG1_REG_14_ & ~n14606_1;
  assign n16226_1 = ~P3_REG1_REG_14_ & n14606_1;
  assign n16227 = ~P3_REG1_REG_13_ & n14540;
  assign n16228 = P3_REG1_REG_13_ & ~n14540;
  assign n16229 = P3_REG1_REG_12_ & ~n14474;
  assign n16230 = P3_REG1_REG_11_ & ~n14404;
  assign n16231_1 = ~P3_REG1_REG_12_ & n14474;
  assign n16232 = ~n16227 & ~n16231_1;
  assign n16233 = n16230 & n16232;
  assign n16234 = ~n16228 & ~n16229;
  assign n16235 = ~n16233 & n16234;
  assign n16236_1 = ~n16227 & ~n16235;
  assign n16237 = ~P3_REG1_REG_11_ & n14404;
  assign n16238 = ~P3_REG1_REG_10_ & n14352;
  assign n16239 = P3_REG1_REG_10_ & ~n14352;
  assign n16240 = P3_REG1_REG_9_ & ~n14273;
  assign n16241_1 = P3_REG1_REG_8_ & ~n14205;
  assign n16242 = ~P3_REG1_REG_9_ & n14273;
  assign n16243 = ~n16238 & ~n16242;
  assign n16244 = n16241_1 & n16243;
  assign n16245 = ~n16239 & ~n16240;
  assign n16246_1 = ~n16244 & n16245;
  assign n16247 = ~n16238 & ~n16246_1;
  assign n16248 = ~P3_REG1_REG_8_ & n14205;
  assign n16249 = P3_REG1_REG_6_ & ~n14063;
  assign n16250 = P3_REG1_REG_7_ & n16249;
  assign n16251_1 = ~P3_REG1_REG_7_ & ~n16249;
  assign n16252 = ~n14136_1 & ~n16251_1;
  assign n16253 = ~P3_REG1_REG_6_ & n14063;
  assign n16254 = ~P3_REG1_REG_7_ & n14136_1;
  assign n16255 = ~n16253 & ~n16254;
  assign n16256_1 = P3_REG1_REG_4_ & ~n13941_1;
  assign n16257 = P3_REG1_REG_5_ & n16256_1;
  assign n16258 = ~P3_REG1_REG_5_ & ~n16256_1;
  assign n16259 = ~n14011_1 & ~n16258;
  assign n16260 = ~P3_REG1_REG_4_ & n13941_1;
  assign n16261_1 = ~P3_REG1_REG_5_ & n14011_1;
  assign n16262 = ~n16260 & ~n16261_1;
  assign n16263 = P3_REG1_REG_3_ & ~n13875;
  assign n16264 = ~P3_REG1_REG_3_ & n13875;
  assign n16265 = P3_REG1_REG_2_ & ~n13810;
  assign n16266_1 = ~n16264 & n16265;
  assign n16267 = ~P3_REG1_REG_2_ & n13810;
  assign n16268 = ~n16264 & ~n16267;
  assign n16269 = P3_REG1_REG_0_ & ~n13668;
  assign n16270 = ~P3_REG1_REG_1_ & n13754;
  assign n16271_1 = n16269 & ~n16270;
  assign n16272 = P3_REG1_REG_1_ & ~n13754;
  assign n16273 = ~n16271_1 & ~n16272;
  assign n16274 = n16268 & ~n16273;
  assign n16275 = ~n16263 & ~n16266_1;
  assign n16276_1 = ~n16274 & n16275;
  assign n16277 = n16262 & ~n16276_1;
  assign n16278 = ~n16257 & ~n16259;
  assign n16279 = ~n16277 & n16278;
  assign n16280 = n16255 & ~n16279;
  assign n16281_1 = ~n16250 & ~n16252;
  assign n16282 = ~n16280 & n16281_1;
  assign n16283 = n16243 & ~n16248;
  assign n16284 = ~n16282 & n16283;
  assign n16285 = ~n16247 & ~n16284;
  assign n16286_1 = n16232 & ~n16237;
  assign n16287 = ~n16285 & n16286_1;
  assign n16288 = ~n16236_1 & ~n16287;
  assign n16289 = ~n16226_1 & ~n16288;
  assign n16290 = ~n16225 & ~n16289;
  assign n16291_1 = ~n16224 & ~n16290;
  assign n16292 = ~n16223 & ~n16291_1;
  assign n16293 = n16222 & ~n16292;
  assign n16294 = ~n16217 & ~n16219;
  assign n16295 = ~n16293 & n16294;
  assign n16296_1 = P3_REG1_REG_18_ & ~n14863;
  assign n16297 = n16295 & ~n16296_1;
  assign n16298 = ~n16212 & ~n16215;
  assign n16299 = ~n16297 & n16298;
  assign n16300 = ~n16212 & ~n16295;
  assign n16301_1 = n16215 & ~n16296_1;
  assign n16302 = ~n16300 & n16301_1;
  assign n16303 = ~n16299 & ~n16302;
  assign n16304 = n16211_1 & n16303;
  assign n16305 = ~n16208 & ~n16210;
  assign n16306_1 = ~n16304 & n16305;
  assign n16307 = n13525 & ~n16109;
  assign n16308 = ~n13716_1 & ~n13725;
  assign n16309 = ~n13733 & n16308;
  assign n16310 = ~n13721_1 & ~n15720;
  assign n16311_1 = ~n13719 & n16310;
  assign n16312 = ~n13727 & ~n13730;
  assign n16313 = ~n15697 & n16312;
  assign n16314 = n16309 & n16311_1;
  assign n16315 = n16313 & n16314;
  assign n16316_1 = n15708 & n16315;
  assign n16317 = ~n15698 & n16316_1;
  assign n16318 = n13664 & ~n16317;
  assign n16319 = ~n13593 & n16318;
  assign n16320 = n16111_1 & ~n16317;
  assign n16321_1 = n16204 & n16320;
  assign n16322 = n13661_1 & ~n16317;
  assign n16323 = n16303 & n16322;
  assign n16324 = ~n16319 & ~n16321_1;
  assign n16325 = ~n16323 & n16324;
  assign n16326_1 = n16307 & ~n16325;
  assign n16327 = n16207 & n16306_1;
  assign n1601 = n16326_1 | ~n16327;
  assign n16329 = P3_REG2_REG_18_ & n14863;
  assign n16330 = ~P3_REG2_REG_18_ & ~n14863;
  assign n16331_1 = ~n16329 & ~n16330;
  assign n16332 = n16196_1 & ~n16331_1;
  assign n16333 = ~n16196_1 & n16331_1;
  assign n16334 = ~n16332 & ~n16333;
  assign n16335 = n16112 & ~n16334;
  assign n16336_1 = P3_REG3_REG_18_ & ~P3_STATE_REG;
  assign n16337 = ~n16335 & ~n16336_1;
  assign n16338 = P3_ADDR_REG_18_ & n16109;
  assign n16339 = ~n14863 & n16209;
  assign n16340 = P3_REG1_REG_18_ & n14863;
  assign n16341_1 = ~P3_REG1_REG_18_ & ~n14863;
  assign n16342 = ~n16340 & ~n16341_1;
  assign n16343 = n16295 & ~n16342;
  assign n16344 = ~n16295 & n16342;
  assign n16345 = ~n16343 & ~n16344;
  assign n16346_1 = n16211_1 & ~n16345;
  assign n16347 = ~n16338 & ~n16339;
  assign n16348 = ~n16346_1 & n16347;
  assign n16349 = ~n14863 & n16318;
  assign n16350 = n16320 & ~n16334;
  assign n16351_1 = n16322 & ~n16345;
  assign n16352 = ~n16349 & ~n16350;
  assign n16353 = ~n16351_1 & n16352;
  assign n16354 = n16307 & ~n16353;
  assign n16355 = n16337 & n16348;
  assign n1606 = n16354 | ~n16355;
  assign n16357 = P3_REG2_REG_17_ & ~n14795;
  assign n16358 = ~n16117 & n16193;
  assign n16359 = n16123 & ~n16357;
  assign n16360 = ~n16358 & n16359;
  assign n16361_1 = P3_REG2_REG_17_ & n14795;
  assign n16362 = ~P3_REG2_REG_17_ & ~n14795;
  assign n16363 = ~n16121_1 & ~n16193;
  assign n16364 = ~n16361_1 & ~n16362;
  assign n16365 = ~n16117 & n16364;
  assign n16366_1 = ~n16363 & n16365;
  assign n16367 = ~n16360 & ~n16366_1;
  assign n16368 = n16112 & n16367;
  assign n16369 = P3_REG3_REG_17_ & ~P3_STATE_REG;
  assign n16370 = ~n16368 & ~n16369;
  assign n16371_1 = P3_ADDR_REG_17_ & n16109;
  assign n16372 = ~n14795 & n16209;
  assign n16373 = P3_REG1_REG_17_ & ~n14795;
  assign n16374 = ~n16216_1 & n16292;
  assign n16375 = n16222 & ~n16373;
  assign n16376_1 = ~n16374 & n16375;
  assign n16377 = P3_REG1_REG_17_ & n14795;
  assign n16378 = ~P3_REG1_REG_17_ & ~n14795;
  assign n16379 = ~n16220 & ~n16292;
  assign n16380 = ~n16377 & ~n16378;
  assign n16381_1 = ~n16216_1 & n16380;
  assign n16382 = ~n16379 & n16381_1;
  assign n16383 = ~n16376_1 & ~n16382;
  assign n16384 = n16211_1 & n16383;
  assign n16385 = ~n16371_1 & ~n16372;
  assign n16386_1 = ~n16384 & n16385;
  assign n16387 = ~n14795 & n16318;
  assign n16388 = n16320 & n16367;
  assign n16389 = n16322 & n16383;
  assign n16390 = ~n16387 & ~n16388;
  assign n16391_1 = ~n16389 & n16390;
  assign n16392 = n16307 & ~n16391_1;
  assign n16393 = n16370 & n16386_1;
  assign n1611 = n16392 | ~n16393;
  assign n16395 = P3_REG2_REG_16_ & n14728;
  assign n16396_1 = ~P3_REG2_REG_16_ & ~n14728;
  assign n16397 = ~n16395 & ~n16396_1;
  assign n16398 = n16193 & ~n16397;
  assign n16399 = ~n16117 & ~n16121_1;
  assign n16400 = ~n16193 & ~n16399;
  assign n16401_1 = ~n16398 & ~n16400;
  assign n16402 = n16112 & ~n16401_1;
  assign n16403 = P3_REG3_REG_16_ & ~P3_STATE_REG;
  assign n16404 = ~n16402 & ~n16403;
  assign n16405 = P3_ADDR_REG_16_ & n16109;
  assign n16406_1 = ~n14728 & n16209;
  assign n16407 = P3_REG1_REG_16_ & n14728;
  assign n16408 = ~P3_REG1_REG_16_ & ~n14728;
  assign n16409 = ~n16407 & ~n16408;
  assign n16410 = n16292 & ~n16409;
  assign n16411_1 = ~n16216_1 & ~n16220;
  assign n16412 = ~n16292 & ~n16411_1;
  assign n16413 = ~n16410 & ~n16412;
  assign n16414 = n16211_1 & ~n16413;
  assign n16415 = ~n16405 & ~n16406_1;
  assign n16416_1 = ~n16414 & n16415;
  assign n16417 = ~n14728 & n16318;
  assign n16418 = n16320 & ~n16401_1;
  assign n16419 = n16322 & ~n16413;
  assign n16420 = ~n16417 & ~n16418;
  assign n16421_1 = ~n16419 & n16420;
  assign n16422 = n16307 & ~n16421_1;
  assign n16423 = n16404 & n16416_1;
  assign n1616 = n16422 | ~n16423;
  assign n16425 = P3_REG2_REG_15_ & n14667;
  assign n16426_1 = ~P3_REG2_REG_15_ & ~n14667;
  assign n16427 = ~n16425 & ~n16426_1;
  assign n16428 = n16191_1 & ~n16427;
  assign n16429 = ~n16191_1 & n16427;
  assign n16430 = ~n16428 & ~n16429;
  assign n16431_1 = n16112 & ~n16430;
  assign n16432 = P3_REG3_REG_15_ & ~P3_STATE_REG;
  assign n16433 = ~n16431_1 & ~n16432;
  assign n16434 = P3_ADDR_REG_15_ & n16109;
  assign n16435 = ~n14667 & n16209;
  assign n16436_1 = P3_REG1_REG_15_ & n14667;
  assign n16437 = ~P3_REG1_REG_15_ & ~n14667;
  assign n16438 = ~n16436_1 & ~n16437;
  assign n16439 = n16290 & ~n16438;
  assign n16440 = ~n16290 & n16438;
  assign n16441_1 = ~n16439 & ~n16440;
  assign n16442 = n16211_1 & ~n16441_1;
  assign n16443 = ~n16434 & ~n16435;
  assign n16444 = ~n16442 & n16443;
  assign n16445 = ~n14667 & n16318;
  assign n16446_1 = n16320 & ~n16430;
  assign n16447 = n16322 & ~n16441_1;
  assign n16448 = ~n16445 & ~n16446_1;
  assign n16449 = ~n16447 & n16448;
  assign n16450 = n16307 & ~n16449;
  assign n16451_1 = n16433 & n16444;
  assign n1621 = n16450 | ~n16451_1;
  assign n16453 = P3_REG2_REG_14_ & n14606_1;
  assign n16454 = ~P3_REG2_REG_14_ & ~n14606_1;
  assign n16455 = ~n16453 & ~n16454;
  assign n16456_1 = n16189 & ~n16455;
  assign n16457 = ~n16189 & n16455;
  assign n16458 = ~n16456_1 & ~n16457;
  assign n16459 = n16112 & ~n16458;
  assign n16460 = P3_REG3_REG_14_ & ~P3_STATE_REG;
  assign n16461_1 = ~n16459 & ~n16460;
  assign n16462 = P3_ADDR_REG_14_ & n16109;
  assign n16463 = ~n14606_1 & n16209;
  assign n16464 = P3_REG1_REG_14_ & n14606_1;
  assign n16465 = ~P3_REG1_REG_14_ & ~n14606_1;
  assign n16466_1 = ~n16464 & ~n16465;
  assign n16467 = n16288 & ~n16466_1;
  assign n16468 = ~n16288 & n16466_1;
  assign n16469 = ~n16467 & ~n16468;
  assign n16470 = n16211_1 & ~n16469;
  assign n16471_1 = ~n16462 & ~n16463;
  assign n16472 = ~n16470 & n16471_1;
  assign n16473 = ~n14606_1 & n16318;
  assign n16474 = n16320 & ~n16458;
  assign n16475 = n16322 & ~n16469;
  assign n16476_1 = ~n16473 & ~n16474;
  assign n16477 = ~n16475 & n16476_1;
  assign n16478 = n16307 & ~n16477;
  assign n16479 = n16461_1 & n16472;
  assign n1626 = n16478 | ~n16479;
  assign n16481_1 = ~n16138 & ~n16186_1;
  assign n16482 = ~n16131_1 & ~n16481_1;
  assign n16483 = ~n16130 & n16482;
  assign n16484 = ~n16129 & n16133;
  assign n16485 = ~n16483 & n16484;
  assign n16486_1 = P3_REG2_REG_13_ & n14540;
  assign n16487 = ~P3_REG2_REG_13_ & ~n14540;
  assign n16488 = ~n16132 & ~n16482;
  assign n16489 = ~n16486_1 & ~n16487;
  assign n16490 = ~n16130 & n16489;
  assign n16491_1 = ~n16488 & n16490;
  assign n16492 = ~n16485 & ~n16491_1;
  assign n16493 = n16112 & n16492;
  assign n16494 = P3_REG3_REG_13_ & ~P3_STATE_REG;
  assign n16495 = ~n16493 & ~n16494;
  assign n16496_1 = P3_ADDR_REG_13_ & n16109;
  assign n16497 = ~n14540 & n16209;
  assign n16498 = ~n16237 & ~n16285;
  assign n16499 = ~n16230 & ~n16498;
  assign n16500 = ~n16229 & n16499;
  assign n16501_1 = ~n16228 & n16232;
  assign n16502 = ~n16500 & n16501_1;
  assign n16503 = P3_REG1_REG_13_ & n14540;
  assign n16504 = ~P3_REG1_REG_13_ & ~n14540;
  assign n16505 = ~n16231_1 & ~n16499;
  assign n16506_1 = ~n16503 & ~n16504;
  assign n16507 = ~n16229 & n16506_1;
  assign n16508 = ~n16505 & n16507;
  assign n16509 = ~n16502 & ~n16508;
  assign n16510 = n16211_1 & n16509;
  assign n16511_1 = ~n16496_1 & ~n16497;
  assign n16512 = ~n16510 & n16511_1;
  assign n16513 = ~n14540 & n16318;
  assign n16514 = n16320 & n16492;
  assign n16515 = n16322 & n16509;
  assign n16516_1 = ~n16513 & ~n16514;
  assign n16517 = ~n16515 & n16516_1;
  assign n16518 = n16307 & ~n16517;
  assign n16519 = n16495 & n16512;
  assign n1631 = n16518 | ~n16519;
  assign n16521_1 = P3_REG2_REG_12_ & n14474;
  assign n16522 = ~P3_REG2_REG_12_ & ~n14474;
  assign n16523 = ~n16521_1 & ~n16522;
  assign n16524 = n16482 & ~n16523;
  assign n16525 = ~n16130 & ~n16132;
  assign n16526_1 = ~n16482 & ~n16525;
  assign n16527 = ~n16524 & ~n16526_1;
  assign n16528 = n16112 & ~n16527;
  assign n16529 = P3_REG3_REG_12_ & ~P3_STATE_REG;
  assign n16530 = ~n16528 & ~n16529;
  assign n16531_1 = P3_ADDR_REG_12_ & n16109;
  assign n16532 = ~n14474 & n16209;
  assign n16533 = P3_REG1_REG_12_ & n14474;
  assign n16534 = ~P3_REG1_REG_12_ & ~n14474;
  assign n16535 = ~n16533 & ~n16534;
  assign n16536_1 = n16499 & ~n16535;
  assign n16537 = ~n16229 & ~n16231_1;
  assign n16538 = ~n16499 & ~n16537;
  assign n16539 = ~n16536_1 & ~n16538;
  assign n16540 = n16211_1 & ~n16539;
  assign n16541_1 = ~n16531_1 & ~n16532;
  assign n16542 = ~n16540 & n16541_1;
  assign n16543 = ~n14474 & n16318;
  assign n16544 = n16320 & ~n16527;
  assign n16545 = n16322 & ~n16539;
  assign n16546_1 = ~n16543 & ~n16544;
  assign n16547 = ~n16545 & n16546_1;
  assign n16548 = n16307 & ~n16547;
  assign n16549 = n16530 & n16542;
  assign n1636 = n16548 | ~n16549;
  assign n16551_1 = P3_REG2_REG_11_ & n14404;
  assign n16552 = ~P3_REG2_REG_11_ & ~n14404;
  assign n16553 = ~n16551_1 & ~n16552;
  assign n16554 = n16186_1 & ~n16553;
  assign n16555 = ~n16131_1 & ~n16138;
  assign n16556_1 = ~n16186_1 & ~n16555;
  assign n16557 = ~n16554 & ~n16556_1;
  assign n16558 = n16112 & ~n16557;
  assign n16559 = P3_REG3_REG_11_ & ~P3_STATE_REG;
  assign n16560 = ~n16558 & ~n16559;
  assign n16561_1 = P3_ADDR_REG_11_ & n16109;
  assign n16562 = ~n14404 & n16209;
  assign n16563 = P3_REG1_REG_11_ & n14404;
  assign n16564 = ~P3_REG1_REG_11_ & ~n14404;
  assign n16565 = ~n16563 & ~n16564;
  assign n16566_1 = n16285 & ~n16565;
  assign n16567 = ~n16230 & ~n16237;
  assign n16568 = ~n16285 & ~n16567;
  assign n16569 = ~n16566_1 & ~n16568;
  assign n16570 = n16211_1 & ~n16569;
  assign n16571_1 = ~n16561_1 & ~n16562;
  assign n16572 = ~n16570 & n16571_1;
  assign n16573 = ~n14404 & n16318;
  assign n16574 = n16320 & ~n16557;
  assign n16575 = n16322 & ~n16569;
  assign n16576_1 = ~n16573 & ~n16574;
  assign n16577 = ~n16575 & n16576_1;
  assign n16578 = n16307 & ~n16577;
  assign n16579 = n16560 & n16572;
  assign n1641 = n16578 | ~n16579;
  assign n16581_1 = ~n16149 & ~n16183;
  assign n16582 = ~n16142 & ~n16581_1;
  assign n16583 = ~n16141_1 & n16582;
  assign n16584 = ~n16140 & n16144;
  assign n16585 = ~n16583 & n16584;
  assign n16586_1 = P3_REG2_REG_10_ & n14352;
  assign n16587 = ~P3_REG2_REG_10_ & ~n14352;
  assign n16588 = ~n16143 & ~n16582;
  assign n16589 = ~n16586_1 & ~n16587;
  assign n16590 = ~n16141_1 & n16589;
  assign n16591_1 = ~n16588 & n16590;
  assign n16592 = ~n16585 & ~n16591_1;
  assign n16593 = n16112 & n16592;
  assign n16594 = P3_REG3_REG_10_ & ~P3_STATE_REG;
  assign n16595 = ~n16593 & ~n16594;
  assign n16596_1 = P3_ADDR_REG_10_ & n16109;
  assign n16597 = ~n14352 & n16209;
  assign n16598 = ~n16248 & ~n16282;
  assign n16599 = ~n16241_1 & ~n16598;
  assign n16600 = ~n16240 & n16599;
  assign n16601_1 = ~n16239 & n16243;
  assign n16602 = ~n16600 & n16601_1;
  assign n16603 = P3_REG1_REG_10_ & n14352;
  assign n16604 = ~P3_REG1_REG_10_ & ~n14352;
  assign n16605 = ~n16242 & ~n16599;
  assign n16606_1 = ~n16603 & ~n16604;
  assign n16607 = ~n16240 & n16606_1;
  assign n16608 = ~n16605 & n16607;
  assign n16609 = ~n16602 & ~n16608;
  assign n16610 = n16211_1 & n16609;
  assign n16611_1 = ~n16596_1 & ~n16597;
  assign n16612 = ~n16610 & n16611_1;
  assign n16613 = ~n14352 & n16318;
  assign n16614 = n16320 & n16592;
  assign n16615 = n16322 & n16609;
  assign n16616_1 = ~n16613 & ~n16614;
  assign n16617 = ~n16615 & n16616_1;
  assign n16618 = n16307 & ~n16617;
  assign n16619 = n16595 & n16612;
  assign n1646 = n16618 | ~n16619;
  assign n16621_1 = P3_REG2_REG_9_ & n14273;
  assign n16622 = ~P3_REG2_REG_9_ & ~n14273;
  assign n16623 = ~n16621_1 & ~n16622;
  assign n16624 = n16582 & ~n16623;
  assign n16625 = ~n16141_1 & ~n16143;
  assign n16626_1 = ~n16582 & ~n16625;
  assign n16627 = ~n16624 & ~n16626_1;
  assign n16628 = n16112 & ~n16627;
  assign n16629 = P3_REG3_REG_9_ & ~P3_STATE_REG;
  assign n16630 = ~n16628 & ~n16629;
  assign n16631_1 = P3_ADDR_REG_9_ & n16109;
  assign n16632 = ~n14273 & n16209;
  assign n16633 = P3_REG1_REG_9_ & n14273;
  assign n16634 = ~P3_REG1_REG_9_ & ~n14273;
  assign n16635 = ~n16633 & ~n16634;
  assign n16636_1 = n16599 & ~n16635;
  assign n16637 = ~n16240 & ~n16242;
  assign n16638 = ~n16599 & ~n16637;
  assign n16639 = ~n16636_1 & ~n16638;
  assign n16640 = n16211_1 & ~n16639;
  assign n16641_1 = ~n16631_1 & ~n16632;
  assign n16642 = ~n16640 & n16641_1;
  assign n16643 = ~n14273 & n16318;
  assign n16644 = n16320 & ~n16627;
  assign n16645 = n16322 & ~n16639;
  assign n16646_1 = ~n16643 & ~n16644;
  assign n16647 = ~n16645 & n16646_1;
  assign n16648 = n16307 & ~n16647;
  assign n16649 = n16630 & n16642;
  assign n1651 = n16648 | ~n16649;
  assign n16651_1 = P3_REG2_REG_8_ & n14205;
  assign n16652 = ~P3_REG2_REG_8_ & ~n14205;
  assign n16653 = ~n16651_1 & ~n16652;
  assign n16654 = n16183 & ~n16653;
  assign n16655 = ~n16142 & ~n16149;
  assign n16656_1 = ~n16183 & ~n16655;
  assign n16657 = ~n16654 & ~n16656_1;
  assign n16658 = n16112 & ~n16657;
  assign n16659 = P3_REG3_REG_8_ & ~P3_STATE_REG;
  assign n16660 = ~n16658 & ~n16659;
  assign n16661_1 = P3_ADDR_REG_8_ & n16109;
  assign n16662 = ~n14205 & n16209;
  assign n16663 = P3_REG1_REG_8_ & n14205;
  assign n16664 = ~P3_REG1_REG_8_ & ~n14205;
  assign n16665 = ~n16663 & ~n16664;
  assign n16666_1 = n16282 & ~n16665;
  assign n16667 = ~n16241_1 & ~n16248;
  assign n16668 = ~n16282 & ~n16667;
  assign n16669 = ~n16666_1 & ~n16668;
  assign n16670 = n16211_1 & ~n16669;
  assign n16671_1 = ~n16661_1 & ~n16662;
  assign n16672 = ~n16670 & n16671_1;
  assign n16673 = ~n14205 & n16318;
  assign n16674 = n16320 & ~n16657;
  assign n16675 = n16322 & ~n16669;
  assign n16676_1 = ~n16673 & ~n16674;
  assign n16677 = ~n16675 & n16676_1;
  assign n16678 = n16307 & ~n16677;
  assign n16679 = n16660 & n16672;
  assign n1656 = n16678 | ~n16679;
  assign n16681_1 = P3_REG2_REG_7_ & ~n14136_1;
  assign n16682 = ~n16150 & n16180;
  assign n16683 = n16156_1 & ~n16681_1;
  assign n16684 = ~n16682 & n16683;
  assign n16685 = P3_REG2_REG_7_ & n14136_1;
  assign n16686_1 = ~P3_REG2_REG_7_ & ~n14136_1;
  assign n16687 = ~n16154 & ~n16180;
  assign n16688 = ~n16685 & ~n16686_1;
  assign n16689 = ~n16150 & n16688;
  assign n16690 = ~n16687 & n16689;
  assign n16691_1 = ~n16684 & ~n16690;
  assign n16692 = n16112 & n16691_1;
  assign n16693 = P3_REG3_REG_7_ & ~P3_STATE_REG;
  assign n16694 = ~n16692 & ~n16693;
  assign n16695 = P3_REG1_REG_7_ & ~n14136_1;
  assign n16696_1 = ~n16249 & n16279;
  assign n16697 = n16255 & ~n16695;
  assign n16698 = ~n16696_1 & n16697;
  assign n16699 = P3_REG1_REG_7_ & n14136_1;
  assign n16700 = ~P3_REG1_REG_7_ & ~n14136_1;
  assign n16701_1 = ~n16253 & ~n16279;
  assign n16702 = ~n16699 & ~n16700;
  assign n16703 = ~n16249 & n16702;
  assign n16704 = ~n16701_1 & n16703;
  assign n16705 = ~n16698 & ~n16704;
  assign n16706_1 = n16211_1 & n16705;
  assign n16707 = ~n14136_1 & n16209;
  assign n16708 = P3_ADDR_REG_7_ & n16109;
  assign n16709 = ~n16706_1 & ~n16707;
  assign n16710 = ~n16708 & n16709;
  assign n16711_1 = ~n14136_1 & n16318;
  assign n16712 = n16320 & n16691_1;
  assign n16713 = n16322 & n16705;
  assign n16714 = ~n16711_1 & ~n16712;
  assign n16715 = ~n16713 & n16714;
  assign n16716_1 = n16307 & ~n16715;
  assign n16717 = n16694 & n16710;
  assign n1661 = n16716_1 | ~n16717;
  assign n16719 = P3_REG1_REG_6_ & n14063;
  assign n16720 = ~P3_REG1_REG_6_ & ~n14063;
  assign n16721 = ~n16719 & ~n16720;
  assign n16722 = n16279 & ~n16721;
  assign n16723 = ~n16249 & ~n16253;
  assign n16724 = ~n16279 & ~n16723;
  assign n16725 = ~n16722 & ~n16724;
  assign n16726 = n16211_1 & ~n16725;
  assign n16727 = ~n14063 & n16209;
  assign n16728 = P3_ADDR_REG_6_ & n16109;
  assign n16729 = ~n16726 & ~n16727;
  assign n16730 = ~n16728 & n16729;
  assign n16731 = P3_REG2_REG_6_ & n14063;
  assign n16732 = ~P3_REG2_REG_6_ & ~n14063;
  assign n16733 = ~n16731 & ~n16732;
  assign n16734 = n16180 & ~n16733;
  assign n16735 = ~n16150 & ~n16154;
  assign n16736 = ~n16180 & ~n16735;
  assign n16737 = ~n16734 & ~n16736;
  assign n16738 = n16112 & ~n16737;
  assign n16739 = P3_REG3_REG_6_ & ~P3_STATE_REG;
  assign n16740 = ~n14063 & n16318;
  assign n16741 = n16320 & ~n16737;
  assign n16742 = n16322 & ~n16725;
  assign n16743 = ~n16740 & ~n16741;
  assign n16744 = ~n16742 & n16743;
  assign n16745 = n16307 & ~n16744;
  assign n16746 = ~n16738 & ~n16739;
  assign n16747 = ~n16745 & n16746;
  assign n1666 = ~n16730 | ~n16747;
  assign n16749 = P3_REG1_REG_5_ & ~n14011_1;
  assign n16750 = n16268 & n16271_1;
  assign n16751 = ~n16267 & n16272;
  assign n16752 = ~n16265 & ~n16751;
  assign n16753 = ~n16264 & ~n16752;
  assign n16754 = ~n16263 & ~n16750;
  assign n16755 = ~n16753 & n16754;
  assign n16756 = ~n16256_1 & n16755;
  assign n16757 = n16262 & ~n16749;
  assign n16758 = ~n16756 & n16757;
  assign n16759 = P3_REG1_REG_5_ & n14011_1;
  assign n16760 = ~P3_REG1_REG_5_ & ~n14011_1;
  assign n16761 = ~n16260 & ~n16755;
  assign n16762 = ~n16759 & ~n16760;
  assign n16763 = ~n16256_1 & n16762;
  assign n16764 = ~n16761 & n16763;
  assign n16765 = ~n16758 & ~n16764;
  assign n16766 = n16211_1 & n16765;
  assign n16767 = ~n14011_1 & n16209;
  assign n16768 = P3_ADDR_REG_5_ & n16109;
  assign n16769 = ~n16766 & ~n16767;
  assign n16770 = ~n16768 & n16769;
  assign n16771 = P3_REG2_REG_5_ & ~n14011_1;
  assign n16772 = n16169 & n16172;
  assign n16773 = ~n16168 & n16173;
  assign n16774 = ~n16166_1 & ~n16773;
  assign n16775 = ~n16165 & ~n16774;
  assign n16776 = ~n16164 & ~n16772;
  assign n16777 = ~n16775 & n16776;
  assign n16778 = ~n16157 & n16777;
  assign n16779 = n16163 & ~n16771;
  assign n16780 = ~n16778 & n16779;
  assign n16781 = P3_REG2_REG_5_ & n14011_1;
  assign n16782 = ~P3_REG2_REG_5_ & ~n14011_1;
  assign n16783 = ~n16161_1 & ~n16777;
  assign n16784 = ~n16781 & ~n16782;
  assign n16785 = ~n16157 & n16784;
  assign n16786 = ~n16783 & n16785;
  assign n16787 = ~n16780 & ~n16786;
  assign n16788 = n16112 & n16787;
  assign n16789 = P3_REG3_REG_5_ & ~P3_STATE_REG;
  assign n16790 = ~n14011_1 & n16318;
  assign n16791 = n16320 & n16787;
  assign n16792 = n16322 & n16765;
  assign n16793 = ~n16790 & ~n16791;
  assign n16794 = ~n16792 & n16793;
  assign n16795 = n16307 & ~n16794;
  assign n16796 = ~n16788 & ~n16789;
  assign n16797 = ~n16795 & n16796;
  assign n1671 = ~n16770 | ~n16797;
  assign n16799 = P3_REG1_REG_4_ & n13941_1;
  assign n16800 = ~P3_REG1_REG_4_ & ~n13941_1;
  assign n16801 = ~n16799 & ~n16800;
  assign n16802 = n16755 & ~n16801;
  assign n16803 = ~n16256_1 & ~n16260;
  assign n16804 = ~n16755 & ~n16803;
  assign n16805 = ~n16802 & ~n16804;
  assign n16806 = n16211_1 & ~n16805;
  assign n16807 = ~n13941_1 & n16209;
  assign n16808 = P3_ADDR_REG_4_ & n16109;
  assign n16809 = ~n16806 & ~n16807;
  assign n16810 = ~n16808 & n16809;
  assign n16811 = P3_REG3_REG_4_ & ~P3_STATE_REG;
  assign n16812 = P3_REG2_REG_4_ & n13941_1;
  assign n16813 = ~P3_REG2_REG_4_ & ~n13941_1;
  assign n16814 = ~n16812 & ~n16813;
  assign n16815 = n16777 & ~n16814;
  assign n16816 = ~n16157 & ~n16161_1;
  assign n16817 = ~n16777 & ~n16816;
  assign n16818 = ~n16815 & ~n16817;
  assign n16819 = n16112 & ~n16818;
  assign n16820 = ~n13941_1 & n16318;
  assign n16821 = n16320 & ~n16818;
  assign n16822 = n16322 & ~n16805;
  assign n16823 = ~n16820 & ~n16821;
  assign n16824 = ~n16822 & n16823;
  assign n16825 = n16307 & ~n16824;
  assign n2021 = P3_STATE_REG & n16104;
  assign n16827 = P3_REG2_REG_0_ & n16111_1;
  assign n16828 = n13668 & n16827;
  assign n16829 = ~P3_REG2_REG_0_ & ~n13661_1;
  assign n16830 = ~n13664 & ~n16829;
  assign n16831 = ~n13668 & ~n16830;
  assign n16832 = n13587 & ~n13593;
  assign n16833 = ~n13584 & ~n13587;
  assign n16834 = ~n16832 & ~n16833;
  assign n16835 = ~n13523 & n13672;
  assign n16836 = n16834 & ~n16835;
  assign n16837 = ~n13523 & ~n16836;
  assign n16838 = n13523 & ~n13668;
  assign n16839 = ~n13523 & ~n16310;
  assign n16840 = ~n13671_1 & n16839;
  assign n16841 = ~n16838 & ~n16840;
  assign n16842 = ~n13673 & ~n13716_1;
  assign n16843 = ~n13725 & n16842;
  assign n16844 = ~n13523 & ~n16843;
  assign n16845 = ~n13523 & n16832;
  assign n16846 = ~n16844 & ~n16845;
  assign n16847 = ~n13707 & ~n16846;
  assign n16848 = n16841 & ~n16847;
  assign n16849 = n16837 & n16848;
  assign n16850 = ~n16837 & ~n16848;
  assign n16851 = ~n16849 & ~n16850;
  assign n16852 = ~n13707 & n16839;
  assign n16853 = P3_REG1_REG_0_ & n13523;
  assign n16854 = ~n16852 & ~n16853;
  assign n16855 = ~n16835 & n16846;
  assign n16856 = ~n13671_1 & ~n16855;
  assign n16857 = n16854 & ~n16856;
  assign n16858 = ~n16837 & ~n16857;
  assign n16859 = n16837 & n16857;
  assign n16860 = ~n16858 & ~n16859;
  assign n16861 = ~n16851 & n16860;
  assign n16862 = n16851 & ~n16860;
  assign n16863 = ~n16861 & ~n16862;
  assign n16864 = n13661_1 & ~n13664;
  assign n16865 = ~n16863 & n16864;
  assign n16866 = ~n16828 & ~n16831;
  assign n16867 = ~n16865 & n16866;
  assign n16868 = n2021 & ~n16867;
  assign n16869 = ~n16825 & ~n16868;
  assign n16870 = ~n16811 & ~n16819;
  assign n16871 = n16869 & n16870;
  assign n1676 = ~n16810 | ~n16871;
  assign n16873 = ~n16267 & n16271_1;
  assign n16874 = n16752 & ~n16873;
  assign n16875 = P3_REG1_REG_3_ & n13875;
  assign n16876 = ~P3_REG1_REG_3_ & ~n13875;
  assign n16877 = ~n16875 & ~n16876;
  assign n16878 = n16874 & ~n16877;
  assign n16879 = ~n16263 & ~n16264;
  assign n16880 = ~n16874 & ~n16879;
  assign n16881 = ~n16878 & ~n16880;
  assign n16882 = n16211_1 & ~n16881;
  assign n16883 = ~n13875 & n16209;
  assign n16884 = P3_ADDR_REG_3_ & n16109;
  assign n16885 = ~n16882 & ~n16883;
  assign n16886 = ~n16884 & n16885;
  assign n16887 = ~n16168 & n16172;
  assign n16888 = n16774 & ~n16887;
  assign n16889 = P3_REG2_REG_3_ & n13875;
  assign n16890 = ~P3_REG2_REG_3_ & ~n13875;
  assign n16891 = ~n16889 & ~n16890;
  assign n16892 = n16888 & ~n16891;
  assign n16893 = ~n16164 & ~n16165;
  assign n16894 = ~n16888 & ~n16893;
  assign n16895 = ~n16892 & ~n16894;
  assign n16896 = n16112 & ~n16895;
  assign n16897 = P3_REG3_REG_3_ & ~P3_STATE_REG;
  assign n16898 = ~n13875 & n16318;
  assign n16899 = n16320 & ~n16895;
  assign n16900 = n16322 & ~n16881;
  assign n16901 = ~n16898 & ~n16899;
  assign n16902 = ~n16900 & n16901;
  assign n16903 = n16307 & ~n16902;
  assign n16904 = ~n16896 & ~n16897;
  assign n16905 = ~n16903 & n16904;
  assign n1681 = ~n16886 | ~n16905;
  assign n16907 = ~n16265 & ~n16267;
  assign n16908 = ~n16273 & n16907;
  assign n16909 = P3_REG1_REG_2_ & n13810;
  assign n16910 = ~P3_REG1_REG_2_ & ~n13810;
  assign n16911 = ~n16909 & ~n16910;
  assign n16912 = ~n16272 & n16911;
  assign n16913 = ~n16271_1 & n16912;
  assign n16914 = ~n16908 & ~n16913;
  assign n16915 = n16211_1 & n16914;
  assign n16916 = ~n13810 & n16209;
  assign n16917 = P3_ADDR_REG_2_ & n16109;
  assign n16918 = ~n16915 & ~n16916;
  assign n16919 = ~n16917 & n16918;
  assign n16920 = P3_REG3_REG_2_ & ~P3_STATE_REG;
  assign n16921 = ~n16166_1 & ~n16168;
  assign n16922 = ~n16174 & n16921;
  assign n16923 = P3_REG2_REG_2_ & n13810;
  assign n16924 = ~P3_REG2_REG_2_ & ~n13810;
  assign n16925 = n16174 & ~n16923;
  assign n16926 = ~n16924 & n16925;
  assign n16927 = ~n16922 & ~n16926;
  assign n16928 = n16112 & n16927;
  assign n16929 = ~n13810 & n16318;
  assign n16930 = n16320 & n16927;
  assign n16931 = n16322 & n16914;
  assign n16932 = ~n16929 & ~n16930;
  assign n16933 = ~n16931 & n16932;
  assign n16934 = n16307 & ~n16933;
  assign n16935 = ~n16868 & ~n16934;
  assign n16936 = ~n16920 & ~n16928;
  assign n16937 = n16935 & n16936;
  assign n1686 = ~n16919 | ~n16937;
  assign n16939 = ~n16270 & ~n16272;
  assign n16940 = ~n16269 & n16939;
  assign n16941 = n16269 & ~n16939;
  assign n16942 = ~n16940 & ~n16941;
  assign n16943 = n16211_1 & ~n16942;
  assign n16944 = ~n13754 & n16209;
  assign n16945 = P3_ADDR_REG_1_ & n16109;
  assign n16946 = ~n16943 & ~n16944;
  assign n16947 = ~n16945 & n16946;
  assign n16948 = ~n16171_1 & ~n16173;
  assign n16949 = ~n16170 & n16948;
  assign n16950 = n16170 & ~n16948;
  assign n16951 = ~n16949 & ~n16950;
  assign n16952 = n16112 & ~n16951;
  assign n16953 = P3_REG3_REG_1_ & ~P3_STATE_REG;
  assign n16954 = ~n13754 & n16318;
  assign n16955 = n16320 & ~n16951;
  assign n16956 = n16322 & ~n16942;
  assign n16957 = ~n16954 & ~n16955;
  assign n16958 = ~n16956 & n16957;
  assign n16959 = n16307 & ~n16958;
  assign n16960 = ~n16952 & ~n16953;
  assign n16961 = ~n16959 & n16960;
  assign n1691 = ~n16947 | ~n16961;
  assign n16963 = P3_REG1_REG_0_ & n13668;
  assign n16964 = ~P3_REG1_REG_0_ & ~n13668;
  assign n16965 = ~n16963 & ~n16964;
  assign n16966 = n16211_1 & ~n16965;
  assign n16967 = ~n13668 & n16209;
  assign n16968 = P3_ADDR_REG_0_ & n16109;
  assign n16969 = ~n16966 & ~n16967;
  assign n16970 = ~n16968 & n16969;
  assign n16971 = P3_REG2_REG_0_ & n13668;
  assign n16972 = ~P3_REG2_REG_0_ & ~n13668;
  assign n16973 = ~n16971 & ~n16972;
  assign n16974 = n16112 & ~n16973;
  assign n16975 = P3_REG3_REG_0_ & ~P3_STATE_REG;
  assign n16976 = ~n13668 & n16318;
  assign n16977 = n16320 & ~n16973;
  assign n16978 = n16322 & ~n16965;
  assign n16979 = ~n16976 & ~n16977;
  assign n16980 = ~n16978 & n16979;
  assign n16981 = n16307 & ~n16980;
  assign n16982 = ~n16974 & ~n16975;
  assign n16983 = ~n16981 & n16982;
  assign n1696 = ~n16970 | ~n16983;
  assign n16985 = ~n13707 & n2021;
  assign n16986 = P3_DATAO_REG_0_ & ~n2021;
  assign n1701 = n16985 | n16986;
  assign n16988 = ~n13697 & n2021;
  assign n16989 = P3_DATAO_REG_1_ & ~n2021;
  assign n1706 = n16988 | n16989;
  assign n16991 = ~n13750 & n2021;
  assign n16992 = P3_DATAO_REG_2_ & ~n2021;
  assign n1711 = n16991 | n16992;
  assign n16994 = ~n13806_1 & n2021;
  assign n16995 = P3_DATAO_REG_3_ & ~n2021;
  assign n1716 = n16994 | n16995;
  assign n16997 = ~n13871_1 & n2021;
  assign n16998 = P3_DATAO_REG_4_ & ~n2021;
  assign n1721 = n16997 | n16998;
  assign n17000 = ~n13937 & n2021;
  assign n17001 = P3_DATAO_REG_5_ & ~n2021;
  assign n1726 = n17000 | n17001;
  assign n17003 = ~n14007 & n2021;
  assign n17004 = P3_DATAO_REG_6_ & ~n2021;
  assign n1731 = n17003 | n17004;
  assign n17006 = ~n14098 & n2021;
  assign n17007 = P3_DATAO_REG_7_ & ~n2021;
  assign n1736 = n17006 | n17007;
  assign n17009 = ~n14165 & n2021;
  assign n17010 = P3_DATAO_REG_8_ & ~n2021;
  assign n1741 = n17009 | n17010;
  assign n17012 = ~n14224 & n2021;
  assign n17013 = P3_DATAO_REG_9_ & ~n2021;
  assign n1746 = n17012 | n17013;
  assign n17015 = ~n14292 & n2021;
  assign n17016 = P3_DATAO_REG_10_ & ~n2021;
  assign n1751 = n17015 | n17016;
  assign n17018 = ~n14348 & n2021;
  assign n17019 = P3_DATAO_REG_11_ & ~n2021;
  assign n1756 = n17018 | n17019;
  assign n17021 = ~n14458 & n2021;
  assign n17022 = P3_DATAO_REG_12_ & ~n2021;
  assign n1761 = n17021 | n17022;
  assign n17024 = ~n14524 & n2021;
  assign n17025 = P3_DATAO_REG_13_ & ~n2021;
  assign n1766 = n17024 | n17025;
  assign n17027 = ~n14588 & n2021;
  assign n17028 = P3_DATAO_REG_14_ & ~n2021;
  assign n1771 = n17027 | n17028;
  assign n17030 = ~n14651_1 & n2021;
  assign n17031 = P3_DATAO_REG_15_ & ~n2021;
  assign n1776 = n17030 | n17031;
  assign n17033 = ~n14712 & n2021;
  assign n17034 = P3_DATAO_REG_16_ & ~n2021;
  assign n1781 = n17033 | n17034;
  assign n17036 = ~n14779 & n2021;
  assign n17037 = P3_DATAO_REG_17_ & ~n2021;
  assign n1786 = n17036 | n17037;
  assign n17039 = ~n14846_1 & n2021;
  assign n17040 = P3_DATAO_REG_18_ & ~n2021;
  assign n1791 = n17039 | n17040;
  assign n17042 = ~n14912 & n2021;
  assign n17043 = P3_DATAO_REG_19_ & ~n2021;
  assign n1796 = n17042 | n17043;
  assign n17045 = ~n14974 & n2021;
  assign n17046 = P3_DATAO_REG_20_ & ~n2021;
  assign n1801 = n17045 | n17046;
  assign n17048 = ~n15033 & n2021;
  assign n17049 = P3_DATAO_REG_21_ & ~n2021;
  assign n1806 = n17048 | n17049;
  assign n17051 = ~n15090 & n2021;
  assign n17052 = P3_DATAO_REG_22_ & ~n2021;
  assign n1811 = n17051 | n17052;
  assign n17054 = ~n15150 & n2021;
  assign n17055 = P3_DATAO_REG_23_ & ~n2021;
  assign n1816 = n17054 | n17055;
  assign n17057 = ~n15207 & n2021;
  assign n17058 = P3_DATAO_REG_24_ & ~n2021;
  assign n1821 = n17057 | n17058;
  assign n17060 = ~n15269 & n2021;
  assign n17061 = P3_DATAO_REG_25_ & ~n2021;
  assign n1826 = n17060 | n17061;
  assign n17063 = ~n15324 & n2021;
  assign n17064 = P3_DATAO_REG_26_ & ~n2021;
  assign n1831 = n17063 | n17064;
  assign n17066 = ~n15382 & n2021;
  assign n17067 = P3_DATAO_REG_27_ & ~n2021;
  assign n1836 = n17066 | n17067;
  assign n17069 = ~n15439 & n2021;
  assign n17070 = P3_DATAO_REG_28_ & ~n2021;
  assign n1841 = n17069 | n17070;
  assign n17072 = ~n15501_1 & n2021;
  assign n17073 = P3_DATAO_REG_29_ & ~n2021;
  assign n1846 = n17072 | n17073;
  assign n17075 = ~n15555 & n2021;
  assign n17076 = P3_DATAO_REG_30_ & ~n2021;
  assign n1851 = n17075 | n17076;
  assign n17078 = ~n15578 & n2021;
  assign n17079 = P3_DATAO_REG_31_ & ~n2021;
  assign n1856 = n17078 | n17079;
  assign n17081 = ~n13512 & ~n13581_1;
  assign n17082 = P3_STATE_REG & ~n17081;
  assign n17083 = ~n16104 & n17082;
  assign n17084 = ~n13581_1 & n13721_1;
  assign n17085 = n16111_1 & n17084;
  assign n17086 = n13512 & ~n17085;
  assign n17087 = n17083 & ~n17086;
  assign n17088 = P3_B_REG & ~n17087;
  assign n17089 = n13675 & n14988;
  assign n17090 = ~n15555 & n15578;
  assign n17091 = ~n15578 & ~n17090;
  assign n17092 = n15555 & ~n15578;
  assign n17093 = ~n17090 & ~n17092;
  assign n17094 = n17090 & n17093;
  assign n17095 = ~n17091 & ~n17094;
  assign n17096 = ~n13512 & n13593;
  assign n17097 = ~n17081 & ~n17096;
  assign n17098 = ~n17095 & ~n17097;
  assign n17099 = ~n17089 & ~n17098;
  assign n17100 = n13675 & ~n17095;
  assign n17101 = n14988 & ~n17097;
  assign n17102 = ~n17100 & ~n17101;
  assign n17103 = ~n17099 & n17102;
  assign n17104 = n17099 & ~n17102;
  assign n17105 = ~n17103 & ~n17104;
  assign n17106 = ~n15555 & ~n17090;
  assign n17107 = n15555 & n17090;
  assign n17108 = ~n17106 & ~n17107;
  assign n17109 = ~n17097 & ~n17108;
  assign n17110 = ~n17089 & ~n17109;
  assign n17111 = n13675 & ~n17108;
  assign n17112 = ~n17101 & ~n17111;
  assign n17113 = ~n17110 & n17112;
  assign n17114 = n17110 & ~n17112;
  assign n17115 = ~n13512 & ~n17089;
  assign n17116 = ~n15501_1 & ~n17090;
  assign n17117 = ~n15501_1 & n17090;
  assign n17118 = ~n17116 & ~n17117;
  assign n17119 = ~n17097 & ~n17118;
  assign n17120 = n17115 & ~n17119;
  assign n17121 = n13675 & ~n17118;
  assign n17122 = n13512 & ~n15439;
  assign n17123 = ~n17101 & ~n17121;
  assign n17124 = ~n17122 & n17123;
  assign n17125 = ~n17114 & ~n17120;
  assign n17126 = n17124 & n17125;
  assign n17127 = ~n17113 & ~n17126;
  assign n17128 = n17105 & ~n17127;
  assign n17129 = n13512 & ~n15269;
  assign n17130 = ~n17101 & ~n17129;
  assign n17131 = ~n15324 & ~n17090;
  assign n17132 = ~n15324 & n17090;
  assign n17133 = ~n17131 & ~n17132;
  assign n17134 = n13675 & ~n17133;
  assign n17135 = n17130 & ~n17134;
  assign n17136 = ~n17097 & ~n17133;
  assign n17137 = n17115 & ~n17136;
  assign n17138 = ~n17135 & n17137;
  assign n17139 = n13512 & ~n15324;
  assign n17140 = ~n17101 & ~n17139;
  assign n17141 = ~n15382 & ~n17090;
  assign n17142 = ~n15382 & n17090;
  assign n17143 = ~n17141 & ~n17142;
  assign n17144 = n13675 & ~n17143;
  assign n17145 = n17140 & ~n17144;
  assign n17146 = ~n17097 & ~n17143;
  assign n17147 = n17115 & ~n17146;
  assign n17148 = ~n17145 & n17147;
  assign n17149 = n17105 & ~n17114;
  assign n17150 = ~n17138 & n17149;
  assign n17151 = ~n17148 & n17150;
  assign n17152 = ~n15269 & ~n17090;
  assign n17153 = ~n15269 & n17090;
  assign n17154 = ~n17152 & ~n17153;
  assign n17155 = ~n17097 & ~n17154;
  assign n17156 = n17115 & ~n17155;
  assign n17157 = n13512 & ~n15207;
  assign n17158 = ~n17101 & ~n17157;
  assign n17159 = n13675 & ~n17154;
  assign n17160 = n17158 & ~n17159;
  assign n17161 = ~n17156 & n17160;
  assign n17162 = n17135 & ~n17137;
  assign n17163 = ~n17161 & ~n17162;
  assign n17164 = n13512 & ~n15382;
  assign n17165 = ~n17101 & ~n17164;
  assign n17166 = ~n15439 & ~n17090;
  assign n17167 = ~n15439 & n17090;
  assign n17168 = ~n17166 & ~n17167;
  assign n17169 = n13675 & ~n17168;
  assign n17170 = n17165 & ~n17169;
  assign n17171 = ~n17097 & ~n17168;
  assign n17172 = n17115 & ~n17171;
  assign n17173 = ~n17170 & n17172;
  assign n17174 = n17120 & ~n17124;
  assign n17175 = ~n17173 & ~n17174;
  assign n17176 = n17151 & ~n17163;
  assign n17177 = n17175 & n17176;
  assign n17178 = ~n17128 & ~n17177;
  assign n17179 = ~n15033 & ~n17090;
  assign n17180 = ~n15033 & n17090;
  assign n17181 = ~n17179 & ~n17180;
  assign n17182 = ~n17097 & ~n17181;
  assign n17183 = n17115 & ~n17182;
  assign n17184 = n13512 & ~n14974;
  assign n17185 = ~n17101 & ~n17184;
  assign n17186 = n13675 & ~n17181;
  assign n17187 = n17185 & ~n17186;
  assign n17188 = ~n17183 & n17187;
  assign n17189 = ~n14974 & ~n17090;
  assign n17190 = ~n14974 & n17090;
  assign n17191 = ~n17189 & ~n17190;
  assign n17192 = ~n17097 & ~n17191;
  assign n17193 = n17115 & ~n17192;
  assign n17194 = n13512 & ~n14912;
  assign n17195 = ~n17101 & ~n17194;
  assign n17196 = n13675 & ~n17191;
  assign n17197 = n17195 & ~n17196;
  assign n17198 = ~n17193 & n17197;
  assign n17199 = n13675 & ~n14929;
  assign n17200 = ~n13512 & ~n17199;
  assign n17201 = ~n14912 & ~n17090;
  assign n17202 = ~n14912 & n17090;
  assign n17203 = ~n17201 & ~n17202;
  assign n17204 = ~n17097 & ~n17203;
  assign n17205 = n17200 & ~n17204;
  assign n17206 = n13512 & ~n14846_1;
  assign n17207 = ~n14929 & ~n17097;
  assign n17208 = ~n17206 & ~n17207;
  assign n17209 = n13675 & ~n17203;
  assign n17210 = n17208 & ~n17209;
  assign n17211 = ~n17205 & n17210;
  assign n17212 = n13512 & ~n14651_1;
  assign n17213 = ~n14731_1 & ~n17097;
  assign n17214 = ~n17212 & ~n17213;
  assign n17215 = ~n14712 & ~n17090;
  assign n17216 = ~n14712 & n17090;
  assign n17217 = ~n17215 & ~n17216;
  assign n17218 = n13675 & ~n17217;
  assign n17219 = n17214 & ~n17218;
  assign n17220 = n13675 & ~n14731_1;
  assign n17221 = ~n13512 & ~n17220;
  assign n17222 = ~n17097 & ~n17217;
  assign n17223 = n17221 & ~n17222;
  assign n17224 = ~n17219 & n17223;
  assign n17225 = n13675 & ~n14866_1;
  assign n17226 = ~n13512 & ~n17225;
  assign n17227 = ~n14846_1 & ~n17090;
  assign n17228 = ~n14846_1 & n17090;
  assign n17229 = ~n17227 & ~n17228;
  assign n17230 = ~n17097 & ~n17229;
  assign n17231 = n17226 & ~n17230;
  assign n17232 = n13512 & ~n14779;
  assign n17233 = ~n14866_1 & ~n17097;
  assign n17234 = ~n17232 & ~n17233;
  assign n17235 = n13675 & ~n17229;
  assign n17236 = n17234 & ~n17235;
  assign n17237 = ~n17231 & n17236;
  assign n17238 = n13675 & ~n14798;
  assign n17239 = ~n13512 & ~n17238;
  assign n17240 = ~n14779 & ~n17090;
  assign n17241 = ~n14779 & n17090;
  assign n17242 = ~n17240 & ~n17241;
  assign n17243 = ~n17097 & ~n17242;
  assign n17244 = n17239 & ~n17243;
  assign n17245 = n13512 & ~n14712;
  assign n17246 = ~n14798 & ~n17097;
  assign n17247 = ~n17245 & ~n17246;
  assign n17248 = n13675 & ~n17242;
  assign n17249 = n17247 & ~n17248;
  assign n17250 = ~n17244 & n17249;
  assign n17251 = ~n17237 & ~n17250;
  assign n17252 = n17224 & n17251;
  assign n17253 = n13675 & ~n14670;
  assign n17254 = ~n13512 & ~n17253;
  assign n17255 = ~n14651_1 & ~n17090;
  assign n17256 = ~n14651_1 & n17090;
  assign n17257 = ~n17255 & ~n17256;
  assign n17258 = ~n17097 & ~n17257;
  assign n17259 = n17254 & ~n17258;
  assign n17260 = n13512 & ~n14588;
  assign n17261 = ~n14670 & ~n17097;
  assign n17262 = ~n17260 & ~n17261;
  assign n17263 = n13675 & ~n17257;
  assign n17264 = n17262 & ~n17263;
  assign n17265 = ~n17259 & n17264;
  assign n17266 = n17219 & ~n17223;
  assign n17267 = ~n17265 & ~n17266;
  assign n17268 = n13675 & ~n14609;
  assign n17269 = ~n13512 & ~n17268;
  assign n17270 = ~n14588 & ~n17090;
  assign n17271 = ~n14588 & n17090;
  assign n17272 = ~n17270 & ~n17271;
  assign n17273 = ~n17097 & ~n17272;
  assign n17274 = n17269 & ~n17273;
  assign n17275 = n13512 & ~n14524;
  assign n17276 = ~n14609 & ~n17097;
  assign n17277 = ~n17275 & ~n17276;
  assign n17278 = n13675 & ~n17272;
  assign n17279 = n17277 & ~n17278;
  assign n17280 = ~n17274 & n17279;
  assign n17281 = n13675 & ~n14543;
  assign n17282 = ~n13512 & ~n17281;
  assign n17283 = ~n14524 & ~n17090;
  assign n17284 = ~n14524 & n17090;
  assign n17285 = ~n17283 & ~n17284;
  assign n17286 = ~n17097 & ~n17285;
  assign n17287 = n17282 & ~n17286;
  assign n17288 = n13512 & ~n14458;
  assign n17289 = ~n14543 & ~n17097;
  assign n17290 = ~n17288 & ~n17289;
  assign n17291 = n13675 & ~n17285;
  assign n17292 = n17290 & ~n17291;
  assign n17293 = ~n17287 & n17292;
  assign n17294 = n17287 & ~n17292;
  assign n17295 = n13512 & ~n14292;
  assign n17296 = ~n14407 & ~n17097;
  assign n17297 = ~n17295 & ~n17296;
  assign n17298 = ~n14348 & ~n17090;
  assign n17299 = ~n14348 & n17090;
  assign n17300 = ~n17298 & ~n17299;
  assign n17301 = n13675 & ~n17300;
  assign n17302 = n17297 & ~n17301;
  assign n17303 = n13675 & ~n14407;
  assign n17304 = ~n13512 & ~n17303;
  assign n17305 = ~n17097 & ~n17300;
  assign n17306 = n17304 & ~n17305;
  assign n17307 = ~n17302 & n17306;
  assign n17308 = n13675 & ~n14477;
  assign n17309 = ~n13512 & ~n17308;
  assign n17310 = ~n14458 & ~n17090;
  assign n17311 = ~n14458 & n17090;
  assign n17312 = ~n17310 & ~n17311;
  assign n17313 = ~n17097 & ~n17312;
  assign n17314 = n17309 & ~n17313;
  assign n17315 = n13512 & ~n14348;
  assign n17316 = ~n14477 & ~n17097;
  assign n17317 = ~n17315 & ~n17316;
  assign n17318 = n13675 & ~n17312;
  assign n17319 = n17317 & ~n17318;
  assign n17320 = ~n17314 & n17319;
  assign n17321 = n17307 & ~n17320;
  assign n17322 = ~n17294 & ~n17321;
  assign n17323 = n13512 & ~n14165;
  assign n17324 = ~n14276_1 & ~n17097;
  assign n17325 = ~n17323 & ~n17324;
  assign n17326 = ~n14224 & ~n17090;
  assign n17327 = ~n14224 & n17090;
  assign n17328 = ~n17326 & ~n17327;
  assign n17329 = n13675 & ~n17328;
  assign n17330 = n17325 & ~n17329;
  assign n17331 = n13675 & ~n14276_1;
  assign n17332 = ~n13512 & ~n17331;
  assign n17333 = ~n17097 & ~n17328;
  assign n17334 = n17332 & ~n17333;
  assign n17335 = ~n17330 & n17334;
  assign n17336 = n13512 & ~n14098;
  assign n17337 = ~n14208 & ~n17097;
  assign n17338 = ~n17336 & ~n17337;
  assign n17339 = ~n14165 & ~n17090;
  assign n17340 = ~n14165 & n17090;
  assign n17341 = ~n17339 & ~n17340;
  assign n17342 = n13675 & ~n17341;
  assign n17343 = n17338 & ~n17342;
  assign n17344 = n13675 & ~n14208;
  assign n17345 = ~n13512 & ~n17344;
  assign n17346 = ~n17097 & ~n17341;
  assign n17347 = n17345 & ~n17346;
  assign n17348 = ~n17343 & n17347;
  assign n17349 = ~n17335 & ~n17348;
  assign n17350 = n13512 & ~n14007;
  assign n17351 = ~n14139 & ~n17097;
  assign n17352 = ~n17350 & ~n17351;
  assign n17353 = ~n14098 & ~n17090;
  assign n17354 = ~n14098 & n17090;
  assign n17355 = ~n17353 & ~n17354;
  assign n17356 = n13675 & ~n17355;
  assign n17357 = n17352 & ~n17356;
  assign n17358 = n13675 & ~n14139;
  assign n17359 = ~n13512 & ~n17358;
  assign n17360 = ~n17097 & ~n17355;
  assign n17361 = n17359 & ~n17360;
  assign n17362 = ~n17357 & n17361;
  assign n17363 = n13512 & ~n13937;
  assign n17364 = ~n14066_1 & ~n17097;
  assign n17365 = ~n17363 & ~n17364;
  assign n17366 = ~n14007 & ~n17090;
  assign n17367 = ~n14007 & n17090;
  assign n17368 = ~n17366 & ~n17367;
  assign n17369 = n13675 & ~n17368;
  assign n17370 = n17365 & ~n17369;
  assign n17371 = n13675 & ~n14066_1;
  assign n17372 = ~n13512 & ~n17371;
  assign n17373 = ~n17097 & ~n17368;
  assign n17374 = n17372 & ~n17373;
  assign n17375 = ~n17370 & n17374;
  assign n17376 = ~n17362 & ~n17375;
  assign n17377 = n17349 & n17376;
  assign n17378 = n13675 & ~n13944;
  assign n17379 = ~n13512 & ~n17378;
  assign n17380 = ~n13871_1 & ~n17090;
  assign n17381 = ~n13871_1 & n17090;
  assign n17382 = ~n17380 & ~n17381;
  assign n17383 = ~n17097 & ~n17382;
  assign n17384 = n17379 & ~n17383;
  assign n17385 = n13512 & ~n13806_1;
  assign n17386 = ~n13944 & ~n17097;
  assign n17387 = ~n17385 & ~n17386;
  assign n17388 = n13675 & ~n17382;
  assign n17389 = n17387 & ~n17388;
  assign n17390 = ~n17384 & n17389;
  assign n17391 = n13675 & ~n13878;
  assign n17392 = ~n13512 & ~n17391;
  assign n17393 = ~n13806_1 & ~n17090;
  assign n17394 = ~n13806_1 & n17090;
  assign n17395 = ~n17393 & ~n17394;
  assign n17396 = ~n17097 & ~n17395;
  assign n17397 = n17392 & ~n17396;
  assign n17398 = n13512 & ~n13750;
  assign n17399 = ~n13878 & ~n17097;
  assign n17400 = ~n17398 & ~n17399;
  assign n17401 = n13675 & ~n17395;
  assign n17402 = n17400 & ~n17401;
  assign n17403 = ~n17397 & n17402;
  assign n17404 = n13675 & ~n13813;
  assign n17405 = ~n13512 & ~n17404;
  assign n17406 = ~n13750 & ~n17090;
  assign n17407 = ~n13750 & n17090;
  assign n17408 = ~n17406 & ~n17407;
  assign n17409 = ~n17097 & ~n17408;
  assign n17410 = n17405 & ~n17409;
  assign n17411 = n13512 & ~n13697;
  assign n17412 = ~n13813 & ~n17097;
  assign n17413 = ~n17411 & ~n17412;
  assign n17414 = n13675 & ~n17408;
  assign n17415 = n17413 & ~n17414;
  assign n17416 = ~n17410 & n17415;
  assign n17417 = n13675 & ~n13757;
  assign n17418 = ~n13512 & ~n17417;
  assign n17419 = ~n13697 & ~n17090;
  assign n17420 = ~n13697 & n17090;
  assign n17421 = ~n17419 & ~n17420;
  assign n17422 = ~n17097 & ~n17421;
  assign n17423 = n17418 & ~n17422;
  assign n17424 = n13512 & ~n13707;
  assign n17425 = ~n13757 & ~n17097;
  assign n17426 = ~n17424 & ~n17425;
  assign n17427 = n13675 & ~n17421;
  assign n17428 = n17426 & ~n17427;
  assign n17429 = ~n17423 & n17428;
  assign n17430 = n17410 & ~n17415;
  assign n17431 = n17429 & ~n17430;
  assign n17432 = ~n17416 & ~n17431;
  assign n17433 = n17397 & ~n17402;
  assign n17434 = ~n17432 & ~n17433;
  assign n17435 = ~n17403 & ~n17434;
  assign n17436 = n17384 & ~n17389;
  assign n17437 = ~n17435 & ~n17436;
  assign n17438 = ~n17390 & ~n17437;
  assign n17439 = n13512 & ~n13871_1;
  assign n17440 = ~n14014 & ~n17097;
  assign n17441 = ~n17439 & ~n17440;
  assign n17442 = ~n13937 & ~n17090;
  assign n17443 = ~n13937 & n17090;
  assign n17444 = ~n17442 & ~n17443;
  assign n17445 = n13675 & ~n17444;
  assign n17446 = n17441 & ~n17445;
  assign n17447 = n13675 & ~n14014;
  assign n17448 = ~n13512 & ~n17447;
  assign n17449 = ~n17097 & ~n17444;
  assign n17450 = n17448 & ~n17449;
  assign n17451 = ~n17446 & n17450;
  assign n17452 = ~n17438 & ~n17451;
  assign n17453 = n17370 & ~n17374;
  assign n17454 = n17446 & ~n17450;
  assign n17455 = ~n17453 & ~n17454;
  assign n17456 = ~n13671_1 & n13675;
  assign n17457 = ~n13512 & ~n17456;
  assign n17458 = ~n13707 & ~n17090;
  assign n17459 = ~n13707 & n17090;
  assign n17460 = ~n17458 & ~n17459;
  assign n17461 = ~n17097 & ~n17460;
  assign n17462 = n17457 & ~n17461;
  assign n17463 = ~n13512 & n13675;
  assign n17464 = n17462 & n17463;
  assign n17465 = n17423 & ~n17428;
  assign n17466 = n13675 & ~n17460;
  assign n17467 = ~n13671_1 & ~n17097;
  assign n17468 = ~n17466 & ~n17467;
  assign n17469 = ~n17462 & ~n17463;
  assign n17470 = ~n17468 & ~n17469;
  assign n17471 = ~n17464 & ~n17465;
  assign n17472 = ~n17470 & n17471;
  assign n17473 = ~n17430 & ~n17433;
  assign n17474 = ~n17451 & n17473;
  assign n17475 = ~n17436 & n17474;
  assign n17476 = n17472 & n17475;
  assign n17477 = n17455 & ~n17476;
  assign n17478 = ~n17452 & n17477;
  assign n17479 = n17377 & ~n17478;
  assign n17480 = n17357 & ~n17361;
  assign n17481 = n17349 & n17480;
  assign n17482 = n17343 & ~n17347;
  assign n17483 = ~n17335 & n17482;
  assign n17484 = n13675 & ~n14355;
  assign n17485 = ~n13512 & ~n17484;
  assign n17486 = ~n14292 & ~n17090;
  assign n17487 = ~n14292 & n17090;
  assign n17488 = ~n17486 & ~n17487;
  assign n17489 = ~n17097 & ~n17488;
  assign n17490 = n17485 & ~n17489;
  assign n17491 = n13512 & ~n14224;
  assign n17492 = ~n14355 & ~n17097;
  assign n17493 = ~n17491 & ~n17492;
  assign n17494 = n13675 & ~n17488;
  assign n17495 = n17493 & ~n17494;
  assign n17496 = ~n17490 & n17495;
  assign n17497 = n17330 & ~n17334;
  assign n17498 = ~n17496 & ~n17497;
  assign n17499 = ~n17481 & ~n17483;
  assign n17500 = n17498 & n17499;
  assign n17501 = n17302 & ~n17306;
  assign n17502 = ~n17320 & ~n17501;
  assign n17503 = ~n17479 & n17500;
  assign n17504 = n17502 & n17503;
  assign n17505 = n17490 & ~n17495;
  assign n17506 = n17502 & n17505;
  assign n17507 = n17314 & ~n17319;
  assign n17508 = ~n17506 & ~n17507;
  assign n17509 = n17322 & ~n17504;
  assign n17510 = n17508 & n17509;
  assign n17511 = ~n17293 & ~n17510;
  assign n17512 = n17274 & ~n17279;
  assign n17513 = ~n17511 & ~n17512;
  assign n17514 = ~n17280 & ~n17513;
  assign n17515 = n17259 & ~n17264;
  assign n17516 = ~n17514 & ~n17515;
  assign n17517 = n17267 & ~n17516;
  assign n17518 = n17251 & n17517;
  assign n17519 = n17244 & ~n17249;
  assign n17520 = ~n17237 & n17519;
  assign n17521 = n17231 & ~n17236;
  assign n17522 = n17205 & ~n17210;
  assign n17523 = ~n17520 & ~n17521;
  assign n17524 = ~n17522 & n17523;
  assign n17525 = ~n17252 & ~n17518;
  assign n17526 = n17524 & n17525;
  assign n17527 = ~n17211 & ~n17526;
  assign n17528 = n17193 & ~n17197;
  assign n17529 = ~n17527 & ~n17528;
  assign n17530 = ~n17198 & ~n17529;
  assign n17531 = n17183 & ~n17187;
  assign n17532 = ~n17530 & ~n17531;
  assign n17533 = ~n15090 & ~n17090;
  assign n17534 = ~n15090 & n17090;
  assign n17535 = ~n17533 & ~n17534;
  assign n17536 = ~n17097 & ~n17535;
  assign n17537 = n17115 & ~n17536;
  assign n17538 = n13512 & ~n15033;
  assign n17539 = ~n17101 & ~n17538;
  assign n17540 = n13675 & ~n17535;
  assign n17541 = n17539 & ~n17540;
  assign n17542 = ~n17537 & n17541;
  assign n17543 = ~n15207 & ~n17090;
  assign n17544 = ~n15207 & n17090;
  assign n17545 = ~n17543 & ~n17544;
  assign n17546 = ~n17097 & ~n17545;
  assign n17547 = n17115 & ~n17546;
  assign n17548 = n13512 & ~n15150;
  assign n17549 = ~n17101 & ~n17548;
  assign n17550 = n13675 & ~n17545;
  assign n17551 = n17549 & ~n17550;
  assign n17552 = ~n17547 & n17551;
  assign n17553 = ~n15150 & ~n17090;
  assign n17554 = ~n15150 & n17090;
  assign n17555 = ~n17553 & ~n17554;
  assign n17556 = ~n17097 & ~n17555;
  assign n17557 = n17115 & ~n17556;
  assign n17558 = n13512 & ~n15090;
  assign n17559 = ~n17101 & ~n17558;
  assign n17560 = n13675 & ~n17555;
  assign n17561 = n17559 & ~n17560;
  assign n17562 = ~n17557 & n17561;
  assign n17563 = ~n17552 & ~n17562;
  assign n17564 = ~n17188 & ~n17532;
  assign n17565 = ~n17542 & n17564;
  assign n17566 = n17563 & n17565;
  assign n17567 = n17557 & ~n17561;
  assign n17568 = ~n17552 & n17567;
  assign n17569 = ~n17173 & ~n17568;
  assign n17570 = n17156 & ~n17160;
  assign n17571 = n17547 & ~n17551;
  assign n17572 = ~n17570 & ~n17571;
  assign n17573 = n17537 & ~n17541;
  assign n17574 = n17563 & n17573;
  assign n17575 = n17572 & ~n17574;
  assign n17576 = n17151 & n17575;
  assign n17577 = ~n17174 & ~n17566;
  assign n17578 = n17569 & n17577;
  assign n17579 = n17576 & n17578;
  assign n17580 = n13512 & ~n13675;
  assign n17581 = n17102 & n17580;
  assign n17582 = ~n17099 & n17581;
  assign n17583 = ~n17102 & ~n17580;
  assign n17584 = n17099 & n17583;
  assign n17585 = ~n17582 & ~n17584;
  assign n17586 = n17145 & ~n17147;
  assign n17587 = ~n17170 & ~n17586;
  assign n17588 = n17172 & ~n17586;
  assign n17589 = ~n17174 & ~n17588;
  assign n17590 = ~n17173 & n17589;
  assign n17591 = n17149 & ~n17587;
  assign n17592 = n17590 & n17591;
  assign n17593 = n17585 & ~n17592;
  assign n17594 = n17178 & ~n17579;
  assign n17595 = n17593 & n17594;
  assign n17596 = n13525 & n17085;
  assign n17597 = n17595 & n17596;
  assign n17598 = ~n17088 & ~n17597;
  assign n17599 = ~n13512 & n13581_1;
  assign n17600 = n17595 & n17599;
  assign n17601 = ~n13587 & n17600;
  assign n17602 = ~n14988 & n15324;
  assign n17603 = ~n15349 & ~n17602;
  assign n17604 = ~n15298 & ~n17603;
  assign n17605 = ~n15177 & ~n15178;
  assign n17606 = ~n15114 & ~n15118;
  assign n17607 = ~n15236_1 & ~n15237;
  assign n17608 = ~n17605 & ~n17606;
  assign n17609 = ~n17607 & n17608;
  assign n17610 = ~n15243 & n17609;
  assign n17611 = n17604 & n17610;
  assign n17612 = ~n14020 & ~n14021_1;
  assign n17613 = ~n13894 & ~n17612;
  assign n17614 = ~n13822 & n17613;
  assign n17615 = ~n14141_1 & ~n14142;
  assign n17616 = ~n14084 & ~n17615;
  assign n17617 = ~n14497 & n17616;
  assign n17618 = n17614 & n17617;
  assign n17619 = ~n14752 & n17618;
  assign n17620 = n13671_1 & n13707;
  assign n17621 = ~n13766_1 & ~n17620;
  assign n17622 = ~n14681_1 & ~n14682;
  assign n17623 = ~n13765 & ~n17621;
  assign n17624 = ~n17622 & n17623;
  assign n17625 = ~n14554 & ~n14555;
  assign n17626 = ~n14238 & ~n14302;
  assign n17627 = ~n17625 & n17626;
  assign n17628 = ~n14745 & ~n14746_1;
  assign n17629 = n17624 & n17627;
  assign n17630 = ~n17628 & n17629;
  assign n17631 = ~n14813 & ~n14815;
  assign n17632 = ~n15467 & ~n15473;
  assign n17633 = n17619 & n17630;
  assign n17634 = ~n17631 & n17633;
  assign n17635 = ~n14886_1 & n17634;
  assign n17636 = ~n17632 & n17635;
  assign n17637 = ~n14356_1 & ~n14357;
  assign n17638 = ~n13961_1 & ~n17637;
  assign n17639 = ~n14431_1 & n17638;
  assign n17640 = ~n14947 & n17639;
  assign n17641 = ~n14988 & n15555;
  assign n17642 = n14988 & ~n15555;
  assign n17643 = ~n17641 & ~n17642;
  assign n17644 = ~n14988 & n15578;
  assign n17645 = n14988 & ~n15578;
  assign n17646 = ~n17644 & ~n17645;
  assign n17647 = ~n17643 & ~n17646;
  assign n17648 = ~n14999 & ~n15001_1;
  assign n17649 = ~n14988 & n15501_1;
  assign n17650 = n14988 & ~n15501_1;
  assign n17651 = ~n17649 & ~n17650;
  assign n17652 = ~n14988 & n15439;
  assign n17653 = ~n15517 & ~n17652;
  assign n17654 = n17640 & n17647;
  assign n17655 = ~n17648 & n17654;
  assign n17656 = ~n17651 & n17655;
  assign n17657 = ~n17653 & n17656;
  assign n17658 = n17611 & n17636;
  assign n17659 = n17657 & n17658;
  assign n17660 = n17096 & n17659;
  assign n17661 = ~n13512 & ~n13593;
  assign n17662 = ~n17659 & n17661;
  assign n17663 = ~n17660 & ~n17662;
  assign n17664 = n13587 & ~n17663;
  assign n17665 = ~n14988 & ~n17095;
  assign n17666 = n14988 & n17108;
  assign n17667 = ~n17665 & ~n17666;
  assign n17668 = n14988 & n17143;
  assign n17669 = n14988 & n17133;
  assign n17670 = n14988 & n17545;
  assign n17671 = ~n14988 & ~n17555;
  assign n17672 = n14988 & n17154;
  assign n17673 = ~n17670 & n17671;
  assign n17674 = ~n17672 & n17673;
  assign n17675 = ~n14670 & n17257;
  assign n17676 = ~n14609 & n17272;
  assign n17677 = n14477 & ~n17312;
  assign n17678 = ~n14543 & n17285;
  assign n17679 = n17677 & ~n17678;
  assign n17680 = n14407 & ~n17300;
  assign n17681 = ~n14477 & n17312;
  assign n17682 = ~n17678 & ~n17681;
  assign n17683 = n17680 & n17682;
  assign n17684 = ~n17679 & ~n17683;
  assign n17685 = ~n14407 & n17300;
  assign n17686 = ~n14355 & n17488;
  assign n17687 = ~n17685 & ~n17686;
  assign n17688 = ~n14276_1 & n17328;
  assign n17689 = ~n14208 & n17341;
  assign n17690 = n14208 & ~n17341;
  assign n17691 = n14139 & ~n17355;
  assign n17692 = ~n17690 & ~n17691;
  assign n17693 = n14066_1 & ~n17368;
  assign n17694 = ~n14139 & n17355;
  assign n17695 = n17693 & ~n17694;
  assign n17696 = n17692 & ~n17695;
  assign n17697 = ~n14014 & n17444;
  assign n17698 = ~n13944 & n17382;
  assign n17699 = ~n13878 & n17395;
  assign n17700 = n13944 & ~n17382;
  assign n17701 = n17699 & ~n17700;
  assign n17702 = ~n14066_1 & n17368;
  assign n17703 = ~n17694 & ~n17702;
  assign n17704 = ~n17698 & ~n17701;
  assign n17705 = n17703 & n17704;
  assign n17706 = n14014 & ~n17444;
  assign n17707 = n17703 & n17706;
  assign n17708 = ~n17705 & ~n17707;
  assign n17709 = ~n17697 & ~n17708;
  assign n17710 = n17696 & ~n17709;
  assign n17711 = ~n17689 & ~n17710;
  assign n17712 = n14276_1 & ~n17328;
  assign n17713 = ~n17711 & ~n17712;
  assign n17714 = ~n17688 & ~n17713;
  assign n17715 = n14355 & ~n17488;
  assign n17716 = ~n17714 & ~n17715;
  assign n17717 = ~n13813 & n17408;
  assign n17718 = n13878 & ~n17395;
  assign n17719 = ~n17700 & ~n17718;
  assign n17720 = ~n17691 & n17719;
  assign n17721 = ~n17690 & n17720;
  assign n17722 = ~n17695 & ~n17707;
  assign n17723 = ~n17712 & n17722;
  assign n17724 = n17721 & n17723;
  assign n17725 = ~n17715 & n17724;
  assign n17726 = n17717 & n17725;
  assign n17727 = ~n13671_1 & n17460;
  assign n17728 = n13757 & ~n17727;
  assign n17729 = n13813 & ~n17408;
  assign n17730 = ~n17728 & ~n17729;
  assign n17731 = ~n13757 & n17727;
  assign n17732 = ~n17421 & ~n17731;
  assign n17733 = n17730 & ~n17732;
  assign n17734 = n17725 & n17733;
  assign n17735 = ~n17726 & ~n17734;
  assign n17736 = n17687 & ~n17716;
  assign n17737 = n17735 & n17736;
  assign n17738 = n17682 & n17737;
  assign n17739 = n14543 & ~n17285;
  assign n17740 = n14609 & ~n17272;
  assign n17741 = ~n17739 & ~n17740;
  assign n17742 = n17684 & ~n17738;
  assign n17743 = n17741 & n17742;
  assign n17744 = ~n17676 & ~n17743;
  assign n17745 = n14670 & ~n17257;
  assign n17746 = ~n17744 & ~n17745;
  assign n17747 = ~n17675 & ~n17746;
  assign n17748 = n14731_1 & ~n17217;
  assign n17749 = n14929 & ~n17203;
  assign n17750 = n14866_1 & ~n17229;
  assign n17751 = ~n14929 & n17203;
  assign n17752 = n17750 & ~n17751;
  assign n17753 = ~n17749 & ~n17752;
  assign n17754 = n14798 & ~n17242;
  assign n17755 = ~n14866_1 & n17229;
  assign n17756 = ~n17751 & ~n17755;
  assign n17757 = n17754 & n17756;
  assign n17758 = ~n14988 & ~n17191;
  assign n17759 = ~n14988 & ~n17535;
  assign n17760 = ~n14988 & ~n17181;
  assign n17761 = ~n17759 & ~n17760;
  assign n17762 = n17753 & ~n17757;
  assign n17763 = ~n17758 & n17762;
  assign n17764 = n17761 & n17763;
  assign n17765 = ~n17747 & ~n17748;
  assign n17766 = n17764 & n17765;
  assign n17767 = ~n14731_1 & n17217;
  assign n17768 = ~n14798 & n17242;
  assign n17769 = ~n17767 & ~n17768;
  assign n17770 = n17756 & n17769;
  assign n17771 = n17764 & ~n17770;
  assign n17772 = n14988 & n17555;
  assign n17773 = n14988 & n17535;
  assign n17774 = ~n17772 & ~n17773;
  assign n17775 = n14988 & n17191;
  assign n17776 = n17761 & n17775;
  assign n17777 = n14988 & n17181;
  assign n17778 = ~n17759 & n17777;
  assign n17779 = ~n17776 & ~n17778;
  assign n17780 = ~n17670 & n17779;
  assign n17781 = ~n17672 & n17780;
  assign n17782 = ~n17766 & ~n17771;
  assign n17783 = n17774 & n17782;
  assign n17784 = n17781 & n17783;
  assign n17785 = ~n14988 & ~n17154;
  assign n17786 = ~n14988 & ~n17545;
  assign n17787 = ~n17785 & ~n17786;
  assign n17788 = ~n17672 & ~n17787;
  assign n17789 = ~n14988 & ~n17133;
  assign n17790 = ~n17788 & ~n17789;
  assign n17791 = ~n17674 & ~n17784;
  assign n17792 = n17790 & n17791;
  assign n17793 = ~n17669 & ~n17792;
  assign n17794 = ~n14988 & ~n17143;
  assign n17795 = ~n17793 & ~n17794;
  assign n17796 = ~n17668 & ~n17795;
  assign n17797 = n14988 & ~n17796;
  assign n17798 = ~n14988 & ~n17668;
  assign n17799 = ~n17795 & n17798;
  assign n17800 = n17168 & ~n17799;
  assign n17801 = n14988 & n17118;
  assign n17802 = n17667 & ~n17797;
  assign n17803 = ~n17800 & n17802;
  assign n17804 = ~n17801 & n17803;
  assign n17805 = n14988 & n17095;
  assign n17806 = ~n14988 & ~n17108;
  assign n17807 = ~n17665 & n17806;
  assign n17808 = ~n17805 & ~n17807;
  assign n17809 = ~n14988 & n17667;
  assign n17810 = ~n17118 & n17809;
  assign n17811 = n17808 & ~n17810;
  assign n17812 = ~n17804 & n17811;
  assign n17813 = n13679 & n17096;
  assign n17814 = n17812 & n17813;
  assign n17815 = ~n17601 & ~n17664;
  assign n17816 = ~n17814 & n17815;
  assign n17817 = ~n13584 & ~n17816;
  assign n17818 = n15164 & ~n15222;
  assign n17819 = ~n15221_1 & ~n17818;
  assign n17820 = ~n15283 & n17819;
  assign n17821 = ~n15338 & n17820;
  assign n17822 = ~n14233 & ~n14295;
  assign n17823 = n14408 & ~n14479;
  assign n17824 = ~n14148 & n17822;
  assign n17825 = ~n14363 & n17824;
  assign n17826 = ~n17823 & n17825;
  assign n17827 = ~n14069 & n17826;
  assign n17828 = n14027 & ~n14068;
  assign n17829 = n17827 & ~n17828;
  assign n17830 = ~n14478 & ~n14544;
  assign n17831 = ~n14610 & ~n14671_1;
  assign n17832 = n14799 & ~n14868;
  assign n17833 = ~n14867 & ~n14930;
  assign n17834 = ~n14989 & ~n17832;
  assign n17835 = n17833 & n17834;
  assign n17836 = ~n14732 & n17835;
  assign n17837 = ~n15049 & n17836;
  assign n17838 = n17831 & n17837;
  assign n17839 = n17830 & n17838;
  assign n17840 = ~n15165 & ~n15222;
  assign n17841 = n15104 & n17840;
  assign n17842 = n17839 & ~n17841;
  assign n17843 = n17829 & n17842;
  assign n17844 = n17821 & n17843;
  assign n17845 = ~n14988 & ~n15555;
  assign n17846 = n14988 & n15578;
  assign n17847 = ~n17845 & ~n17846;
  assign n17848 = ~n15521_1 & n17847;
  assign n17849 = ~n15396_1 & n17848;
  assign n17850 = n13806_1 & ~n13951_1;
  assign n17851 = ~n15453 & n17850;
  assign n17852 = ~n13878 & n17844;
  assign n17853 = n17849 & n17852;
  assign n17854 = n17851 & n17853;
  assign n17855 = ~n14014 & n17827;
  assign n17856 = n17821 & n17855;
  assign n17857 = n13937 & ~n15453;
  assign n17858 = n17842 & n17856;
  assign n17859 = n17849 & n17858;
  assign n17860 = n17857 & n17859;
  assign n17861 = n14007 & ~n15453;
  assign n17862 = n17826 & n17842;
  assign n17863 = n17821 & n17862;
  assign n17864 = ~n14066_1 & n17863;
  assign n17865 = n17849 & n17864;
  assign n17866 = n17861 & n17865;
  assign n17867 = n14651_1 & ~n15453;
  assign n17868 = ~n14670 & n17837;
  assign n17869 = n17821 & n17868;
  assign n17870 = ~n17841 & n17869;
  assign n17871 = n17849 & n17870;
  assign n17872 = n17867 & n17871;
  assign n17873 = ~n17866 & ~n17872;
  assign n17874 = ~n14139 & n17822;
  assign n17875 = ~n14363 & ~n17823;
  assign n17876 = n17842 & n17875;
  assign n17877 = n17821 & n17876;
  assign n17878 = n14098 & n17849;
  assign n17879 = n17874 & n17877;
  assign n17880 = ~n15453 & n17879;
  assign n17881 = n17878 & n17880;
  assign n17882 = ~n14989 & ~n15049;
  assign n17883 = ~n17841 & n17882;
  assign n17884 = n17821 & n17883;
  assign n17885 = n14912 & n17849;
  assign n17886 = ~n14929 & n17884;
  assign n17887 = ~n15453 & n17886;
  assign n17888 = n17885 & n17887;
  assign n17889 = n14524 & ~n15453;
  assign n17890 = ~n14543 & n17838;
  assign n17891 = n17821 & n17890;
  assign n17892 = ~n17841 & n17891;
  assign n17893 = n17849 & n17892;
  assign n17894 = n17889 & n17893;
  assign n17895 = ~n17881 & ~n17888;
  assign n17896 = ~n17894 & n17895;
  assign n17897 = ~n17854 & ~n17860;
  assign n17898 = n17873 & n17897;
  assign n17899 = n17896 & n17898;
  assign n17900 = ~n13889 & ~n13951_1;
  assign n17901 = ~n13827 & n17900;
  assign n17902 = ~n13757 & n17901;
  assign n17903 = n13697 & n17849;
  assign n17904 = n17844 & n17902;
  assign n17905 = ~n15453 & n17904;
  assign n17906 = n17903 & n17905;
  assign n17907 = ~n15284 & ~n15339;
  assign n17908 = ~n15338 & ~n15453;
  assign n17909 = n17849 & ~n17907;
  assign n17910 = n17908 & n17909;
  assign n17911 = ~n14988 & ~n15578;
  assign n17912 = ~n13587 & ~n13671_1;
  assign n17913 = ~n13707 & ~n17912;
  assign n17914 = n13587 & n13671_1;
  assign n17915 = ~n17828 & ~n17913;
  assign n17916 = ~n13774 & n17915;
  assign n17917 = n17901 & n17916;
  assign n17918 = ~n17914 & n17917;
  assign n17919 = n17827 & n17918;
  assign n17920 = n17821 & n17919;
  assign n17921 = ~n15104 & ~n15453;
  assign n17922 = n17839 & n17920;
  assign n17923 = n17849 & n17922;
  assign n17924 = n17921 & n17923;
  assign n17925 = ~n17911 & ~n17924;
  assign n17926 = n14348 & n17849;
  assign n17927 = ~n14407 & n17842;
  assign n17928 = n17821 & n17927;
  assign n17929 = ~n15453 & n17928;
  assign n17930 = n17926 & n17929;
  assign n17931 = n14458 & ~n14544;
  assign n17932 = ~n17841 & n17931;
  assign n17933 = ~n15453 & n17932;
  assign n17934 = ~n14477 & n17838;
  assign n17935 = n17821 & n17934;
  assign n17936 = n17849 & n17935;
  assign n17937 = n17933 & n17936;
  assign n17938 = ~n17930 & ~n17937;
  assign n17939 = n14224 & n17849;
  assign n17940 = ~n14276_1 & n17877;
  assign n17941 = ~n15453 & n17940;
  assign n17942 = n17939 & n17941;
  assign n17943 = ~n17906 & ~n17910;
  assign n17944 = n17925 & n17943;
  assign n17945 = n17938 & n17944;
  assign n17946 = ~n17942 & n17945;
  assign n17947 = n13871_1 & n17849;
  assign n17948 = ~n13944 & n17844;
  assign n17949 = ~n15453 & n17948;
  assign n17950 = n17947 & n17949;
  assign n17951 = n14165 & ~n14295;
  assign n17952 = ~n15453 & n17951;
  assign n17953 = ~n14208 & n17877;
  assign n17954 = n17849 & n17953;
  assign n17955 = n17952 & n17954;
  assign n17956 = n13750 & n17900;
  assign n17957 = ~n15453 & n17956;
  assign n17958 = ~n13813 & n17843;
  assign n17959 = n17821 & n17958;
  assign n17960 = n17849 & n17959;
  assign n17961 = n17957 & n17960;
  assign n17962 = n14292 & ~n15453;
  assign n17963 = ~n14355 & n17842;
  assign n17964 = n17821 & n17963;
  assign n17965 = ~n17823 & n17964;
  assign n17966 = n17849 & n17965;
  assign n17967 = n17962 & n17966;
  assign n17968 = n14588 & ~n14671_1;
  assign n17969 = ~n17841 & n17968;
  assign n17970 = ~n15453 & n17969;
  assign n17971 = ~n14609 & n17837;
  assign n17972 = n17821 & n17971;
  assign n17973 = n17849 & n17972;
  assign n17974 = n17970 & n17973;
  assign n17975 = ~n14731_1 & n17833;
  assign n17976 = ~n17832 & n17849;
  assign n17977 = n14712 & ~n15453;
  assign n17978 = n17884 & n17975;
  assign n17979 = n17976 & n17978;
  assign n17980 = n17977 & n17979;
  assign n17981 = n14974 & ~n15049;
  assign n17982 = ~n17841 & n17981;
  assign n17983 = ~n15453 & n17982;
  assign n17984 = n14988 & n17821;
  assign n17985 = n17849 & n17984;
  assign n17986 = n17983 & n17985;
  assign n17987 = ~n17980 & ~n17986;
  assign n17988 = ~n17967 & ~n17974;
  assign n17989 = n17987 & n17988;
  assign n17990 = n14846_1 & ~n14930;
  assign n17991 = ~n15453 & n17990;
  assign n17992 = ~n14866_1 & n17884;
  assign n17993 = n17849 & n17992;
  assign n17994 = n17991 & n17993;
  assign n17995 = n15227 & n17840;
  assign n17996 = ~n17841 & ~n17995;
  assign n17997 = ~n15453 & n17996;
  assign n17998 = n17821 & n17997;
  assign n17999 = n17849 & n17998;
  assign n18000 = ~n14798 & n17833;
  assign n18001 = n14779 & n17849;
  assign n18002 = n17884 & n18000;
  assign n18003 = ~n15453 & n18002;
  assign n18004 = n18001 & n18003;
  assign n18005 = n14988 & ~n17845;
  assign n18006 = ~n15521_1 & n18005;
  assign n18007 = n15439 & n18006;
  assign n18008 = ~n17846 & n18007;
  assign n18009 = n14988 & n15555;
  assign n18010 = n15501_1 & n18005;
  assign n18011 = ~n18009 & ~n18010;
  assign n18012 = ~n17846 & ~n18011;
  assign n18013 = n14988 & ~n15521_1;
  assign n18014 = ~n17845 & n18013;
  assign n18015 = n15382 & n18014;
  assign n18016 = ~n17846 & n18015;
  assign n18017 = ~n15453 & n18016;
  assign n18018 = ~n18008 & ~n18012;
  assign n18019 = ~n18017 & n18018;
  assign n18020 = ~n17994 & ~n17999;
  assign n18021 = ~n18004 & n18020;
  assign n18022 = n18019 & n18021;
  assign n18023 = ~n17950 & ~n17955;
  assign n18024 = ~n17961 & n18023;
  assign n18025 = n17989 & n18024;
  assign n18026 = n18022 & n18025;
  assign n18027 = n17899 & n17946;
  assign n18028 = n18026 & n18027;
  assign n18029 = n17096 & ~n18028;
  assign n18030 = n13584 & n18029;
  assign n18031 = ~n13512 & n13732;
  assign n18032 = n18028 & n18031;
  assign n18033 = n13725 & n17081;
  assign n18034 = ~n17595 & n18033;
  assign n18035 = ~n18032 & ~n18034;
  assign n18036 = ~n17817 & ~n18030;
  assign n18037 = n18035 & n18036;
  assign n18038 = P3_STATE_REG & ~n18037;
  assign n1861 = ~n17598 | n18038;
  assign n18040 = n13525 & ~n15708;
  assign n18041 = ~n13574 & ~n13578;
  assign n18042 = n13656_1 & n18041;
  assign n18043 = n18040 & ~n18042;
  assign n18044 = n13512 & ~n15699;
  assign n18045 = ~n16104 & n18044;
  assign n18046 = ~n13727 & ~n13733;
  assign n18047 = ~n13730 & n18046;
  assign n18048 = n13587 & ~n18047;
  assign n18049 = ~n13719 & ~n15720;
  assign n18050 = ~n13725 & n18049;
  assign n18051 = n13581_1 & ~n18050;
  assign n18052 = ~n13717 & ~n13722;
  assign n18053 = ~n15697 & n18052;
  assign n18054 = ~n18048 & ~n18051;
  assign n18055 = n18053 & n18054;
  assign n18056 = ~n18042 & ~n18055;
  assign n18057 = n18045 & ~n18056;
  assign n18058 = P3_STATE_REG & ~n18057;
  assign n18059 = ~n18043 & ~n18058;
  assign n18060 = ~n14647 & ~n18059;
  assign n18061 = n18040 & n18042;
  assign n18062 = n13525 & n15698;
  assign n18063 = ~n18061 & ~n18062;
  assign n18064 = ~n14670 & ~n18063;
  assign n18065 = n13525 & n17084;
  assign n18066 = ~n14647 & ~n18042;
  assign n18067 = ~n13664 & n18042;
  assign n18068 = ~n14588 & n18067;
  assign n18069 = n13664 & n18042;
  assign n18070 = ~n14712 & n18069;
  assign n18071 = ~n18066 & ~n18068;
  assign n18072 = ~n18070 & n18071;
  assign n18073 = n18065 & ~n18072;
  assign n18074 = ~n14588 & ~n16846;
  assign n18075 = ~n14609 & n16839;
  assign n18076 = ~n18074 & ~n18075;
  assign n18077 = ~n14588 & n16839;
  assign n18078 = ~n14609 & ~n16855;
  assign n18079 = ~n18077 & ~n18078;
  assign n18080 = ~n16837 & ~n18079;
  assign n18081 = n16837 & n18079;
  assign n18082 = ~n18080 & ~n18081;
  assign n18083 = ~n18076 & ~n18082;
  assign n18084 = n18076 & n18082;
  assign n18085 = ~n14524 & n16839;
  assign n18086 = ~n14543 & ~n16855;
  assign n18087 = ~n18085 & ~n18086;
  assign n18088 = ~n16837 & ~n18087;
  assign n18089 = n16837 & n18087;
  assign n18090 = ~n18088 & ~n18089;
  assign n18091 = ~n14524 & ~n16846;
  assign n18092 = ~n14543 & n16839;
  assign n18093 = ~n18091 & ~n18092;
  assign n18094 = n18090 & n18093;
  assign n18095 = ~n18090 & ~n18093;
  assign n18096 = ~n14458 & ~n16846;
  assign n18097 = ~n14477 & n16839;
  assign n18098 = ~n18096 & ~n18097;
  assign n18099 = ~n14458 & n16839;
  assign n18100 = ~n14477 & ~n16855;
  assign n18101 = ~n18099 & ~n18100;
  assign n18102 = ~n16837 & ~n18101;
  assign n18103 = n16837 & n18101;
  assign n18104 = ~n18102 & ~n18103;
  assign n18105 = ~n18098 & ~n18104;
  assign n18106 = ~n18095 & ~n18105;
  assign n18107 = ~n14348 & ~n16846;
  assign n18108 = ~n14407 & n16839;
  assign n18109 = ~n18107 & ~n18108;
  assign n18110 = ~n14348 & n16839;
  assign n18111 = ~n14407 & ~n16855;
  assign n18112 = ~n18110 & ~n18111;
  assign n18113 = ~n16837 & ~n18112;
  assign n18114 = n16837 & n18112;
  assign n18115 = ~n18113 & ~n18114;
  assign n18116 = ~n18109 & ~n18115;
  assign n18117 = n18098 & n18104;
  assign n18118 = ~n18094 & ~n18117;
  assign n18119 = n18116 & n18118;
  assign n18120 = n18106 & ~n18119;
  assign n18121 = ~n18094 & ~n18120;
  assign n18122 = n18109 & n18115;
  assign n18123 = n18118 & ~n18122;
  assign n18124 = ~n14292 & ~n16846;
  assign n18125 = ~n14355 & n16839;
  assign n18126 = ~n18124 & ~n18125;
  assign n18127 = ~n14292 & n16839;
  assign n18128 = ~n14355 & ~n16855;
  assign n18129 = ~n18127 & ~n18128;
  assign n18130 = ~n16837 & ~n18129;
  assign n18131 = n16837 & n18129;
  assign n18132 = ~n18130 & ~n18131;
  assign n18133 = ~n18126 & ~n18132;
  assign n18134 = n18126 & n18132;
  assign n18135 = ~n14224 & ~n16846;
  assign n18136 = ~n14276_1 & n16839;
  assign n18137 = ~n18135 & ~n18136;
  assign n18138 = ~n14165 & ~n16846;
  assign n18139 = ~n14208 & n16839;
  assign n18140 = ~n18138 & ~n18139;
  assign n18141 = ~n14165 & n16839;
  assign n18142 = ~n14208 & ~n16855;
  assign n18143 = ~n18141 & ~n18142;
  assign n18144 = ~n16837 & ~n18143;
  assign n18145 = n16837 & n18143;
  assign n18146 = ~n18144 & ~n18145;
  assign n18147 = ~n18140 & ~n18146;
  assign n18148 = n18140 & n18146;
  assign n18149 = ~n14098 & ~n16846;
  assign n18150 = ~n14139 & n16839;
  assign n18151 = ~n18149 & ~n18150;
  assign n18152 = ~n14007 & ~n16846;
  assign n18153 = ~n14066_1 & n16839;
  assign n18154 = ~n18152 & ~n18153;
  assign n18155 = ~n14007 & n16839;
  assign n18156 = ~n14066_1 & ~n16855;
  assign n18157 = ~n18155 & ~n18156;
  assign n18158 = ~n16837 & ~n18157;
  assign n18159 = n16837 & n18157;
  assign n18160 = ~n18158 & ~n18159;
  assign n18161 = ~n18154 & ~n18160;
  assign n18162 = ~n18151 & n18161;
  assign n18163 = ~n14098 & n16839;
  assign n18164 = ~n14139 & ~n16855;
  assign n18165 = ~n18163 & ~n18164;
  assign n18166 = ~n16837 & ~n18165;
  assign n18167 = n16837 & n18165;
  assign n18168 = ~n18166 & ~n18167;
  assign n18169 = n18151 & ~n18161;
  assign n18170 = ~n18168 & ~n18169;
  assign n18171 = ~n18162 & ~n18170;
  assign n18172 = n18154 & n18160;
  assign n18173 = n18151 & n18168;
  assign n18174 = ~n18172 & ~n18173;
  assign n18175 = ~n13937 & ~n16846;
  assign n18176 = ~n14014 & n16839;
  assign n18177 = ~n18175 & ~n18176;
  assign n18178 = ~n13937 & n16839;
  assign n18179 = ~n14014 & ~n16855;
  assign n18180 = ~n18178 & ~n18179;
  assign n18181 = ~n16837 & ~n18180;
  assign n18182 = n16837 & n18180;
  assign n18183 = ~n18181 & ~n18182;
  assign n18184 = ~n18177 & ~n18183;
  assign n18185 = n18177 & n18183;
  assign n18186 = ~n13871_1 & ~n16846;
  assign n18187 = ~n13944 & n16839;
  assign n18188 = ~n18186 & ~n18187;
  assign n18189 = ~n13806_1 & ~n16846;
  assign n18190 = ~n13878 & n16839;
  assign n18191 = ~n18189 & ~n18190;
  assign n18192 = ~n13750 & ~n16846;
  assign n18193 = ~n13813 & n16839;
  assign n18194 = ~n18192 & ~n18193;
  assign n18195 = ~n13750 & n16839;
  assign n18196 = ~n13813 & ~n16855;
  assign n18197 = ~n18195 & ~n18196;
  assign n18198 = ~n16837 & ~n18197;
  assign n18199 = n16837 & n18197;
  assign n18200 = ~n18198 & ~n18199;
  assign n18201 = ~n18194 & ~n18200;
  assign n18202 = ~n18191 & n18201;
  assign n18203 = ~n13806_1 & n16839;
  assign n18204 = ~n13878 & ~n16855;
  assign n18205 = ~n18203 & ~n18204;
  assign n18206 = ~n16837 & ~n18205;
  assign n18207 = n16837 & n18205;
  assign n18208 = ~n18206 & ~n18207;
  assign n18209 = n18191 & ~n18201;
  assign n18210 = ~n18208 & ~n18209;
  assign n18211 = ~n18202 & ~n18210;
  assign n18212 = n18194 & n18200;
  assign n18213 = n18191 & n18208;
  assign n18214 = ~n18212 & ~n18213;
  assign n18215 = ~n13697 & ~n16846;
  assign n18216 = ~n13757 & n16839;
  assign n18217 = ~n18215 & ~n18216;
  assign n18218 = ~n13697 & n16839;
  assign n18219 = ~n13757 & ~n16855;
  assign n18220 = ~n18218 & ~n18219;
  assign n18221 = ~n16837 & ~n18220;
  assign n18222 = n16837 & n18220;
  assign n18223 = ~n18221 & ~n18222;
  assign n18224 = ~n18217 & ~n18223;
  assign n18225 = n18217 & n18223;
  assign n18226 = n16837 & ~n16848;
  assign n18227 = ~n16837 & n16848;
  assign n18228 = ~n16860 & ~n18227;
  assign n18229 = ~n18226 & ~n18228;
  assign n18230 = ~n18225 & ~n18229;
  assign n18231 = ~n18224 & ~n18230;
  assign n18232 = n18214 & ~n18231;
  assign n18233 = n18211 & ~n18232;
  assign n18234 = ~n18188 & ~n18233;
  assign n18235 = ~n13871_1 & n16839;
  assign n18236 = ~n13944 & ~n16855;
  assign n18237 = ~n18235 & ~n18236;
  assign n18238 = ~n16837 & ~n18237;
  assign n18239 = n16837 & n18237;
  assign n18240 = ~n18238 & ~n18239;
  assign n18241 = n18188 & n18233;
  assign n18242 = ~n18240 & ~n18241;
  assign n18243 = ~n18234 & ~n18242;
  assign n18244 = ~n18185 & ~n18243;
  assign n18245 = ~n18184 & ~n18244;
  assign n18246 = n18174 & ~n18245;
  assign n18247 = n18171 & ~n18246;
  assign n18248 = ~n18148 & ~n18247;
  assign n18249 = ~n18147 & ~n18248;
  assign n18250 = ~n18137 & ~n18249;
  assign n18251 = ~n14224 & n16839;
  assign n18252 = ~n14276_1 & ~n16855;
  assign n18253 = ~n18251 & ~n18252;
  assign n18254 = ~n16837 & ~n18253;
  assign n18255 = n16837 & n18253;
  assign n18256 = ~n18254 & ~n18255;
  assign n18257 = n18137 & n18249;
  assign n18258 = ~n18256 & ~n18257;
  assign n18259 = ~n18250 & ~n18258;
  assign n18260 = ~n18134 & ~n18259;
  assign n18261 = ~n18133 & ~n18260;
  assign n18262 = n18123 & ~n18261;
  assign n18263 = ~n18121 & ~n18262;
  assign n18264 = ~n18084 & ~n18263;
  assign n18265 = ~n18083 & ~n18264;
  assign n18266 = ~n14651_1 & n16839;
  assign n18267 = ~n14670 & ~n16855;
  assign n18268 = ~n18266 & ~n18267;
  assign n18269 = ~n16837 & ~n18268;
  assign n18270 = n16837 & n18268;
  assign n18271 = ~n18269 & ~n18270;
  assign n18272 = ~n14651_1 & ~n16846;
  assign n18273 = ~n14670 & n16839;
  assign n18274 = ~n18272 & ~n18273;
  assign n18275 = ~n18271 & n18274;
  assign n18276 = n18271 & ~n18274;
  assign n18277 = ~n18275 & ~n18276;
  assign n18278 = n18265 & ~n18277;
  assign n18279 = ~n18265 & n18277;
  assign n18280 = ~n18278 & ~n18279;
  assign n18281 = n13525 & ~n18055;
  assign n18282 = n18042 & n18281;
  assign n18283 = ~n18280 & n18282;
  assign n18284 = ~n18060 & ~n18064;
  assign n18285 = ~n16432 & n18284;
  assign n18286 = ~n18073 & n18285;
  assign n1866 = n18283 | ~n18286;
  assign n18288 = ~n15708 & ~n18042;
  assign n18289 = n18057 & ~n18288;
  assign n18290 = P3_STATE_REG & ~n18289;
  assign n18291 = ~n15320 & n18290;
  assign n18292 = ~n15708 & n18042;
  assign n18293 = ~n15698 & ~n18292;
  assign n18294 = n13525 & ~n18293;
  assign n18295 = n14988 & n18294;
  assign n18296 = P3_REG3_REG_26_ & ~P3_STATE_REG;
  assign n18297 = ~n15320 & ~n18042;
  assign n18298 = ~n15269 & n18067;
  assign n18299 = ~n15382 & n18069;
  assign n18300 = ~n18297 & ~n18298;
  assign n18301 = ~n18299 & n18300;
  assign n18302 = n18065 & ~n18301;
  assign n18303 = ~n15207 & ~n16846;
  assign n18304 = n14988 & n16839;
  assign n18305 = ~n18303 & ~n18304;
  assign n18306 = ~n15207 & n16839;
  assign n18307 = n14988 & ~n16855;
  assign n18308 = ~n18306 & ~n18307;
  assign n18309 = ~n16837 & ~n18308;
  assign n18310 = n16837 & n18308;
  assign n18311 = ~n18309 & ~n18310;
  assign n18312 = ~n18305 & ~n18311;
  assign n18313 = n18305 & n18311;
  assign n18314 = ~n15150 & ~n16846;
  assign n18315 = ~n18304 & ~n18314;
  assign n18316 = ~n15150 & n16839;
  assign n18317 = ~n18307 & ~n18316;
  assign n18318 = ~n16837 & ~n18317;
  assign n18319 = n16837 & n18317;
  assign n18320 = ~n18318 & ~n18319;
  assign n18321 = ~n18315 & ~n18320;
  assign n18322 = n18315 & n18320;
  assign n18323 = ~n15090 & ~n16846;
  assign n18324 = ~n18304 & ~n18323;
  assign n18325 = ~n15090 & n16839;
  assign n18326 = ~n18307 & ~n18325;
  assign n18327 = ~n16837 & ~n18326;
  assign n18328 = n16837 & n18326;
  assign n18329 = ~n18327 & ~n18328;
  assign n18330 = ~n18324 & ~n18329;
  assign n18331 = n18324 & n18329;
  assign n18332 = ~n14912 & n16839;
  assign n18333 = ~n14929 & ~n16855;
  assign n18334 = ~n18332 & ~n18333;
  assign n18335 = ~n16837 & ~n18334;
  assign n18336 = n16837 & n18334;
  assign n18337 = ~n18335 & ~n18336;
  assign n18338 = ~n14912 & ~n16846;
  assign n18339 = ~n14929 & n16839;
  assign n18340 = ~n18338 & ~n18339;
  assign n18341 = n18337 & n18340;
  assign n18342 = ~n14846_1 & ~n16846;
  assign n18343 = ~n14866_1 & n16839;
  assign n18344 = ~n18342 & ~n18343;
  assign n18345 = ~n14846_1 & n16839;
  assign n18346 = ~n14866_1 & ~n16855;
  assign n18347 = ~n18345 & ~n18346;
  assign n18348 = ~n16837 & ~n18347;
  assign n18349 = n16837 & n18347;
  assign n18350 = ~n18348 & ~n18349;
  assign n18351 = ~n18344 & ~n18350;
  assign n18352 = n18344 & n18350;
  assign n18353 = ~n14779 & ~n16846;
  assign n18354 = ~n14798 & n16839;
  assign n18355 = ~n18353 & ~n18354;
  assign n18356 = ~n14712 & ~n16846;
  assign n18357 = ~n14731_1 & n16839;
  assign n18358 = ~n18356 & ~n18357;
  assign n18359 = ~n14712 & n16839;
  assign n18360 = ~n14731_1 & ~n16855;
  assign n18361 = ~n18359 & ~n18360;
  assign n18362 = ~n16837 & ~n18361;
  assign n18363 = n16837 & n18361;
  assign n18364 = ~n18362 & ~n18363;
  assign n18365 = ~n18358 & ~n18364;
  assign n18366 = ~n18355 & n18365;
  assign n18367 = ~n14779 & n16839;
  assign n18368 = ~n14798 & ~n16855;
  assign n18369 = ~n18367 & ~n18368;
  assign n18370 = ~n16837 & ~n18369;
  assign n18371 = n16837 & n18369;
  assign n18372 = ~n18370 & ~n18371;
  assign n18373 = n18355 & ~n18365;
  assign n18374 = ~n18372 & ~n18373;
  assign n18375 = ~n18366 & ~n18374;
  assign n18376 = n18358 & n18364;
  assign n18377 = n18355 & n18372;
  assign n18378 = ~n18376 & ~n18377;
  assign n18379 = ~n18271 & ~n18274;
  assign n18380 = n18271 & n18274;
  assign n18381 = ~n18265 & ~n18380;
  assign n18382 = ~n18379 & ~n18381;
  assign n18383 = n18378 & ~n18382;
  assign n18384 = n18375 & ~n18383;
  assign n18385 = ~n18352 & ~n18384;
  assign n18386 = ~n18351 & ~n18385;
  assign n18387 = ~n14974 & n16839;
  assign n18388 = ~n18307 & ~n18387;
  assign n18389 = ~n16837 & ~n18388;
  assign n18390 = n16837 & n18388;
  assign n18391 = ~n18389 & ~n18390;
  assign n18392 = ~n14974 & ~n16846;
  assign n18393 = ~n18304 & ~n18392;
  assign n18394 = n18391 & n18393;
  assign n18395 = ~n15033 & n16839;
  assign n18396 = ~n18307 & ~n18395;
  assign n18397 = ~n16837 & ~n18396;
  assign n18398 = n16837 & n18396;
  assign n18399 = ~n18397 & ~n18398;
  assign n18400 = ~n15033 & ~n16846;
  assign n18401 = ~n18304 & ~n18400;
  assign n18402 = n18399 & n18401;
  assign n18403 = ~n18394 & ~n18402;
  assign n18404 = ~n18341 & ~n18386;
  assign n18405 = n18403 & n18404;
  assign n18406 = ~n18399 & ~n18401;
  assign n18407 = ~n18391 & ~n18393;
  assign n18408 = ~n18337 & ~n18340;
  assign n18409 = n18403 & n18408;
  assign n18410 = ~n18407 & ~n18409;
  assign n18411 = ~n18402 & ~n18410;
  assign n18412 = ~n18405 & ~n18406;
  assign n18413 = ~n18411 & n18412;
  assign n18414 = ~n18331 & ~n18413;
  assign n18415 = ~n18330 & ~n18414;
  assign n18416 = ~n18322 & ~n18415;
  assign n18417 = ~n18321 & ~n18416;
  assign n18418 = ~n18313 & ~n18417;
  assign n18419 = ~n18312 & ~n18418;
  assign n18420 = ~n15269 & ~n16846;
  assign n18421 = ~n18304 & ~n18420;
  assign n18422 = ~n15269 & n16839;
  assign n18423 = ~n18307 & ~n18422;
  assign n18424 = ~n16837 & ~n18423;
  assign n18425 = n16837 & n18423;
  assign n18426 = ~n18424 & ~n18425;
  assign n18427 = ~n18421 & ~n18426;
  assign n18428 = n18419 & ~n18427;
  assign n18429 = ~n15324 & ~n16846;
  assign n18430 = ~n18304 & ~n18429;
  assign n18431 = ~n15324 & n16839;
  assign n18432 = ~n18307 & ~n18431;
  assign n18433 = ~n16837 & ~n18432;
  assign n18434 = n16837 & n18432;
  assign n18435 = ~n18433 & ~n18434;
  assign n18436 = ~n18430 & ~n18435;
  assign n18437 = n18421 & n18426;
  assign n18438 = ~n18430 & ~n18437;
  assign n18439 = ~n18435 & ~n18437;
  assign n18440 = ~n18438 & ~n18439;
  assign n18441 = ~n18428 & ~n18436;
  assign n18442 = ~n18440 & n18441;
  assign n18443 = n18430 & ~n18435;
  assign n18444 = ~n18430 & n18435;
  assign n18445 = ~n18443 & ~n18444;
  assign n18446 = ~n18427 & n18445;
  assign n18447 = ~n18419 & ~n18437;
  assign n18448 = n18446 & ~n18447;
  assign n18449 = ~n18442 & ~n18448;
  assign n18450 = n18282 & n18449;
  assign n18451 = ~n18291 & ~n18295;
  assign n18452 = ~n18296 & n18451;
  assign n18453 = ~n18302 & n18452;
  assign n1871 = n18450 | ~n18453;
  assign n18455 = ~n14000 & ~n18059;
  assign n18456 = ~n14066_1 & ~n18063;
  assign n18457 = ~n14098 & n18069;
  assign n18458 = ~n13937 & n18067;
  assign n18459 = ~n14000 & ~n18042;
  assign n18460 = ~n18457 & ~n18458;
  assign n18461 = ~n18459 & n18460;
  assign n18462 = n18065 & ~n18461;
  assign n18463 = n18154 & ~n18160;
  assign n18464 = ~n18154 & n18160;
  assign n18465 = ~n18463 & ~n18464;
  assign n18466 = n18245 & ~n18465;
  assign n18467 = ~n18161 & ~n18172;
  assign n18468 = ~n18245 & ~n18467;
  assign n18469 = ~n18466 & ~n18468;
  assign n18470 = n18282 & ~n18469;
  assign n18471 = ~n18455 & ~n18456;
  assign n18472 = ~n16739 & n18471;
  assign n18473 = ~n18462 & n18472;
  assign n1876 = n18470 | ~n18473;
  assign n18475 = ~n14842 & ~n18059;
  assign n18476 = ~n14866_1 & ~n18063;
  assign n18477 = ~n14842 & ~n18042;
  assign n18478 = ~n14779 & n18067;
  assign n18479 = ~n14912 & n18069;
  assign n18480 = ~n18477 & ~n18478;
  assign n18481 = ~n18479 & n18480;
  assign n18482 = n18065 & ~n18481;
  assign n18483 = n18344 & ~n18350;
  assign n18484 = ~n18344 & n18350;
  assign n18485 = ~n18483 & ~n18484;
  assign n18486 = n18384 & ~n18485;
  assign n18487 = ~n18384 & n18485;
  assign n18488 = ~n18486 & ~n18487;
  assign n18489 = n18282 & ~n18488;
  assign n18490 = ~n18475 & ~n18476;
  assign n18491 = ~n16336_1 & n18490;
  assign n18492 = ~n18482 & n18491;
  assign n1881 = n18489 | ~n18492;
  assign n18494 = n18194 & ~n18200;
  assign n18495 = ~n18194 & n18200;
  assign n18496 = ~n18494 & ~n18495;
  assign n18497 = n18231 & ~n18496;
  assign n18498 = ~n18201 & ~n18212;
  assign n18499 = ~n18231 & ~n18498;
  assign n18500 = ~n18497 & ~n18499;
  assign n18501 = n18282 & ~n18500;
  assign n18502 = ~n16920 & ~n18501;
  assign n18503 = ~n13813 & ~n18063;
  assign n18504 = n18502 & ~n18503;
  assign n18505 = P3_REG3_REG_2_ & ~n18059;
  assign n18506 = ~n13806_1 & n18069;
  assign n18507 = ~n13697 & n18067;
  assign n18508 = P3_REG3_REG_2_ & ~n18042;
  assign n18509 = ~n18506 & ~n18507;
  assign n18510 = ~n18508 & n18509;
  assign n18511 = n18065 & ~n18510;
  assign n18512 = n18504 & ~n18505;
  assign n1886 = n18511 | ~n18512;
  assign n18514 = ~n14344 & ~n18059;
  assign n18515 = ~n14407 & ~n18063;
  assign n18516 = ~n14458 & n18069;
  assign n18517 = ~n14292 & n18067;
  assign n18518 = ~n14344 & ~n18042;
  assign n18519 = ~n18516 & ~n18517;
  assign n18520 = ~n18518 & n18519;
  assign n18521 = n18065 & ~n18520;
  assign n18522 = n18109 & ~n18115;
  assign n18523 = ~n18109 & n18115;
  assign n18524 = ~n18522 & ~n18523;
  assign n18525 = n18261 & ~n18524;
  assign n18526 = ~n18116 & ~n18122;
  assign n18527 = ~n18261 & ~n18526;
  assign n18528 = ~n18525 & ~n18527;
  assign n18529 = n18282 & ~n18528;
  assign n18530 = ~n18514 & ~n18515;
  assign n18531 = ~n16559 & n18530;
  assign n18532 = ~n18521 & n18531;
  assign n1891 = n18529 | ~n18532;
  assign n18534 = ~n15086_1 & n18290;
  assign n18535 = P3_REG3_REG_22_ & ~P3_STATE_REG;
  assign n18536 = ~n15086_1 & ~n18042;
  assign n18537 = ~n15033 & n18067;
  assign n18538 = ~n15150 & n18069;
  assign n18539 = ~n18536 & ~n18537;
  assign n18540 = ~n18538 & n18539;
  assign n18541 = n18065 & ~n18540;
  assign n18542 = n18324 & ~n18329;
  assign n18543 = ~n18324 & n18329;
  assign n18544 = ~n18542 & ~n18543;
  assign n18545 = n18413 & ~n18544;
  assign n18546 = ~n18413 & n18544;
  assign n18547 = ~n18545 & ~n18546;
  assign n18548 = n18282 & ~n18547;
  assign n18549 = ~n18295 & ~n18534;
  assign n18550 = ~n18535 & n18549;
  assign n18551 = ~n18541 & n18550;
  assign n1896 = n18548 | ~n18551;
  assign n18553 = ~n14520 & ~n18059;
  assign n18554 = ~n14543 & ~n18063;
  assign n18555 = ~n14520 & ~n18042;
  assign n18556 = ~n14458 & n18067;
  assign n18557 = ~n14588 & n18069;
  assign n18558 = ~n18555 & ~n18556;
  assign n18559 = ~n18557 & n18558;
  assign n18560 = n18065 & ~n18559;
  assign n18561 = ~n18095 & n18118;
  assign n18562 = ~n18122 & ~n18261;
  assign n18563 = ~n18116 & ~n18562;
  assign n18564 = ~n18105 & n18563;
  assign n18565 = n18561 & ~n18564;
  assign n18566 = ~n18090 & n18093;
  assign n18567 = n18090 & ~n18093;
  assign n18568 = ~n18566 & ~n18567;
  assign n18569 = ~n18105 & n18568;
  assign n18570 = ~n18117 & ~n18563;
  assign n18571 = n18569 & ~n18570;
  assign n18572 = ~n18565 & ~n18571;
  assign n18573 = n18282 & n18572;
  assign n18574 = ~n18553 & ~n18554;
  assign n18575 = ~n16494 & n18574;
  assign n18576 = ~n18560 & n18575;
  assign n1901 = n18573 | ~n18576;
  assign n18578 = ~n14970 & n18290;
  assign n18579 = P3_REG3_REG_20_ & ~P3_STATE_REG;
  assign n18580 = ~n14970 & ~n18042;
  assign n18581 = ~n14912 & n18067;
  assign n18582 = ~n15033 & n18069;
  assign n18583 = ~n18580 & ~n18581;
  assign n18584 = ~n18582 & n18583;
  assign n18585 = n18065 & ~n18584;
  assign n18586 = ~n18391 & n18393;
  assign n18587 = n18391 & ~n18393;
  assign n18588 = ~n18586 & ~n18587;
  assign n18589 = ~n18404 & ~n18408;
  assign n18590 = ~n18588 & n18589;
  assign n18591 = ~n18394 & ~n18407;
  assign n18592 = ~n18589 & ~n18591;
  assign n18593 = ~n18590 & ~n18592;
  assign n18594 = n18282 & ~n18593;
  assign n18595 = ~n18295 & ~n18578;
  assign n18596 = ~n18579 & n18595;
  assign n18597 = ~n18585 & n18596;
  assign n1906 = n18594 | ~n18597;
  assign n18599 = ~n16863 & n18282;
  assign n18600 = ~n16975 & ~n18599;
  assign n18601 = ~n18040 & ~n18065;
  assign n18602 = ~n18042 & ~n18601;
  assign n18603 = ~n18058 & ~n18602;
  assign n18604 = P3_REG3_REG_0_ & ~n18603;
  assign n18605 = ~n13671_1 & ~n18063;
  assign n18606 = ~n13697 & n18065;
  assign n18607 = n18069 & n18606;
  assign n18608 = ~n18605 & ~n18607;
  assign n18609 = n18600 & ~n18604;
  assign n1911 = ~n18608 | ~n18609;
  assign n18611 = ~n14220 & ~n18059;
  assign n18612 = ~n14276_1 & ~n18063;
  assign n18613 = ~n14292 & n18069;
  assign n18614 = ~n14165 & n18067;
  assign n18615 = ~n14220 & ~n18042;
  assign n18616 = ~n18613 & ~n18614;
  assign n18617 = ~n18615 & n18616;
  assign n18618 = n18065 & ~n18617;
  assign n18619 = n18137 & ~n18256;
  assign n18620 = ~n18137 & n18256;
  assign n18621 = ~n18619 & ~n18620;
  assign n18622 = n18249 & ~n18621;
  assign n18623 = ~n18249 & n18621;
  assign n18624 = ~n18622 & ~n18623;
  assign n18625 = n18282 & ~n18624;
  assign n18626 = ~n18611 & ~n18612;
  assign n18627 = ~n16629 & n18626;
  assign n18628 = ~n18618 & n18627;
  assign n1916 = n18625 | ~n18628;
  assign n18630 = n18188 & ~n18240;
  assign n18631 = ~n18188 & n18240;
  assign n18632 = ~n18630 & ~n18631;
  assign n18633 = n18233 & ~n18632;
  assign n18634 = ~n18233 & n18632;
  assign n18635 = ~n18633 & ~n18634;
  assign n18636 = n18282 & ~n18635;
  assign n18637 = ~n16811 & ~n18636;
  assign n18638 = ~n13944 & ~n18063;
  assign n18639 = n18637 & ~n18638;
  assign n18640 = ~n13864 & ~n18059;
  assign n18641 = ~n13937 & n18069;
  assign n18642 = ~n13806_1 & n18067;
  assign n18643 = ~n13864 & ~n18042;
  assign n18644 = ~n18641 & ~n18642;
  assign n18645 = ~n18643 & n18644;
  assign n18646 = n18065 & ~n18645;
  assign n18647 = n18639 & ~n18640;
  assign n1921 = n18646 | ~n18647;
  assign n18649 = ~n15203 & n18290;
  assign n18650 = P3_REG3_REG_24_ & ~P3_STATE_REG;
  assign n18651 = ~n15203 & ~n18042;
  assign n18652 = ~n15150 & n18067;
  assign n18653 = ~n15269 & n18069;
  assign n18654 = ~n18651 & ~n18652;
  assign n18655 = ~n18653 & n18654;
  assign n18656 = n18065 & ~n18655;
  assign n18657 = n18305 & ~n18311;
  assign n18658 = ~n18305 & n18311;
  assign n18659 = ~n18657 & ~n18658;
  assign n18660 = n18417 & ~n18659;
  assign n18661 = ~n18312 & ~n18313;
  assign n18662 = ~n18417 & ~n18661;
  assign n18663 = ~n18660 & ~n18662;
  assign n18664 = n18282 & ~n18663;
  assign n18665 = ~n18295 & ~n18649;
  assign n18666 = ~n18650 & n18665;
  assign n18667 = ~n18656 & n18666;
  assign n1926 = n18664 | ~n18667;
  assign n18669 = ~n14775 & ~n18059;
  assign n18670 = ~n14798 & ~n18063;
  assign n18671 = ~n14775 & ~n18042;
  assign n18672 = ~n14712 & n18067;
  assign n18673 = ~n14846_1 & n18069;
  assign n18674 = ~n18671 & ~n18672;
  assign n18675 = ~n18673 & n18674;
  assign n18676 = n18065 & ~n18675;
  assign n18677 = ~n18355 & ~n18372;
  assign n18678 = n18378 & ~n18677;
  assign n18679 = ~n18365 & n18382;
  assign n18680 = n18678 & ~n18679;
  assign n18681 = n18355 & ~n18372;
  assign n18682 = ~n18355 & n18372;
  assign n18683 = ~n18681 & ~n18682;
  assign n18684 = ~n18365 & n18683;
  assign n18685 = ~n18376 & ~n18382;
  assign n18686 = n18684 & ~n18685;
  assign n18687 = ~n18680 & ~n18686;
  assign n18688 = n18282 & n18687;
  assign n18689 = ~n18669 & ~n18670;
  assign n18690 = ~n16369 & n18689;
  assign n18691 = ~n18676 & n18690;
  assign n1931 = n18688 | ~n18691;
  assign n18693 = ~n13930 & ~n18059;
  assign n18694 = ~n14014 & ~n18063;
  assign n18695 = ~n14007 & n18069;
  assign n18696 = ~n13871_1 & n18067;
  assign n18697 = ~n13930 & ~n18042;
  assign n18698 = ~n18695 & ~n18696;
  assign n18699 = ~n18697 & n18698;
  assign n18700 = n18065 & ~n18699;
  assign n18701 = n18177 & ~n18183;
  assign n18702 = ~n18177 & n18183;
  assign n18703 = ~n18701 & ~n18702;
  assign n18704 = n18243 & ~n18703;
  assign n18705 = ~n18243 & n18703;
  assign n18706 = ~n18704 & ~n18705;
  assign n18707 = n18282 & ~n18706;
  assign n18708 = ~n16789 & ~n18707;
  assign n18709 = ~n18693 & ~n18694;
  assign n18710 = ~n18700 & n18709;
  assign n1936 = ~n18708 | ~n18710;
  assign n18712 = ~n14708 & ~n18059;
  assign n18713 = ~n14731_1 & ~n18063;
  assign n18714 = ~n14708 & ~n18042;
  assign n18715 = ~n14651_1 & n18067;
  assign n18716 = ~n14779 & n18069;
  assign n18717 = ~n18714 & ~n18715;
  assign n18718 = ~n18716 & n18717;
  assign n18719 = n18065 & ~n18718;
  assign n18720 = n18358 & ~n18364;
  assign n18721 = ~n18358 & n18364;
  assign n18722 = ~n18720 & ~n18721;
  assign n18723 = n18382 & ~n18722;
  assign n18724 = ~n18365 & ~n18376;
  assign n18725 = ~n18382 & ~n18724;
  assign n18726 = ~n18723 & ~n18725;
  assign n18727 = n18282 & ~n18726;
  assign n18728 = ~n18712 & ~n18713;
  assign n18729 = ~n16403 & n18728;
  assign n18730 = ~n18719 & n18729;
  assign n1941 = n18727 | ~n18730;
  assign n18732 = ~n15265 & n18290;
  assign n18733 = P3_REG3_REG_25_ & ~P3_STATE_REG;
  assign n18734 = ~n15265 & ~n18042;
  assign n18735 = ~n15207 & n18067;
  assign n18736 = ~n15324 & n18069;
  assign n18737 = ~n18734 & ~n18735;
  assign n18738 = ~n18736 & n18737;
  assign n18739 = n18065 & ~n18738;
  assign n18740 = n18421 & ~n18426;
  assign n18741 = ~n18421 & n18426;
  assign n18742 = ~n18740 & ~n18741;
  assign n18743 = n18419 & ~n18742;
  assign n18744 = ~n18427 & ~n18437;
  assign n18745 = ~n18419 & ~n18744;
  assign n18746 = ~n18743 & ~n18745;
  assign n18747 = n18282 & ~n18746;
  assign n18748 = ~n18295 & ~n18732;
  assign n18749 = ~n18733 & n18748;
  assign n18750 = ~n18739 & n18749;
  assign n1946 = n18747 | ~n18750;
  assign n18752 = ~n14454 & ~n18059;
  assign n18753 = ~n14477 & ~n18063;
  assign n18754 = ~n14454 & ~n18042;
  assign n18755 = ~n14348 & n18067;
  assign n18756 = ~n14524 & n18069;
  assign n18757 = ~n18754 & ~n18755;
  assign n18758 = ~n18756 & n18757;
  assign n18759 = n18065 & ~n18758;
  assign n18760 = n18098 & ~n18104;
  assign n18761 = ~n18098 & n18104;
  assign n18762 = ~n18760 & ~n18761;
  assign n18763 = n18563 & ~n18762;
  assign n18764 = ~n18105 & ~n18117;
  assign n18765 = ~n18563 & ~n18764;
  assign n18766 = ~n18763 & ~n18765;
  assign n18767 = n18282 & ~n18766;
  assign n18768 = ~n18752 & ~n18753;
  assign n18769 = ~n16529 & n18768;
  assign n18770 = ~n18759 & n18769;
  assign n1951 = n18767 | ~n18770;
  assign n18772 = ~n15029 & n18290;
  assign n18773 = P3_REG3_REG_21_ & ~P3_STATE_REG;
  assign n18774 = ~n15029 & ~n18042;
  assign n18775 = ~n14974 & n18067;
  assign n18776 = ~n15090 & n18069;
  assign n18777 = ~n18774 & ~n18775;
  assign n18778 = ~n18776 & n18777;
  assign n18779 = n18065 & ~n18778;
  assign n18780 = ~n18407 & n18589;
  assign n18781 = ~n18406 & ~n18780;
  assign n18782 = n18403 & n18781;
  assign n18783 = ~n18399 & n18401;
  assign n18784 = n18399 & ~n18401;
  assign n18785 = ~n18783 & ~n18784;
  assign n18786 = ~n18407 & n18785;
  assign n18787 = ~n18394 & ~n18589;
  assign n18788 = n18786 & ~n18787;
  assign n18789 = ~n18782 & ~n18788;
  assign n18790 = n18282 & n18789;
  assign n18791 = ~n18295 & ~n18772;
  assign n18792 = ~n18773 & n18791;
  assign n18793 = ~n18779 & n18792;
  assign n1956 = n18790 | ~n18793;
  assign n18795 = n18217 & ~n18223;
  assign n18796 = ~n18217 & n18223;
  assign n18797 = ~n18795 & ~n18796;
  assign n18798 = n18229 & ~n18797;
  assign n18799 = ~n18229 & n18797;
  assign n18800 = ~n18798 & ~n18799;
  assign n18801 = n18282 & ~n18800;
  assign n18802 = ~n16953 & ~n18801;
  assign n18803 = ~n13757 & ~n18063;
  assign n18804 = n18802 & ~n18803;
  assign n18805 = P3_REG3_REG_1_ & ~n18059;
  assign n18806 = ~n13750 & n18069;
  assign n18807 = ~n13707 & n18067;
  assign n18808 = P3_REG3_REG_1_ & ~n18042;
  assign n18809 = ~n18806 & ~n18807;
  assign n18810 = ~n18808 & n18809;
  assign n18811 = n18065 & ~n18810;
  assign n18812 = n18804 & ~n18805;
  assign n1961 = n18811 | ~n18812;
  assign n18814 = ~n14158 & ~n18059;
  assign n18815 = ~n14208 & ~n18063;
  assign n18816 = ~n14224 & n18069;
  assign n18817 = ~n14098 & n18067;
  assign n18818 = ~n14158 & ~n18042;
  assign n18819 = ~n18816 & ~n18817;
  assign n18820 = ~n18818 & n18819;
  assign n18821 = n18065 & ~n18820;
  assign n18822 = n18140 & ~n18146;
  assign n18823 = ~n18140 & n18146;
  assign n18824 = ~n18822 & ~n18823;
  assign n18825 = n18247 & ~n18824;
  assign n18826 = ~n18247 & n18824;
  assign n18827 = ~n18825 & ~n18826;
  assign n18828 = n18282 & ~n18827;
  assign n18829 = ~n18814 & ~n18815;
  assign n18830 = ~n16659 & n18829;
  assign n18831 = ~n18821 & n18830;
  assign n1966 = n18828 | ~n18831;
  assign n18833 = ~n15435 & n18290;
  assign n18834 = P3_REG3_REG_28_ & ~P3_STATE_REG;
  assign n18835 = ~n15501_1 & n18069;
  assign n18836 = ~n15382 & n18067;
  assign n18837 = ~n15435 & ~n18042;
  assign n18838 = ~n18835 & ~n18836;
  assign n18839 = ~n18837 & n18838;
  assign n18840 = n18065 & ~n18839;
  assign n18841 = ~n15382 & n16839;
  assign n18842 = ~n18307 & ~n18841;
  assign n18843 = ~n16837 & ~n18842;
  assign n18844 = n16837 & n18842;
  assign n18845 = ~n18843 & ~n18844;
  assign n18846 = ~n15382 & ~n16846;
  assign n18847 = ~n18304 & ~n18846;
  assign n18848 = n18845 & n18847;
  assign n18849 = n18436 & ~n18848;
  assign n18850 = ~n18313 & ~n18848;
  assign n18851 = ~n18417 & ~n18440;
  assign n18852 = n18850 & n18851;
  assign n18853 = ~n18312 & ~n18427;
  assign n18854 = ~n18440 & ~n18853;
  assign n18855 = ~n18848 & n18854;
  assign n18856 = ~n18845 & ~n18847;
  assign n18857 = ~n18855 & ~n18856;
  assign n18858 = ~n15439 & ~n16846;
  assign n18859 = ~n18304 & ~n18858;
  assign n18860 = ~n16837 & ~n18859;
  assign n18861 = n16837 & n18859;
  assign n18862 = ~n18860 & ~n18861;
  assign n18863 = ~n15439 & n16839;
  assign n18864 = ~n18307 & ~n18863;
  assign n18865 = ~n18862 & n18864;
  assign n18866 = n18862 & ~n18864;
  assign n18867 = ~n18865 & ~n18866;
  assign n18868 = ~n18849 & ~n18852;
  assign n18869 = n18857 & n18868;
  assign n18870 = ~n18867 & n18869;
  assign n18871 = n18418 & ~n18440;
  assign n18872 = ~n18436 & ~n18856;
  assign n18873 = ~n18854 & ~n18871;
  assign n18874 = n18872 & n18873;
  assign n18875 = ~n18848 & ~n18874;
  assign n18876 = n18867 & n18875;
  assign n18877 = ~n18870 & ~n18876;
  assign n18878 = n18282 & ~n18877;
  assign n18879 = ~n18295 & ~n18833;
  assign n18880 = ~n18834 & n18879;
  assign n18881 = ~n18840 & n18880;
  assign n1971 = n18878 | ~n18881;
  assign n18883 = ~n14908 & ~n18059;
  assign n18884 = ~n14929 & ~n18063;
  assign n18885 = ~n14908 & ~n18042;
  assign n18886 = ~n14846_1 & n18067;
  assign n18887 = ~n14974 & n18069;
  assign n18888 = ~n18885 & ~n18886;
  assign n18889 = ~n18887 & n18888;
  assign n18890 = n18065 & ~n18889;
  assign n18891 = ~n18337 & n18340;
  assign n18892 = n18337 & ~n18340;
  assign n18893 = ~n18891 & ~n18892;
  assign n18894 = n18386 & ~n18893;
  assign n18895 = ~n18341 & ~n18408;
  assign n18896 = ~n18386 & ~n18895;
  assign n18897 = ~n18894 & ~n18896;
  assign n18898 = n18282 & ~n18897;
  assign n18899 = ~n18883 & ~n18884;
  assign n18900 = ~n16206_1 & n18899;
  assign n18901 = ~n18890 & n18900;
  assign n1976 = n18898 | ~n18901;
  assign n18903 = ~n18191 & ~n18208;
  assign n18904 = n18214 & ~n18903;
  assign n18905 = ~n18201 & n18231;
  assign n18906 = n18904 & ~n18905;
  assign n18907 = n18191 & ~n18208;
  assign n18908 = ~n18191 & n18208;
  assign n18909 = ~n18907 & ~n18908;
  assign n18910 = ~n18201 & n18909;
  assign n18911 = ~n18212 & ~n18231;
  assign n18912 = n18910 & ~n18911;
  assign n18913 = ~n18906 & ~n18912;
  assign n18914 = n18282 & n18913;
  assign n18915 = ~n16897 & ~n18914;
  assign n18916 = ~n13878 & ~n18063;
  assign n18917 = n18915 & ~n18916;
  assign n18918 = ~P3_REG3_REG_3_ & ~n18059;
  assign n18919 = ~n13871_1 & n18069;
  assign n18920 = ~n13750 & n18067;
  assign n18921 = ~P3_REG3_REG_3_ & ~n18042;
  assign n18922 = ~n18919 & ~n18920;
  assign n18923 = ~n18921 & n18922;
  assign n18924 = n18065 & ~n18923;
  assign n18925 = n18917 & ~n18918;
  assign n1981 = n18924 | ~n18925;
  assign n18927 = ~n14288 & ~n18059;
  assign n18928 = ~n14355 & ~n18063;
  assign n18929 = ~n14348 & n18069;
  assign n18930 = ~n14224 & n18067;
  assign n18931 = ~n14288 & ~n18042;
  assign n18932 = ~n18929 & ~n18930;
  assign n18933 = ~n18931 & n18932;
  assign n18934 = n18065 & ~n18933;
  assign n18935 = n18126 & ~n18132;
  assign n18936 = ~n18126 & n18132;
  assign n18937 = ~n18935 & ~n18936;
  assign n18938 = n18259 & ~n18937;
  assign n18939 = ~n18259 & n18937;
  assign n18940 = ~n18938 & ~n18939;
  assign n18941 = n18282 & ~n18940;
  assign n18942 = ~n18927 & ~n18928;
  assign n18943 = ~n16594 & n18942;
  assign n18944 = ~n18934 & n18943;
  assign n1986 = n18941 | ~n18944;
  assign n18946 = ~n15146_1 & n18290;
  assign n18947 = P3_REG3_REG_23_ & ~P3_STATE_REG;
  assign n18948 = ~n15146_1 & ~n18042;
  assign n18949 = ~n15090 & n18067;
  assign n18950 = ~n15207 & n18069;
  assign n18951 = ~n18948 & ~n18949;
  assign n18952 = ~n18950 & n18951;
  assign n18953 = n18065 & ~n18952;
  assign n18954 = n18315 & ~n18320;
  assign n18955 = ~n18315 & n18320;
  assign n18956 = ~n18954 & ~n18955;
  assign n18957 = n18415 & ~n18956;
  assign n18958 = ~n18415 & n18956;
  assign n18959 = ~n18957 & ~n18958;
  assign n18960 = n18282 & ~n18959;
  assign n18961 = ~n18295 & ~n18946;
  assign n18962 = ~n18947 & n18961;
  assign n18963 = ~n18953 & n18962;
  assign n1991 = n18960 | ~n18963;
  assign n18965 = ~n14584 & ~n18059;
  assign n18966 = ~n14609 & ~n18063;
  assign n18967 = ~n14584 & ~n18042;
  assign n18968 = ~n14524 & n18067;
  assign n18969 = ~n14651_1 & n18069;
  assign n18970 = ~n18967 & ~n18968;
  assign n18971 = ~n18969 & n18970;
  assign n18972 = n18065 & ~n18971;
  assign n18973 = n18076 & ~n18082;
  assign n18974 = ~n18076 & n18082;
  assign n18975 = ~n18973 & ~n18974;
  assign n18976 = n18263 & ~n18975;
  assign n18977 = ~n18263 & n18975;
  assign n18978 = ~n18976 & ~n18977;
  assign n18979 = n18282 & ~n18978;
  assign n18980 = ~n18965 & ~n18966;
  assign n18981 = ~n16460 & n18980;
  assign n18982 = ~n18972 & n18981;
  assign n1996 = n18979 | ~n18982;
  assign n18984 = ~n15378 & n18290;
  assign n18985 = P3_REG3_REG_27_ & ~P3_STATE_REG;
  assign n18986 = ~n15378 & ~n18042;
  assign n18987 = ~n15324 & n18067;
  assign n18988 = ~n15439 & n18069;
  assign n18989 = ~n18986 & ~n18987;
  assign n18990 = ~n18988 & n18989;
  assign n18991 = n18065 & ~n18990;
  assign n18992 = ~n18436 & n18873;
  assign n18993 = ~n18845 & n18847;
  assign n18994 = n18845 & ~n18847;
  assign n18995 = ~n18993 & ~n18994;
  assign n18996 = n18992 & ~n18995;
  assign n18997 = ~n18992 & n18995;
  assign n18998 = ~n18996 & ~n18997;
  assign n18999 = n18282 & ~n18998;
  assign n19000 = ~n18295 & ~n18984;
  assign n19001 = ~n18985 & n19000;
  assign n19002 = ~n18991 & n19001;
  assign n2001 = n18999 | ~n19002;
  assign n19004 = ~n14091_1 & ~n18059;
  assign n19005 = ~n14139 & ~n18063;
  assign n19006 = ~n14165 & n18069;
  assign n19007 = ~n14007 & n18067;
  assign n19008 = ~n14091_1 & ~n18042;
  assign n19009 = ~n19006 & ~n19007;
  assign n19010 = ~n19008 & n19009;
  assign n19011 = n18065 & ~n19010;
  assign n19012 = ~n18151 & ~n18168;
  assign n19013 = n18174 & ~n19012;
  assign n19014 = ~n18161 & n18245;
  assign n19015 = n19013 & ~n19014;
  assign n19016 = n18151 & ~n18168;
  assign n19017 = ~n18151 & n18168;
  assign n19018 = ~n19016 & ~n19017;
  assign n19019 = ~n18161 & n19018;
  assign n19020 = ~n18172 & ~n18245;
  assign n19021 = n19019 & ~n19020;
  assign n19022 = ~n19015 & ~n19021;
  assign n19023 = n18282 & n19022;
  assign n19024 = ~n19004 & ~n19005;
  assign n19025 = ~n16693 & n19024;
  assign n19026 = ~n19011 & n19025;
  assign n2006 = n19023 | ~n19026;
  assign n19028 = ~P4_IR_REG_31_ & P4_STATE_REG;
  assign n19029 = P4_IR_REG_0_ & n19028;
  assign n19030 = ~P4_STATE_REG & P2_P3_DATAO_REG_0_;
  assign n19031 = ~n19029 & ~n19030;
  assign n19032 = P4_STATE_REG & ~n19028;
  assign n19033 = P4_IR_REG_0_ & n19032;
  assign n2026 = ~n19031 | n19033;
  assign n19035 = P4_IR_REG_1_ & n19028;
  assign n19036 = ~P4_STATE_REG & P2_P3_DATAO_REG_1_;
  assign n19037 = ~n19035 & ~n19036;
  assign n19038 = P4_IR_REG_0_ & ~P4_IR_REG_1_;
  assign n19039 = ~P4_IR_REG_0_ & P4_IR_REG_1_;
  assign n19040 = ~n19038 & ~n19039;
  assign n19041 = n19032 & ~n19040;
  assign n2031 = ~n19037 | n19041;
  assign n19043 = P4_IR_REG_2_ & n19028;
  assign n19044 = ~P4_STATE_REG & P2_P3_DATAO_REG_2_;
  assign n19045 = ~n19043 & ~n19044;
  assign n19046 = ~P4_IR_REG_0_ & ~P4_IR_REG_1_;
  assign n19047 = P4_IR_REG_2_ & ~n19046;
  assign n19048 = ~P4_IR_REG_2_ & n19046;
  assign n19049 = ~n19047 & ~n19048;
  assign n19050 = n19032 & n19049;
  assign n2036 = ~n19045 | n19050;
  assign n19052 = P4_IR_REG_3_ & n19028;
  assign n19053 = ~P4_STATE_REG & P2_P3_DATAO_REG_3_;
  assign n19054 = ~n19052 & ~n19053;
  assign n19055 = P4_IR_REG_3_ & ~n19048;
  assign n19056 = ~P4_IR_REG_3_ & n19048;
  assign n19057 = ~n19055 & ~n19056;
  assign n19058 = n19032 & n19057;
  assign n2041 = ~n19054 | n19058;
  assign n19060 = P4_IR_REG_4_ & n19028;
  assign n19061 = ~P4_STATE_REG & P2_P3_DATAO_REG_4_;
  assign n19062 = ~n19060 & ~n19061;
  assign n19063 = P4_IR_REG_4_ & ~n19056;
  assign n19064 = ~P4_IR_REG_3_ & ~P4_IR_REG_4_;
  assign n19065 = n19048 & n19064;
  assign n19066 = ~n19063 & ~n19065;
  assign n19067 = n19032 & n19066;
  assign n2046 = ~n19062 | n19067;
  assign n19069 = P4_IR_REG_5_ & n19028;
  assign n19070 = ~P4_STATE_REG & P2_P3_DATAO_REG_5_;
  assign n19071 = ~n19069 & ~n19070;
  assign n19072 = ~P4_IR_REG_5_ & n19065;
  assign n19073 = P4_IR_REG_5_ & ~n19065;
  assign n19074 = ~n19072 & ~n19073;
  assign n19075 = n19032 & n19074;
  assign n2051 = ~n19071 | n19075;
  assign n19077 = P4_IR_REG_6_ & n19028;
  assign n19078 = ~P4_STATE_REG & P2_P3_DATAO_REG_6_;
  assign n19079 = ~n19077 & ~n19078;
  assign n19080 = P4_IR_REG_6_ & ~n19072;
  assign n19081 = ~P4_IR_REG_5_ & ~P4_IR_REG_6_;
  assign n19082 = n19065 & n19081;
  assign n19083 = ~n19080 & ~n19082;
  assign n19084 = n19032 & n19083;
  assign n2056 = ~n19079 | n19084;
  assign n19086 = P4_IR_REG_7_ & n19028;
  assign n19087 = ~P4_STATE_REG & P2_P3_DATAO_REG_7_;
  assign n19088 = ~n19086 & ~n19087;
  assign n19089 = P4_IR_REG_7_ & ~n19082;
  assign n19090 = ~P4_IR_REG_7_ & n19082;
  assign n19091 = ~n19089 & ~n19090;
  assign n19092 = n19032 & n19091;
  assign n2061 = ~n19088 | n19092;
  assign n19094 = P4_IR_REG_8_ & n19028;
  assign n19095 = ~P4_STATE_REG & P2_P3_DATAO_REG_8_;
  assign n19096 = ~n19094 & ~n19095;
  assign n19097 = P4_IR_REG_8_ & ~n19090;
  assign n19098 = ~P4_IR_REG_7_ & ~P4_IR_REG_8_;
  assign n19099 = ~P4_IR_REG_5_ & n19064;
  assign n19100 = ~P4_IR_REG_6_ & n19099;
  assign n19101 = n19048 & n19098;
  assign n19102 = n19100 & n19101;
  assign n19103 = ~n19097 & ~n19102;
  assign n19104 = n19032 & n19103;
  assign n2066 = ~n19096 | n19104;
  assign n19106 = P4_IR_REG_9_ & n19028;
  assign n19107 = ~P4_STATE_REG & P2_P3_DATAO_REG_9_;
  assign n19108 = ~n19106 & ~n19107;
  assign n19109 = ~P4_IR_REG_9_ & n19102;
  assign n19110 = P4_IR_REG_9_ & ~n19102;
  assign n19111 = ~n19109 & ~n19110;
  assign n19112 = n19032 & n19111;
  assign n2071 = ~n19108 | n19112;
  assign n19114 = P4_IR_REG_10_ & n19028;
  assign n19115 = ~P4_STATE_REG & P2_P3_DATAO_REG_10_;
  assign n19116 = ~n19114 & ~n19115;
  assign n19117 = P4_IR_REG_10_ & ~n19109;
  assign n19118 = ~P4_IR_REG_9_ & ~P4_IR_REG_10_;
  assign n19119 = n19102 & n19118;
  assign n19120 = ~n19117 & ~n19119;
  assign n19121 = n19032 & n19120;
  assign n2076 = ~n19116 | n19121;
  assign n19123 = P4_IR_REG_11_ & n19028;
  assign n19124 = ~P4_STATE_REG & P2_P3_DATAO_REG_11_;
  assign n19125 = ~n19123 & ~n19124;
  assign n19126 = P4_IR_REG_11_ & ~n19119;
  assign n19127 = ~P4_IR_REG_11_ & n19119;
  assign n19128 = ~n19126 & ~n19127;
  assign n19129 = n19032 & n19128;
  assign n2081 = ~n19125 | n19129;
  assign n19131 = P4_IR_REG_12_ & n19028;
  assign n19132 = ~P4_STATE_REG & P2_P3_DATAO_REG_12_;
  assign n19133 = ~n19131 & ~n19132;
  assign n19134 = P4_IR_REG_12_ & ~n19127;
  assign n19135 = ~P4_IR_REG_9_ & ~P4_IR_REG_12_;
  assign n19136 = ~P4_IR_REG_10_ & n19135;
  assign n19137 = ~P4_IR_REG_11_ & n19136;
  assign n19138 = n19102 & n19137;
  assign n19139 = ~n19134 & ~n19138;
  assign n19140 = n19032 & n19139;
  assign n2086 = ~n19133 | n19140;
  assign n19142 = P4_IR_REG_13_ & n19028;
  assign n19143 = ~P4_STATE_REG & P2_P3_DATAO_REG_13_;
  assign n19144 = ~n19142 & ~n19143;
  assign n19145 = ~P4_IR_REG_13_ & n19138;
  assign n19146 = P4_IR_REG_13_ & ~n19138;
  assign n19147 = ~n19145 & ~n19146;
  assign n19148 = n19032 & n19147;
  assign n2091 = ~n19144 | n19148;
  assign n19150 = P4_IR_REG_14_ & n19028;
  assign n19151 = ~P4_STATE_REG & P2_P3_DATAO_REG_14_;
  assign n19152 = ~n19150 & ~n19151;
  assign n19153 = P4_IR_REG_14_ & ~n19145;
  assign n19154 = ~P4_IR_REG_13_ & ~P4_IR_REG_14_;
  assign n19155 = n19138 & n19154;
  assign n19156 = ~n19153 & ~n19155;
  assign n19157 = n19032 & n19156;
  assign n2096 = ~n19152 | n19157;
  assign n19159 = P4_IR_REG_15_ & n19028;
  assign n19160 = ~P4_STATE_REG & P2_P3_DATAO_REG_15_;
  assign n19161 = ~n19159 & ~n19160;
  assign n19162 = P4_IR_REG_15_ & ~n19155;
  assign n19163 = ~P4_IR_REG_15_ & n19155;
  assign n19164 = ~n19162 & ~n19163;
  assign n19165 = n19032 & n19164;
  assign n2101 = ~n19161 | n19165;
  assign n19167 = P4_IR_REG_16_ & n19028;
  assign n19168 = ~P4_STATE_REG & P2_P3_DATAO_REG_16_;
  assign n19169 = ~n19167 & ~n19168;
  assign n19170 = P4_IR_REG_16_ & ~n19163;
  assign n19171 = ~P4_IR_REG_6_ & ~P4_IR_REG_7_;
  assign n19172 = ~P4_IR_REG_8_ & n19171;
  assign n19173 = ~P4_IR_REG_9_ & n19172;
  assign n19174 = ~P4_IR_REG_2_ & ~P4_IR_REG_3_;
  assign n19175 = ~P4_IR_REG_4_ & n19174;
  assign n19176 = ~P4_IR_REG_5_ & n19175;
  assign n19177 = ~P4_IR_REG_15_ & ~P4_IR_REG_16_;
  assign n19178 = ~P4_IR_REG_1_ & n19177;
  assign n19179 = ~P4_IR_REG_0_ & n19178;
  assign n19180 = ~P4_IR_REG_12_ & n19154;
  assign n19181 = ~P4_IR_REG_10_ & n19180;
  assign n19182 = ~P4_IR_REG_11_ & n19181;
  assign n19183 = n19173 & n19176;
  assign n19184 = n19179 & n19183;
  assign n19185 = n19182 & n19184;
  assign n19186 = ~n19170 & ~n19185;
  assign n19187 = n19032 & n19186;
  assign n2106 = ~n19169 | n19187;
  assign n19189 = P4_IR_REG_17_ & n19028;
  assign n19190 = ~P4_STATE_REG & P2_P3_DATAO_REG_17_;
  assign n19191 = ~n19189 & ~n19190;
  assign n19192 = ~P4_IR_REG_17_ & n19185;
  assign n19193 = P4_IR_REG_17_ & ~n19185;
  assign n19194 = ~n19192 & ~n19193;
  assign n19195 = n19032 & n19194;
  assign n2111 = ~n19191 | n19195;
  assign n19197 = P4_IR_REG_18_ & n19028;
  assign n19198 = ~P4_STATE_REG & P2_P3_DATAO_REG_18_;
  assign n19199 = ~n19197 & ~n19198;
  assign n19200 = P4_IR_REG_18_ & ~n19192;
  assign n19201 = ~P4_IR_REG_17_ & ~P4_IR_REG_18_;
  assign n19202 = n19185 & n19201;
  assign n19203 = ~n19200 & ~n19202;
  assign n19204 = n19032 & n19203;
  assign n2116 = ~n19199 | n19204;
  assign n19206 = P4_IR_REG_19_ & n19028;
  assign n19207 = ~P4_STATE_REG & P2_P3_DATAO_REG_19_;
  assign n19208 = ~n19206 & ~n19207;
  assign n19209 = ~P4_IR_REG_6_ & ~P4_IR_REG_8_;
  assign n19210 = ~P4_IR_REG_7_ & n19209;
  assign n19211 = ~P4_IR_REG_1_ & n19201;
  assign n19212 = ~P4_IR_REG_0_ & n19211;
  assign n19213 = ~P4_IR_REG_15_ & n19154;
  assign n19214 = ~P4_IR_REG_16_ & n19213;
  assign n19215 = n19137 & n19210;
  assign n19216 = n19176 & n19215;
  assign n19217 = n19212 & n19216;
  assign n19218 = n19214 & n19217;
  assign n19219 = ~P4_IR_REG_19_ & ~n19218;
  assign n19220 = P4_IR_REG_19_ & n19202;
  assign n19221 = ~n19219 & ~n19220;
  assign n19222 = n19032 & ~n19221;
  assign n2121 = ~n19208 | n19222;
  assign n19224 = P4_IR_REG_20_ & n19028;
  assign n19225 = ~P4_STATE_REG & P2_P3_DATAO_REG_20_;
  assign n19226 = ~n19224 & ~n19225;
  assign n19227 = ~P4_IR_REG_8_ & ~P4_IR_REG_9_;
  assign n19228 = ~P4_IR_REG_7_ & n19227;
  assign n19229 = ~P4_IR_REG_5_ & n19228;
  assign n19230 = ~P4_IR_REG_6_ & n19229;
  assign n19231 = ~P4_IR_REG_2_ & n19064;
  assign n19232 = ~P4_IR_REG_1_ & n19231;
  assign n19233 = ~P4_IR_REG_0_ & n19232;
  assign n19234 = ~P4_IR_REG_18_ & ~P4_IR_REG_19_;
  assign n19235 = ~P4_IR_REG_17_ & n19234;
  assign n19236 = ~P4_IR_REG_15_ & n19235;
  assign n19237 = ~P4_IR_REG_16_ & n19236;
  assign n19238 = n19230 & n19233;
  assign n19239 = n19237 & n19238;
  assign n19240 = n19182 & n19239;
  assign n19241 = ~P4_IR_REG_20_ & n19240;
  assign n19242 = P4_IR_REG_20_ & ~n19240;
  assign n19243 = ~n19241 & ~n19242;
  assign n19244 = n19032 & n19243;
  assign n2126 = ~n19226 | n19244;
  assign n19246 = P4_IR_REG_21_ & n19028;
  assign n19247 = ~P4_STATE_REG & P2_P3_DATAO_REG_21_;
  assign n19248 = ~n19246 & ~n19247;
  assign n19249 = ~P4_IR_REG_13_ & ~P4_IR_REG_15_;
  assign n19250 = ~P4_IR_REG_14_ & n19249;
  assign n19251 = ~P4_IR_REG_10_ & ~P4_IR_REG_12_;
  assign n19252 = ~P4_IR_REG_11_ & n19251;
  assign n19253 = ~P4_IR_REG_1_ & ~P4_IR_REG_19_;
  assign n19254 = ~P4_IR_REG_18_ & n19253;
  assign n19255 = ~P4_IR_REG_16_ & n19254;
  assign n19256 = ~P4_IR_REG_17_ & n19255;
  assign n19257 = ~P4_IR_REG_0_ & n19231;
  assign n19258 = ~P4_IR_REG_20_ & n19257;
  assign n19259 = n19250 & n19252;
  assign n19260 = n19256 & n19259;
  assign n19261 = n19230 & n19260;
  assign n19262 = n19258 & n19261;
  assign n19263 = P4_IR_REG_21_ & ~n19262;
  assign n19264 = ~P4_IR_REG_2_ & ~P4_IR_REG_4_;
  assign n19265 = ~P4_IR_REG_3_ & n19264;
  assign n19266 = ~P4_IR_REG_0_ & ~P4_IR_REG_21_;
  assign n19267 = ~P4_IR_REG_20_ & n19266;
  assign n19268 = n19265 & n19267;
  assign n19269 = n19230 & n19268;
  assign n19270 = n19256 & n19269;
  assign n19271 = n19259 & n19270;
  assign n19272 = ~n19263 & ~n19271;
  assign n19273 = n19032 & n19272;
  assign n2131 = ~n19248 | n19273;
  assign n19275 = P4_IR_REG_22_ & n19028;
  assign n19276 = ~P4_STATE_REG & P2_P3_DATAO_REG_22_;
  assign n19277 = ~n19275 & ~n19276;
  assign n19278 = ~P4_IR_REG_22_ & n19271;
  assign n19279 = P4_IR_REG_22_ & ~n19271;
  assign n19280 = ~n19278 & ~n19279;
  assign n19281 = n19032 & n19280;
  assign n2136 = ~n19277 | n19281;
  assign n19283 = P4_IR_REG_23_ & n19028;
  assign n19284 = ~P4_STATE_REG & P2_P3_DATAO_REG_23_;
  assign n19285 = ~n19283 & ~n19284;
  assign n19286 = ~P4_IR_REG_23_ & n19278;
  assign n19287 = P4_IR_REG_23_ & ~n19278;
  assign n19288 = ~n19286 & ~n19287;
  assign n19289 = n19032 & n19288;
  assign n2141 = ~n19285 | n19289;
  assign n19291 = P4_IR_REG_24_ & n19028;
  assign n19292 = ~P4_STATE_REG & P2_P3_DATAO_REG_24_;
  assign n19293 = ~n19291 & ~n19292;
  assign n19294 = P4_IR_REG_24_ & ~n19286;
  assign n19295 = ~P4_IR_REG_22_ & ~P4_IR_REG_24_;
  assign n19296 = ~P4_IR_REG_23_ & n19295;
  assign n19297 = n19271 & n19296;
  assign n19298 = ~n19294 & ~n19297;
  assign n19299 = n19032 & n19298;
  assign n2146 = ~n19293 | n19299;
  assign n19301 = P4_IR_REG_25_ & n19028;
  assign n19302 = ~P4_STATE_REG & P2_P3_DATAO_REG_25_;
  assign n19303 = ~n19301 & ~n19302;
  assign n19304 = ~P4_IR_REG_21_ & ~P4_IR_REG_22_;
  assign n19305 = ~P4_IR_REG_23_ & n19304;
  assign n19306 = ~P4_IR_REG_24_ & n19305;
  assign n19307 = ~P4_IR_REG_19_ & n19201;
  assign n19308 = ~P4_IR_REG_20_ & n19307;
  assign n19309 = n19306 & n19308;
  assign n19310 = n19185 & n19309;
  assign n19311 = P4_IR_REG_25_ & ~n19310;
  assign n19312 = ~P4_IR_REG_25_ & n19309;
  assign n19313 = n19185 & n19312;
  assign n19314 = ~n19311 & ~n19313;
  assign n19315 = n19032 & n19314;
  assign n2151 = ~n19303 | n19315;
  assign n19317 = P4_IR_REG_26_ & n19028;
  assign n19318 = ~P4_STATE_REG & P2_P3_DATAO_REG_26_;
  assign n19319 = ~n19317 & ~n19318;
  assign n19320 = P4_IR_REG_26_ & ~n19313;
  assign n19321 = ~P4_IR_REG_26_ & n19313;
  assign n19322 = ~n19320 & ~n19321;
  assign n19323 = n19032 & n19322;
  assign n2156 = ~n19319 | n19323;
  assign n19325 = P4_IR_REG_27_ & n19028;
  assign n19326 = ~P4_STATE_REG & P2_P3_DATAO_REG_27_;
  assign n19327 = ~n19325 & ~n19326;
  assign n19328 = ~P4_IR_REG_25_ & ~P4_IR_REG_26_;
  assign n19329 = n19297 & n19328;
  assign n19330 = ~P4_IR_REG_27_ & n19329;
  assign n19331 = P4_IR_REG_27_ & ~n19329;
  assign n19332 = ~n19330 & ~n19331;
  assign n19333 = n19032 & n19332;
  assign n2161 = ~n19327 | n19333;
  assign n19335 = P4_IR_REG_28_ & n19028;
  assign n19336 = ~P4_STATE_REG & P2_P3_DATAO_REG_28_;
  assign n19337 = ~n19335 & ~n19336;
  assign n19338 = ~P4_IR_REG_24_ & ~P4_IR_REG_25_;
  assign n19339 = ~P4_IR_REG_22_ & ~P4_IR_REG_23_;
  assign n19340 = ~P4_IR_REG_26_ & ~P4_IR_REG_27_;
  assign n19341 = n19338 & n19339;
  assign n19342 = n19340 & n19341;
  assign n19343 = n19271 & n19342;
  assign n19344 = ~P4_IR_REG_28_ & n19343;
  assign n19345 = P4_IR_REG_28_ & ~n19343;
  assign n19346 = ~n19344 & ~n19345;
  assign n19347 = n19032 & n19346;
  assign n2166 = ~n19337 | n19347;
  assign n19349 = P4_IR_REG_29_ & n19028;
  assign n19350 = ~P4_STATE_REG & P2_P3_DATAO_REG_29_;
  assign n19351 = ~n19349 & ~n19350;
  assign n19352 = ~P4_IR_REG_7_ & ~P4_IR_REG_9_;
  assign n19353 = ~P4_IR_REG_8_ & n19352;
  assign n19354 = ~P4_IR_REG_2_ & ~P4_IR_REG_27_;
  assign n19355 = ~P4_IR_REG_28_ & n19354;
  assign n19356 = ~P4_IR_REG_23_ & ~P4_IR_REG_24_;
  assign n19357 = ~P4_IR_REG_25_ & n19356;
  assign n19358 = ~P4_IR_REG_26_ & n19357;
  assign n19359 = n19100 & n19353;
  assign n19360 = n19355 & n19359;
  assign n19361 = n19358 & n19360;
  assign n19362 = ~P4_IR_REG_20_ & ~P4_IR_REG_22_;
  assign n19363 = ~P4_IR_REG_21_ & n19362;
  assign n19364 = ~P4_IR_REG_1_ & n19234;
  assign n19365 = ~P4_IR_REG_0_ & n19364;
  assign n19366 = ~P4_IR_REG_14_ & ~P4_IR_REG_15_;
  assign n19367 = ~P4_IR_REG_16_ & n19366;
  assign n19368 = ~P4_IR_REG_17_ & n19367;
  assign n19369 = ~P4_IR_REG_10_ & ~P4_IR_REG_11_;
  assign n19370 = ~P4_IR_REG_12_ & n19369;
  assign n19371 = ~P4_IR_REG_13_ & n19370;
  assign n19372 = n19363 & n19365;
  assign n19373 = n19368 & n19372;
  assign n19374 = n19371 & n19373;
  assign n19375 = n19361 & n19374;
  assign n19376 = ~P4_IR_REG_29_ & n19375;
  assign n19377 = P4_IR_REG_29_ & ~n19375;
  assign n19378 = ~n19376 & ~n19377;
  assign n19379 = n19032 & n19378;
  assign n2171 = ~n19351 | n19379;
  assign n19381 = P4_IR_REG_30_ & n19028;
  assign n19382 = ~P4_STATE_REG & P2_P3_DATAO_REG_30_;
  assign n19383 = ~n19381 & ~n19382;
  assign n19384 = ~P4_IR_REG_27_ & ~P4_IR_REG_28_;
  assign n19385 = ~P4_IR_REG_29_ & n19384;
  assign n19386 = ~P4_IR_REG_2_ & n19385;
  assign n19387 = n19359 & n19386;
  assign n19388 = n19358 & n19387;
  assign n19389 = n19374 & n19388;
  assign n19390 = ~P4_IR_REG_30_ & n19389;
  assign n19391 = P4_IR_REG_30_ & ~n19389;
  assign n19392 = ~n19390 & ~n19391;
  assign n19393 = n19032 & n19392;
  assign n2176 = ~n19383 | n19393;
  assign n19395 = P4_IR_REG_31_ & n19028;
  assign n19396 = ~P4_STATE_REG & P2_P3_DATAO_REG_31_;
  assign n19397 = ~n19395 & ~n19396;
  assign n19398 = ~P4_IR_REG_30_ & n19385;
  assign n19399 = n19321 & n19398;
  assign n19400 = ~P4_IR_REG_31_ & n19399;
  assign n19401 = P4_IR_REG_31_ & ~n19399;
  assign n19402 = ~n19400 & ~n19401;
  assign n19403 = n19032 & n19402;
  assign n2181 = ~n19397 | n19403;
  assign n19405 = P4_IR_REG_31_ & n19288;
  assign n19406 = P4_IR_REG_23_ & ~P4_IR_REG_31_;
  assign n19407 = ~n19405 & ~n19406;
  assign n19408 = P4_IR_REG_31_ & n19298;
  assign n19409 = P4_IR_REG_24_ & ~P4_IR_REG_31_;
  assign n19410 = ~n19408 & ~n19409;
  assign n19411 = P4_IR_REG_31_ & n19314;
  assign n19412 = P4_IR_REG_25_ & ~P4_IR_REG_31_;
  assign n19413 = ~n19411 & ~n19412;
  assign n19414 = P4_IR_REG_31_ & n19322;
  assign n19415 = P4_IR_REG_26_ & ~P4_IR_REG_31_;
  assign n19416 = ~n19414 & ~n19415;
  assign n19417 = ~n19410 & ~n19413;
  assign n19418 = ~n19416 & n19417;
  assign n19419 = n19407 & ~n19418;
  assign n19420 = P4_STATE_REG & n19419;
  assign n19421 = n19413 & ~n19416;
  assign n19422 = n19410 & n19421;
  assign n19423 = P4_B_REG & n19422;
  assign n19424 = ~P4_B_REG & ~n19410;
  assign n19425 = ~n19423 & ~n19424;
  assign n19426 = ~n19416 & n19425;
  assign n19427 = n19420 & ~n19426;
  assign n19428 = n19410 & ~n19421;
  assign n19429 = n19427 & ~n19428;
  assign n19430 = P4_D_REG_0_ & ~n19427;
  assign n2186 = n19429 | n19430;
  assign n19432 = n19413 & ~n19421;
  assign n19433 = n19427 & ~n19432;
  assign n19434 = P4_D_REG_1_ & ~n19427;
  assign n2191 = n19433 | n19434;
  assign n2196 = P4_D_REG_2_ & ~n19427;
  assign n2201 = P4_D_REG_3_ & ~n19427;
  assign n2206 = P4_D_REG_4_ & ~n19427;
  assign n2211 = P4_D_REG_5_ & ~n19427;
  assign n2216 = P4_D_REG_6_ & ~n19427;
  assign n2221 = P4_D_REG_7_ & ~n19427;
  assign n2226 = P4_D_REG_8_ & ~n19427;
  assign n2231 = P4_D_REG_9_ & ~n19427;
  assign n2236 = P4_D_REG_10_ & ~n19427;
  assign n2241 = P4_D_REG_11_ & ~n19427;
  assign n2246 = P4_D_REG_12_ & ~n19427;
  assign n2251 = P4_D_REG_13_ & ~n19427;
  assign n2256 = P4_D_REG_14_ & ~n19427;
  assign n2261 = P4_D_REG_15_ & ~n19427;
  assign n2266 = P4_D_REG_16_ & ~n19427;
  assign n2271 = P4_D_REG_17_ & ~n19427;
  assign n2276 = P4_D_REG_18_ & ~n19427;
  assign n2281 = P4_D_REG_19_ & ~n19427;
  assign n2286 = P4_D_REG_20_ & ~n19427;
  assign n2291 = P4_D_REG_21_ & ~n19427;
  assign n2296 = P4_D_REG_22_ & ~n19427;
  assign n2301 = P4_D_REG_23_ & ~n19427;
  assign n2306 = P4_D_REG_24_ & ~n19427;
  assign n2311 = P4_D_REG_25_ & ~n19427;
  assign n2316 = P4_D_REG_26_ & ~n19427;
  assign n2321 = P4_D_REG_27_ & ~n19427;
  assign n2326 = P4_D_REG_28_ & ~n19427;
  assign n2331 = P4_D_REG_29_ & ~n19427;
  assign n2336 = P4_D_REG_30_ & ~n19427;
  assign n2341 = P4_D_REG_31_ & ~n19427;
  assign n19466 = P4_D_REG_0_ & n19426;
  assign n19467 = n19410 & n19416;
  assign n19468 = ~n19426 & ~n19467;
  assign n19469 = ~n19466 & ~n19468;
  assign n19470 = n19420 & n19469;
  assign n19471 = ~n19426 & ~n19432;
  assign n19472 = P4_D_REG_1_ & n19426;
  assign n19473 = ~n19471 & ~n19472;
  assign n19474 = P4_IR_REG_31_ & n19243;
  assign n19475 = P4_IR_REG_20_ & ~P4_IR_REG_31_;
  assign n19476 = ~n19474 & ~n19475;
  assign n19477 = P4_IR_REG_31_ & ~n19221;
  assign n19478 = P4_IR_REG_19_ & ~P4_IR_REG_31_;
  assign n19479 = ~n19477 & ~n19478;
  assign n19480 = n19476 & n19479;
  assign n19481 = P4_IR_REG_31_ & n19272;
  assign n19482 = P4_IR_REG_21_ & ~P4_IR_REG_31_;
  assign n19483 = ~n19481 & ~n19482;
  assign n19484 = ~n19476 & n19483;
  assign n19485 = P4_IR_REG_31_ & n19280;
  assign n19486 = P4_IR_REG_22_ & ~P4_IR_REG_31_;
  assign n19487 = ~n19485 & ~n19486;
  assign n19488 = ~n19483 & n19487;
  assign n19489 = n19483 & ~n19487;
  assign n19490 = ~n19480 & ~n19484;
  assign n19491 = ~n19488 & n19490;
  assign n19492 = ~n19489 & n19491;
  assign n19493 = n19473 & ~n19492;
  assign n19494 = P4_D_REG_8_ & n19426;
  assign n19495 = P4_D_REG_7_ & n19426;
  assign n19496 = P4_D_REG_9_ & n19426;
  assign n19497 = ~n19494 & ~n19495;
  assign n19498 = ~n19496 & n19497;
  assign n19499 = P4_D_REG_6_ & n19426;
  assign n19500 = P4_D_REG_5_ & n19426;
  assign n19501 = P4_D_REG_4_ & n19426;
  assign n19502 = P4_D_REG_3_ & n19426;
  assign n19503 = ~n19499 & ~n19500;
  assign n19504 = ~n19501 & n19503;
  assign n19505 = ~n19502 & n19504;
  assign n19506 = P4_D_REG_31_ & n19426;
  assign n19507 = P4_D_REG_30_ & n19426;
  assign n19508 = P4_D_REG_2_ & n19426;
  assign n19509 = P4_D_REG_29_ & n19426;
  assign n19510 = ~n19506 & ~n19507;
  assign n19511 = ~n19508 & n19510;
  assign n19512 = ~n19509 & n19511;
  assign n19513 = P4_D_REG_28_ & n19426;
  assign n19514 = P4_D_REG_27_ & n19426;
  assign n19515 = P4_D_REG_26_ & n19426;
  assign n19516 = P4_D_REG_25_ & n19426;
  assign n19517 = ~n19513 & ~n19514;
  assign n19518 = ~n19515 & n19517;
  assign n19519 = ~n19516 & n19518;
  assign n19520 = n19498 & n19505;
  assign n19521 = n19512 & n19520;
  assign n19522 = n19519 & n19521;
  assign n19523 = P4_D_REG_23_ & n19426;
  assign n19524 = P4_D_REG_22_ & n19426;
  assign n19525 = P4_D_REG_24_ & n19426;
  assign n19526 = ~n19523 & ~n19524;
  assign n19527 = ~n19525 & n19526;
  assign n19528 = P4_D_REG_21_ & n19426;
  assign n19529 = P4_D_REG_20_ & n19426;
  assign n19530 = P4_D_REG_19_ & n19426;
  assign n19531 = P4_D_REG_18_ & n19426;
  assign n19532 = ~n19528 & ~n19529;
  assign n19533 = ~n19530 & n19532;
  assign n19534 = ~n19531 & n19533;
  assign n19535 = P4_D_REG_17_ & n19426;
  assign n19536 = P4_D_REG_16_ & n19426;
  assign n19537 = P4_D_REG_15_ & n19426;
  assign n19538 = P4_D_REG_14_ & n19426;
  assign n19539 = ~n19535 & ~n19536;
  assign n19540 = ~n19537 & n19539;
  assign n19541 = ~n19538 & n19540;
  assign n19542 = P4_D_REG_13_ & n19426;
  assign n19543 = P4_D_REG_12_ & n19426;
  assign n19544 = P4_D_REG_11_ & n19426;
  assign n19545 = P4_D_REG_10_ & n19426;
  assign n19546 = ~n19542 & ~n19543;
  assign n19547 = ~n19544 & n19546;
  assign n19548 = ~n19545 & n19547;
  assign n19549 = n19527 & n19534;
  assign n19550 = n19541 & n19549;
  assign n19551 = n19548 & n19550;
  assign n19552 = n19522 & n19551;
  assign n19553 = n19493 & n19552;
  assign n19554 = n19470 & n19553;
  assign n19555 = P4_IR_REG_31_ & n19332;
  assign n19556 = P4_IR_REG_27_ & ~P4_IR_REG_31_;
  assign n19557 = ~n19555 & ~n19556;
  assign n19558 = P4_IR_REG_31_ & n19346;
  assign n19559 = P4_IR_REG_28_ & ~P4_IR_REG_31_;
  assign n19560 = ~n19558 & ~n19559;
  assign n19561 = n19557 & n19560;
  assign n19562 = P4_IR_REG_0_ & P4_IR_REG_31_;
  assign n19563 = P4_IR_REG_0_ & ~P4_IR_REG_31_;
  assign n19564 = ~n19562 & ~n19563;
  assign n19565 = n19561 & ~n19564;
  assign n19566 = P2_P3_DATAO_REG_0_ & ~n19561;
  assign n19567 = ~n19565 & ~n19566;
  assign n19568 = n19484 & n19487;
  assign n19569 = ~n19567 & n19568;
  assign n19570 = n19476 & n19487;
  assign n19571 = n19483 & n19570;
  assign n19572 = ~n19567 & n19571;
  assign n19573 = ~n19483 & ~n19487;
  assign n19574 = n19560 & n19573;
  assign n19575 = P4_IR_REG_31_ & n19392;
  assign n19576 = P4_IR_REG_30_ & ~P4_IR_REG_31_;
  assign n19577 = ~n19575 & ~n19576;
  assign n19578 = P4_IR_REG_31_ & n19378;
  assign n19579 = P4_IR_REG_29_ & ~P4_IR_REG_31_;
  assign n19580 = ~n19578 & ~n19579;
  assign n19581 = ~n19577 & ~n19580;
  assign n19582 = P4_REG3_REG_1_ & n19581;
  assign n19583 = n19577 & n19580;
  assign n19584 = P4_REG0_REG_1_ & n19583;
  assign n19585 = n19577 & ~n19580;
  assign n19586 = P4_REG1_REG_1_ & n19585;
  assign n19587 = ~n19577 & n19580;
  assign n19588 = P4_REG2_REG_1_ & n19587;
  assign n19589 = ~n19582 & ~n19584;
  assign n19590 = ~n19586 & n19589;
  assign n19591 = ~n19588 & n19590;
  assign n19592 = n19574 & ~n19591;
  assign n19593 = P4_REG3_REG_0_ & n19581;
  assign n19594 = P4_REG2_REG_0_ & n19587;
  assign n19595 = P4_REG1_REG_0_ & n19585;
  assign n19596 = P4_REG0_REG_0_ & n19583;
  assign n19597 = ~n19593 & ~n19594;
  assign n19598 = ~n19595 & n19597;
  assign n19599 = ~n19596 & n19598;
  assign n19600 = ~n19567 & n19599;
  assign n19601 = n19567 & ~n19599;
  assign n19602 = ~n19600 & ~n19601;
  assign n19603 = ~n19479 & n19487;
  assign n19604 = n19476 & n19603;
  assign n19605 = ~n19602 & n19604;
  assign n19606 = ~n19569 & ~n19572;
  assign n19607 = ~n19592 & n19606;
  assign n19608 = ~n19605 & n19607;
  assign n19609 = n19476 & ~n19487;
  assign n19610 = n19479 & n19609;
  assign n19611 = n19483 & n19610;
  assign n19612 = ~n19602 & n19611;
  assign n19613 = ~n19476 & ~n19483;
  assign n19614 = n19479 & n19613;
  assign n19615 = ~n19602 & n19614;
  assign n19616 = n19480 & ~n19483;
  assign n19617 = n19487 & n19616;
  assign n19618 = ~n19602 & n19617;
  assign n19619 = ~n19479 & n19613;
  assign n19620 = ~n19602 & n19619;
  assign n19621 = ~n19476 & ~n19487;
  assign n19622 = n19479 & n19621;
  assign n19623 = ~n19602 & n19622;
  assign n19624 = ~n19620 & ~n19623;
  assign n19625 = ~n19479 & n19621;
  assign n19626 = ~n19602 & n19625;
  assign n19627 = ~n19479 & n19609;
  assign n19628 = ~n19602 & n19627;
  assign n19629 = ~n19626 & ~n19628;
  assign n19630 = ~n19612 & ~n19615;
  assign n19631 = ~n19618 & n19630;
  assign n19632 = n19624 & n19631;
  assign n19633 = n19629 & n19632;
  assign n19634 = n19608 & n19633;
  assign n19635 = n19554 & ~n19634;
  assign n19636 = P4_REG0_REG_0_ & ~n19554;
  assign n2346 = n19635 | n19636;
  assign n19638 = P4_IR_REG_31_ & ~n19040;
  assign n19639 = P4_IR_REG_1_ & ~P4_IR_REG_31_;
  assign n19640 = ~n19638 & ~n19639;
  assign n19641 = n19561 & ~n19640;
  assign n19642 = P2_P3_DATAO_REG_1_ & ~n19561;
  assign n19643 = ~n19641 & ~n19642;
  assign n19644 = n19568 & ~n19643;
  assign n19645 = ~n19591 & ~n19643;
  assign n19646 = n19591 & n19643;
  assign n19647 = ~n19645 & ~n19646;
  assign n19648 = ~n19567 & ~n19599;
  assign n19649 = n19647 & ~n19648;
  assign n19650 = ~n19647 & n19648;
  assign n19651 = ~n19649 & ~n19650;
  assign n19652 = n19604 & ~n19651;
  assign n19653 = P4_REG3_REG_2_ & n19581;
  assign n19654 = P4_REG0_REG_2_ & n19583;
  assign n19655 = P4_REG1_REG_2_ & n19585;
  assign n19656 = P4_REG2_REG_2_ & n19587;
  assign n19657 = ~n19653 & ~n19654;
  assign n19658 = ~n19655 & n19657;
  assign n19659 = ~n19656 & n19658;
  assign n19660 = n19574 & ~n19659;
  assign n19661 = ~n19567 & n19643;
  assign n19662 = n19567 & ~n19643;
  assign n19663 = ~n19661 & ~n19662;
  assign n19664 = n19571 & ~n19663;
  assign n19665 = ~n19644 & ~n19652;
  assign n19666 = ~n19660 & n19665;
  assign n19667 = ~n19664 & n19666;
  assign n19668 = ~n19591 & n19643;
  assign n19669 = n19591 & ~n19643;
  assign n19670 = ~n19668 & ~n19669;
  assign n19671 = ~n19600 & ~n19670;
  assign n19672 = n19600 & n19670;
  assign n19673 = ~n19671 & ~n19672;
  assign n19674 = n19627 & ~n19673;
  assign n19675 = ~n19560 & n19573;
  assign n19676 = ~n19599 & n19675;
  assign n19677 = n19622 & ~n19651;
  assign n19678 = n19625 & ~n19673;
  assign n19679 = ~n19677 & ~n19678;
  assign n19680 = n19617 & ~n19651;
  assign n19681 = n19611 & ~n19651;
  assign n19682 = n19614 & ~n19673;
  assign n19683 = n19619 & ~n19673;
  assign n19684 = ~n19682 & ~n19683;
  assign n19685 = ~n19680 & ~n19681;
  assign n19686 = n19684 & n19685;
  assign n19687 = ~n19674 & ~n19676;
  assign n19688 = n19679 & n19687;
  assign n19689 = n19686 & n19688;
  assign n19690 = n19667 & n19689;
  assign n19691 = n19554 & ~n19690;
  assign n19692 = P4_REG0_REG_1_ & ~n19554;
  assign n2351 = n19691 | n19692;
  assign n19694 = P4_IR_REG_31_ & n19049;
  assign n19695 = P4_IR_REG_2_ & ~P4_IR_REG_31_;
  assign n19696 = ~n19694 & ~n19695;
  assign n19697 = n19561 & ~n19696;
  assign n19698 = P2_P3_DATAO_REG_2_ & ~n19561;
  assign n19699 = ~n19697 & ~n19698;
  assign n19700 = n19568 & ~n19699;
  assign n19701 = ~n19659 & ~n19699;
  assign n19702 = n19659 & n19699;
  assign n19703 = ~n19701 & ~n19702;
  assign n19704 = ~n19646 & n19648;
  assign n19705 = ~n19645 & ~n19704;
  assign n19706 = n19703 & ~n19705;
  assign n19707 = n19659 & ~n19699;
  assign n19708 = ~n19659 & n19699;
  assign n19709 = ~n19707 & ~n19708;
  assign n19710 = ~n19645 & n19709;
  assign n19711 = ~n19704 & n19710;
  assign n19712 = ~n19706 & ~n19711;
  assign n19713 = n19604 & n19712;
  assign n19714 = ~P4_REG3_REG_3_ & n19581;
  assign n19715 = P4_REG0_REG_3_ & n19583;
  assign n19716 = P4_REG1_REG_3_ & n19585;
  assign n19717 = P4_REG2_REG_3_ & n19587;
  assign n19718 = ~n19714 & ~n19715;
  assign n19719 = ~n19716 & n19718;
  assign n19720 = ~n19717 & n19719;
  assign n19721 = n19574 & ~n19720;
  assign n19722 = n19567 & n19643;
  assign n19723 = ~n19699 & ~n19722;
  assign n19724 = n19699 & n19722;
  assign n19725 = ~n19723 & ~n19724;
  assign n19726 = n19571 & n19725;
  assign n19727 = ~n19700 & ~n19713;
  assign n19728 = ~n19721 & n19727;
  assign n19729 = ~n19726 & n19728;
  assign n19730 = ~n19600 & ~n19669;
  assign n19731 = ~n19668 & ~n19730;
  assign n19732 = n19709 & n19731;
  assign n19733 = ~n19709 & ~n19731;
  assign n19734 = ~n19732 & ~n19733;
  assign n19735 = n19627 & ~n19734;
  assign n19736 = ~n19591 & n19675;
  assign n19737 = n19622 & n19712;
  assign n19738 = n19625 & ~n19734;
  assign n19739 = ~n19737 & ~n19738;
  assign n19740 = n19617 & n19712;
  assign n19741 = n19611 & n19712;
  assign n19742 = n19614 & ~n19734;
  assign n19743 = n19619 & ~n19734;
  assign n19744 = ~n19742 & ~n19743;
  assign n19745 = ~n19740 & ~n19741;
  assign n19746 = n19744 & n19745;
  assign n19747 = ~n19735 & ~n19736;
  assign n19748 = n19739 & n19747;
  assign n19749 = n19746 & n19748;
  assign n19750 = n19729 & n19749;
  assign n19751 = n19554 & ~n19750;
  assign n19752 = P4_REG0_REG_2_ & ~n19554;
  assign n2356 = n19751 | n19752;
  assign n19754 = ~P4_REG3_REG_4_ & P4_REG3_REG_3_;
  assign n19755 = P4_REG3_REG_4_ & ~P4_REG3_REG_3_;
  assign n19756 = ~n19754 & ~n19755;
  assign n19757 = n19581 & ~n19756;
  assign n19758 = P4_REG0_REG_4_ & n19583;
  assign n19759 = P4_REG1_REG_4_ & n19585;
  assign n19760 = P4_REG2_REG_4_ & n19587;
  assign n19761 = ~n19757 & ~n19758;
  assign n19762 = ~n19759 & n19761;
  assign n19763 = ~n19760 & n19762;
  assign n19764 = n19574 & ~n19763;
  assign n19765 = P4_IR_REG_31_ & n19057;
  assign n19766 = P4_IR_REG_3_ & ~P4_IR_REG_31_;
  assign n19767 = ~n19765 & ~n19766;
  assign n19768 = n19561 & ~n19767;
  assign n19769 = P2_P3_DATAO_REG_3_ & ~n19561;
  assign n19770 = ~n19768 & ~n19769;
  assign n19771 = ~n19724 & ~n19770;
  assign n19772 = n19724 & n19770;
  assign n19773 = ~n19771 & ~n19772;
  assign n19774 = n19571 & n19773;
  assign n19775 = n19568 & ~n19770;
  assign n19776 = n19645 & ~n19702;
  assign n19777 = ~n19701 & ~n19776;
  assign n19778 = ~n19702 & n19704;
  assign n19779 = n19777 & ~n19778;
  assign n19780 = n19720 & ~n19770;
  assign n19781 = ~n19720 & n19770;
  assign n19782 = ~n19780 & ~n19781;
  assign n19783 = n19779 & ~n19782;
  assign n19784 = ~n19720 & ~n19770;
  assign n19785 = n19720 & n19770;
  assign n19786 = ~n19784 & ~n19785;
  assign n19787 = ~n19779 & ~n19786;
  assign n19788 = ~n19783 & ~n19787;
  assign n19789 = n19604 & ~n19788;
  assign n19790 = ~n19764 & ~n19774;
  assign n19791 = ~n19775 & n19790;
  assign n19792 = ~n19789 & n19791;
  assign n19793 = ~n19707 & ~n19782;
  assign n19794 = ~n19708 & n19731;
  assign n19795 = n19793 & ~n19794;
  assign n19796 = ~n19708 & n19782;
  assign n19797 = ~n19707 & ~n19731;
  assign n19798 = n19796 & ~n19797;
  assign n19799 = ~n19795 & ~n19798;
  assign n19800 = n19627 & ~n19799;
  assign n19801 = ~n19659 & n19675;
  assign n19802 = n19622 & ~n19788;
  assign n19803 = n19625 & ~n19799;
  assign n19804 = ~n19802 & ~n19803;
  assign n19805 = n19617 & ~n19788;
  assign n19806 = n19611 & ~n19788;
  assign n19807 = n19614 & ~n19799;
  assign n19808 = n19619 & ~n19799;
  assign n19809 = ~n19807 & ~n19808;
  assign n19810 = ~n19805 & ~n19806;
  assign n19811 = n19809 & n19810;
  assign n19812 = ~n19800 & ~n19801;
  assign n19813 = n19804 & n19812;
  assign n19814 = n19811 & n19813;
  assign n19815 = n19792 & n19814;
  assign n19816 = n19554 & ~n19815;
  assign n19817 = P4_REG0_REG_3_ & ~n19554;
  assign n2361 = n19816 | n19817;
  assign n19819 = P4_IR_REG_31_ & n19066;
  assign n19820 = P4_IR_REG_4_ & ~P4_IR_REG_31_;
  assign n19821 = ~n19819 & ~n19820;
  assign n19822 = n19561 & ~n19821;
  assign n19823 = P2_P3_DATAO_REG_4_ & ~n19561;
  assign n19824 = ~n19822 & ~n19823;
  assign n19825 = n19568 & ~n19824;
  assign n19826 = n19763 & ~n19824;
  assign n19827 = ~n19763 & n19824;
  assign n19828 = ~n19826 & ~n19827;
  assign n19829 = ~n19702 & ~n19785;
  assign n19830 = n19704 & n19829;
  assign n19831 = ~n19784 & ~n19830;
  assign n19832 = ~n19777 & ~n19785;
  assign n19833 = n19831 & ~n19832;
  assign n19834 = ~n19828 & n19833;
  assign n19835 = n19763 & n19824;
  assign n19836 = ~n19763 & ~n19824;
  assign n19837 = ~n19835 & ~n19836;
  assign n19838 = ~n19833 & ~n19837;
  assign n19839 = ~n19834 & ~n19838;
  assign n19840 = n19604 & ~n19839;
  assign n19841 = P4_REG3_REG_4_ & P4_REG3_REG_3_;
  assign n19842 = ~P4_REG3_REG_5_ & n19841;
  assign n19843 = P4_REG3_REG_5_ & ~n19841;
  assign n19844 = ~n19842 & ~n19843;
  assign n19845 = n19581 & ~n19844;
  assign n19846 = P4_REG0_REG_5_ & n19583;
  assign n19847 = P4_REG1_REG_5_ & n19585;
  assign n19848 = P4_REG2_REG_5_ & n19587;
  assign n19849 = ~n19845 & ~n19846;
  assign n19850 = ~n19847 & n19849;
  assign n19851 = ~n19848 & n19850;
  assign n19852 = n19574 & ~n19851;
  assign n19853 = ~n19772 & ~n19824;
  assign n19854 = n19770 & n19824;
  assign n19855 = n19724 & n19854;
  assign n19856 = ~n19853 & ~n19855;
  assign n19857 = n19571 & n19856;
  assign n19858 = ~n19825 & ~n19840;
  assign n19859 = ~n19852 & n19858;
  assign n19860 = ~n19857 & n19859;
  assign n19861 = n19708 & ~n19720;
  assign n19862 = ~n19770 & ~n19861;
  assign n19863 = ~n19708 & n19720;
  assign n19864 = ~n19862 & ~n19863;
  assign n19865 = ~n19707 & ~n19780;
  assign n19866 = ~n19731 & n19865;
  assign n19867 = ~n19864 & ~n19866;
  assign n19868 = n19828 & n19867;
  assign n19869 = ~n19828 & ~n19867;
  assign n19870 = ~n19868 & ~n19869;
  assign n19871 = n19627 & ~n19870;
  assign n19872 = n19675 & ~n19720;
  assign n19873 = n19622 & ~n19839;
  assign n19874 = n19625 & ~n19870;
  assign n19875 = ~n19873 & ~n19874;
  assign n19876 = n19617 & ~n19839;
  assign n19877 = n19611 & ~n19839;
  assign n19878 = n19614 & ~n19870;
  assign n19879 = n19619 & ~n19870;
  assign n19880 = ~n19878 & ~n19879;
  assign n19881 = ~n19876 & ~n19877;
  assign n19882 = n19880 & n19881;
  assign n19883 = ~n19871 & ~n19872;
  assign n19884 = n19875 & n19883;
  assign n19885 = n19882 & n19884;
  assign n19886 = n19860 & n19885;
  assign n19887 = n19554 & ~n19886;
  assign n19888 = P4_REG0_REG_4_ & ~n19554;
  assign n2366 = n19887 | n19888;
  assign n19890 = P4_REG3_REG_5_ & P4_REG3_REG_3_;
  assign n19891 = P4_REG3_REG_4_ & n19890;
  assign n19892 = ~P4_REG3_REG_6_ & n19891;
  assign n19893 = P4_REG3_REG_6_ & ~n19891;
  assign n19894 = ~n19892 & ~n19893;
  assign n19895 = n19581 & ~n19894;
  assign n19896 = P4_REG0_REG_6_ & n19583;
  assign n19897 = P4_REG1_REG_6_ & n19585;
  assign n19898 = P4_REG2_REG_6_ & n19587;
  assign n19899 = ~n19895 & ~n19896;
  assign n19900 = ~n19897 & n19899;
  assign n19901 = ~n19898 & n19900;
  assign n19902 = n19574 & ~n19901;
  assign n19903 = P4_IR_REG_31_ & n19074;
  assign n19904 = P4_IR_REG_5_ & ~P4_IR_REG_31_;
  assign n19905 = ~n19903 & ~n19904;
  assign n19906 = n19561 & ~n19905;
  assign n19907 = P2_P3_DATAO_REG_5_ & ~n19561;
  assign n19908 = ~n19906 & ~n19907;
  assign n19909 = ~n19855 & ~n19908;
  assign n19910 = n19855 & n19908;
  assign n19911 = ~n19909 & ~n19910;
  assign n19912 = n19571 & n19911;
  assign n19913 = n19568 & ~n19908;
  assign n19914 = ~n19851 & ~n19908;
  assign n19915 = n19851 & n19908;
  assign n19916 = ~n19835 & ~n19915;
  assign n19917 = ~n19914 & n19916;
  assign n19918 = n19833 & ~n19836;
  assign n19919 = n19917 & ~n19918;
  assign n19920 = n19851 & ~n19908;
  assign n19921 = ~n19851 & n19908;
  assign n19922 = ~n19920 & ~n19921;
  assign n19923 = ~n19836 & n19922;
  assign n19924 = ~n19833 & ~n19835;
  assign n19925 = n19923 & ~n19924;
  assign n19926 = ~n19919 & ~n19925;
  assign n19927 = n19604 & n19926;
  assign n19928 = ~n19902 & ~n19912;
  assign n19929 = ~n19913 & n19928;
  assign n19930 = ~n19927 & n19929;
  assign n19931 = ~n19826 & ~n19867;
  assign n19932 = ~n19827 & ~n19931;
  assign n19933 = n19922 & n19932;
  assign n19934 = ~n19922 & ~n19932;
  assign n19935 = ~n19933 & ~n19934;
  assign n19936 = n19627 & ~n19935;
  assign n19937 = n19675 & ~n19763;
  assign n19938 = n19622 & n19926;
  assign n19939 = n19625 & ~n19935;
  assign n19940 = ~n19938 & ~n19939;
  assign n19941 = n19617 & n19926;
  assign n19942 = n19611 & n19926;
  assign n19943 = n19614 & ~n19935;
  assign n19944 = n19619 & ~n19935;
  assign n19945 = ~n19943 & ~n19944;
  assign n19946 = ~n19941 & ~n19942;
  assign n19947 = n19945 & n19946;
  assign n19948 = ~n19936 & ~n19937;
  assign n19949 = n19940 & n19948;
  assign n19950 = n19947 & n19949;
  assign n19951 = n19930 & n19950;
  assign n19952 = n19554 & ~n19951;
  assign n19953 = P4_REG0_REG_5_ & ~n19554;
  assign n2371 = n19952 | n19953;
  assign n19955 = P4_REG3_REG_6_ & n19891;
  assign n19956 = ~P4_REG3_REG_7_ & n19955;
  assign n19957 = P4_REG3_REG_7_ & ~n19955;
  assign n19958 = ~n19956 & ~n19957;
  assign n19959 = n19581 & ~n19958;
  assign n19960 = P4_REG0_REG_7_ & n19583;
  assign n19961 = P4_REG1_REG_7_ & n19585;
  assign n19962 = P4_REG2_REG_7_ & n19587;
  assign n19963 = ~n19959 & ~n19960;
  assign n19964 = ~n19961 & n19963;
  assign n19965 = ~n19962 & n19964;
  assign n19966 = n19574 & ~n19965;
  assign n19967 = P4_IR_REG_31_ & n19083;
  assign n19968 = P4_IR_REG_6_ & ~P4_IR_REG_31_;
  assign n19969 = ~n19967 & ~n19968;
  assign n19970 = n19561 & ~n19969;
  assign n19971 = P2_P3_DATAO_REG_6_ & ~n19561;
  assign n19972 = ~n19970 & ~n19971;
  assign n19973 = ~n19910 & ~n19972;
  assign n19974 = n19908 & n19972;
  assign n19975 = n19855 & n19974;
  assign n19976 = ~n19973 & ~n19975;
  assign n19977 = n19571 & n19976;
  assign n19978 = n19568 & ~n19972;
  assign n19979 = n19901 & ~n19972;
  assign n19980 = ~n19901 & n19972;
  assign n19981 = ~n19979 & ~n19980;
  assign n19982 = n19836 & ~n19908;
  assign n19983 = ~n19836 & n19908;
  assign n19984 = ~n19851 & ~n19983;
  assign n19985 = ~n19982 & ~n19984;
  assign n19986 = ~n19785 & n19916;
  assign n19987 = ~n19701 & ~n19784;
  assign n19988 = ~n19702 & ~n19705;
  assign n19989 = n19987 & ~n19988;
  assign n19990 = n19986 & ~n19989;
  assign n19991 = n19985 & ~n19990;
  assign n19992 = ~n19981 & n19991;
  assign n19993 = n19901 & n19972;
  assign n19994 = ~n19901 & ~n19972;
  assign n19995 = ~n19993 & ~n19994;
  assign n19996 = ~n19991 & ~n19995;
  assign n19997 = ~n19992 & ~n19996;
  assign n19998 = n19604 & ~n19997;
  assign n19999 = ~n19966 & ~n19977;
  assign n20000 = ~n19978 & n19999;
  assign n20001 = ~n19998 & n20000;
  assign n20002 = ~n19920 & ~n19981;
  assign n20003 = ~n19921 & n19932;
  assign n20004 = n20002 & ~n20003;
  assign n20005 = ~n19921 & ~n19980;
  assign n20006 = ~n19979 & n20005;
  assign n20007 = ~n19920 & ~n19932;
  assign n20008 = n20006 & ~n20007;
  assign n20009 = ~n20004 & ~n20008;
  assign n20010 = n19627 & ~n20009;
  assign n20011 = n19675 & ~n19851;
  assign n20012 = n19622 & ~n19997;
  assign n20013 = n19625 & ~n20009;
  assign n20014 = ~n20012 & ~n20013;
  assign n20015 = n19617 & ~n19997;
  assign n20016 = n19611 & ~n19997;
  assign n20017 = n19614 & ~n20009;
  assign n20018 = n19619 & ~n20009;
  assign n20019 = ~n20017 & ~n20018;
  assign n20020 = ~n20015 & ~n20016;
  assign n20021 = n20019 & n20020;
  assign n20022 = ~n20010 & ~n20011;
  assign n20023 = n20014 & n20022;
  assign n20024 = n20021 & n20023;
  assign n20025 = n20001 & n20024;
  assign n20026 = n19554 & ~n20025;
  assign n20027 = P4_REG0_REG_6_ & ~n19554;
  assign n2376 = n20026 | n20027;
  assign n20029 = P4_REG3_REG_6_ & P4_REG3_REG_7_;
  assign n20030 = n19891 & n20029;
  assign n20031 = ~P4_REG3_REG_8_ & n20030;
  assign n20032 = P4_REG3_REG_8_ & ~n20030;
  assign n20033 = ~n20031 & ~n20032;
  assign n20034 = n19581 & ~n20033;
  assign n20035 = P4_REG0_REG_8_ & n19583;
  assign n20036 = P4_REG1_REG_8_ & n19585;
  assign n20037 = P4_REG2_REG_8_ & n19587;
  assign n20038 = ~n20034 & ~n20035;
  assign n20039 = ~n20036 & n20038;
  assign n20040 = ~n20037 & n20039;
  assign n20041 = n19574 & ~n20040;
  assign n20042 = P4_IR_REG_31_ & n19091;
  assign n20043 = P4_IR_REG_7_ & ~P4_IR_REG_31_;
  assign n20044 = ~n20042 & ~n20043;
  assign n20045 = n19561 & ~n20044;
  assign n20046 = P2_P3_DATAO_REG_7_ & ~n19561;
  assign n20047 = ~n20045 & ~n20046;
  assign n20048 = ~n19975 & ~n20047;
  assign n20049 = n19975 & n20047;
  assign n20050 = ~n20048 & ~n20049;
  assign n20051 = n19571 & n20050;
  assign n20052 = n19568 & ~n20047;
  assign n20053 = ~n19965 & ~n20047;
  assign n20054 = n19965 & n20047;
  assign n20055 = ~n19993 & ~n20054;
  assign n20056 = ~n20053 & n20055;
  assign n20057 = n19991 & ~n19994;
  assign n20058 = n20056 & ~n20057;
  assign n20059 = n19965 & ~n20047;
  assign n20060 = ~n19965 & n20047;
  assign n20061 = ~n20059 & ~n20060;
  assign n20062 = ~n19994 & n20061;
  assign n20063 = ~n19991 & ~n19993;
  assign n20064 = n20062 & ~n20063;
  assign n20065 = ~n20058 & ~n20064;
  assign n20066 = n19604 & n20065;
  assign n20067 = ~n20041 & ~n20051;
  assign n20068 = ~n20052 & n20067;
  assign n20069 = ~n20066 & n20068;
  assign n20070 = ~n19920 & ~n19979;
  assign n20071 = n19827 & n20070;
  assign n20072 = n20005 & ~n20071;
  assign n20073 = ~n19979 & ~n20072;
  assign n20074 = ~n19826 & n20070;
  assign n20075 = ~n19867 & n20074;
  assign n20076 = ~n20073 & ~n20075;
  assign n20077 = n20061 & n20076;
  assign n20078 = ~n20061 & ~n20076;
  assign n20079 = ~n20077 & ~n20078;
  assign n20080 = n19627 & ~n20079;
  assign n20081 = n19675 & ~n19901;
  assign n20082 = n19622 & n20065;
  assign n20083 = n19625 & ~n20079;
  assign n20084 = ~n20082 & ~n20083;
  assign n20085 = n19617 & n20065;
  assign n20086 = n19611 & n20065;
  assign n20087 = n19614 & ~n20079;
  assign n20088 = n19619 & ~n20079;
  assign n20089 = ~n20087 & ~n20088;
  assign n20090 = ~n20085 & ~n20086;
  assign n20091 = n20089 & n20090;
  assign n20092 = ~n20080 & ~n20081;
  assign n20093 = n20084 & n20092;
  assign n20094 = n20091 & n20093;
  assign n20095 = n20069 & n20094;
  assign n20096 = n19554 & ~n20095;
  assign n20097 = P4_REG0_REG_7_ & ~n19554;
  assign n2381 = n20096 | n20097;
  assign n20099 = P4_REG3_REG_8_ & n20030;
  assign n20100 = ~P4_REG3_REG_9_ & n20099;
  assign n20101 = P4_REG3_REG_9_ & ~n20099;
  assign n20102 = ~n20100 & ~n20101;
  assign n20103 = n19581 & ~n20102;
  assign n20104 = P4_REG0_REG_9_ & n19583;
  assign n20105 = P4_REG1_REG_9_ & n19585;
  assign n20106 = P4_REG2_REG_9_ & n19587;
  assign n20107 = ~n20103 & ~n20104;
  assign n20108 = ~n20105 & n20107;
  assign n20109 = ~n20106 & n20108;
  assign n20110 = n19574 & ~n20109;
  assign n20111 = P4_IR_REG_31_ & n19103;
  assign n20112 = P4_IR_REG_8_ & ~P4_IR_REG_31_;
  assign n20113 = ~n20111 & ~n20112;
  assign n20114 = n19561 & ~n20113;
  assign n20115 = P2_P3_DATAO_REG_8_ & ~n19561;
  assign n20116 = ~n20114 & ~n20115;
  assign n20117 = n20049 & n20116;
  assign n20118 = ~n20049 & ~n20116;
  assign n20119 = ~n20117 & ~n20118;
  assign n20120 = n19571 & n20119;
  assign n20121 = n19568 & ~n20116;
  assign n20122 = n19994 & ~n20047;
  assign n20123 = ~n19994 & n20047;
  assign n20124 = ~n19965 & ~n20123;
  assign n20125 = ~n20122 & ~n20124;
  assign n20126 = ~n19991 & n20055;
  assign n20127 = n20125 & ~n20126;
  assign n20128 = n20040 & ~n20116;
  assign n20129 = ~n20040 & n20116;
  assign n20130 = ~n20128 & ~n20129;
  assign n20131 = n20127 & ~n20130;
  assign n20132 = n20040 & n20116;
  assign n20133 = ~n20040 & ~n20116;
  assign n20134 = ~n20132 & ~n20133;
  assign n20135 = ~n20127 & ~n20134;
  assign n20136 = ~n20131 & ~n20135;
  assign n20137 = n19604 & ~n20136;
  assign n20138 = ~n20110 & ~n20120;
  assign n20139 = ~n20121 & n20138;
  assign n20140 = ~n20137 & n20139;
  assign n20141 = ~n20059 & ~n20130;
  assign n20142 = ~n20060 & n20076;
  assign n20143 = n20141 & ~n20142;
  assign n20144 = ~n20060 & n20130;
  assign n20145 = ~n20059 & ~n20076;
  assign n20146 = n20144 & ~n20145;
  assign n20147 = ~n20143 & ~n20146;
  assign n20148 = n19627 & ~n20147;
  assign n20149 = n19675 & ~n19965;
  assign n20150 = n19622 & ~n20136;
  assign n20151 = n19625 & ~n20147;
  assign n20152 = ~n20150 & ~n20151;
  assign n20153 = n19617 & ~n20136;
  assign n20154 = n19611 & ~n20136;
  assign n20155 = n19614 & ~n20147;
  assign n20156 = n19619 & ~n20147;
  assign n20157 = ~n20155 & ~n20156;
  assign n20158 = ~n20153 & ~n20154;
  assign n20159 = n20157 & n20158;
  assign n20160 = ~n20148 & ~n20149;
  assign n20161 = n20152 & n20160;
  assign n20162 = n20159 & n20161;
  assign n20163 = n20140 & n20162;
  assign n20164 = n19554 & ~n20163;
  assign n20165 = P4_REG0_REG_8_ & ~n19554;
  assign n2386 = n20164 | n20165;
  assign n20167 = P4_REG3_REG_9_ & P4_REG3_REG_8_;
  assign n20168 = n20030 & n20167;
  assign n20169 = ~P4_REG3_REG_10_ & n20168;
  assign n20170 = P4_REG3_REG_10_ & ~n20168;
  assign n20171 = ~n20169 & ~n20170;
  assign n20172 = n19581 & ~n20171;
  assign n20173 = P4_REG0_REG_10_ & n19583;
  assign n20174 = P4_REG1_REG_10_ & n19585;
  assign n20175 = P4_REG2_REG_10_ & n19587;
  assign n20176 = ~n20172 & ~n20173;
  assign n20177 = ~n20174 & n20176;
  assign n20178 = ~n20175 & n20177;
  assign n20179 = n19574 & ~n20178;
  assign n20180 = n20047 & n20116;
  assign n20181 = n19975 & n20180;
  assign n20182 = P4_IR_REG_31_ & n19111;
  assign n20183 = P4_IR_REG_9_ & ~P4_IR_REG_31_;
  assign n20184 = ~n20182 & ~n20183;
  assign n20185 = n19561 & ~n20184;
  assign n20186 = P2_P3_DATAO_REG_9_ & ~n19561;
  assign n20187 = ~n20185 & ~n20186;
  assign n20188 = n20181 & n20187;
  assign n20189 = ~n20181 & ~n20187;
  assign n20190 = ~n20188 & ~n20189;
  assign n20191 = n19571 & n20190;
  assign n20192 = n19568 & ~n20187;
  assign n20193 = n20109 & ~n20187;
  assign n20194 = ~n20109 & n20187;
  assign n20195 = ~n20193 & ~n20194;
  assign n20196 = ~n20127 & ~n20132;
  assign n20197 = ~n20133 & ~n20196;
  assign n20198 = ~n20195 & n20197;
  assign n20199 = n20109 & n20187;
  assign n20200 = ~n20109 & ~n20187;
  assign n20201 = ~n20199 & ~n20200;
  assign n20202 = ~n20197 & ~n20201;
  assign n20203 = ~n20198 & ~n20202;
  assign n20204 = n19604 & ~n20203;
  assign n20205 = ~n20179 & ~n20191;
  assign n20206 = ~n20192 & n20205;
  assign n20207 = ~n20204 & n20206;
  assign n20208 = ~n20040 & n20060;
  assign n20209 = n20040 & ~n20060;
  assign n20210 = n20116 & ~n20209;
  assign n20211 = ~n20208 & ~n20210;
  assign n20212 = ~n20059 & ~n20128;
  assign n20213 = ~n20076 & n20212;
  assign n20214 = n20211 & ~n20213;
  assign n20215 = n20195 & n20214;
  assign n20216 = ~n20195 & ~n20214;
  assign n20217 = ~n20215 & ~n20216;
  assign n20218 = n19627 & ~n20217;
  assign n20219 = n19675 & ~n20040;
  assign n20220 = n19622 & ~n20203;
  assign n20221 = n19625 & ~n20217;
  assign n20222 = ~n20220 & ~n20221;
  assign n20223 = n19617 & ~n20203;
  assign n20224 = n19611 & ~n20203;
  assign n20225 = n19614 & ~n20217;
  assign n20226 = n19619 & ~n20217;
  assign n20227 = ~n20225 & ~n20226;
  assign n20228 = ~n20223 & ~n20224;
  assign n20229 = n20227 & n20228;
  assign n20230 = ~n20218 & ~n20219;
  assign n20231 = n20222 & n20230;
  assign n20232 = n20229 & n20231;
  assign n20233 = n20207 & n20232;
  assign n20234 = n19554 & ~n20233;
  assign n20235 = P4_REG0_REG_9_ & ~n19554;
  assign n2391 = n20234 | n20235;
  assign n20237 = P4_REG3_REG_10_ & n20168;
  assign n20238 = ~P4_REG3_REG_11_ & n20237;
  assign n20239 = P4_REG3_REG_11_ & ~n20237;
  assign n20240 = ~n20238 & ~n20239;
  assign n20241 = n19581 & ~n20240;
  assign n20242 = P4_REG0_REG_11_ & n19583;
  assign n20243 = P4_REG1_REG_11_ & n19585;
  assign n20244 = P4_REG2_REG_11_ & n19587;
  assign n20245 = ~n20241 & ~n20242;
  assign n20246 = ~n20243 & n20245;
  assign n20247 = ~n20244 & n20246;
  assign n20248 = n19574 & ~n20247;
  assign n20249 = P4_IR_REG_31_ & n19120;
  assign n20250 = P4_IR_REG_10_ & ~P4_IR_REG_31_;
  assign n20251 = ~n20249 & ~n20250;
  assign n20252 = n19561 & ~n20251;
  assign n20253 = P2_P3_DATAO_REG_10_ & ~n19561;
  assign n20254 = ~n20252 & ~n20253;
  assign n20255 = n20188 & n20254;
  assign n20256 = ~n20188 & ~n20254;
  assign n20257 = ~n20255 & ~n20256;
  assign n20258 = n19571 & n20257;
  assign n20259 = n19568 & ~n20254;
  assign n20260 = ~n20178 & ~n20254;
  assign n20261 = n20178 & n20254;
  assign n20262 = ~n20199 & ~n20261;
  assign n20263 = ~n20260 & n20262;
  assign n20264 = n20197 & ~n20200;
  assign n20265 = n20263 & ~n20264;
  assign n20266 = n20178 & ~n20254;
  assign n20267 = ~n20178 & n20254;
  assign n20268 = ~n20266 & ~n20267;
  assign n20269 = ~n20200 & n20268;
  assign n20270 = ~n20197 & ~n20199;
  assign n20271 = n20269 & ~n20270;
  assign n20272 = ~n20265 & ~n20271;
  assign n20273 = n19604 & n20272;
  assign n20274 = ~n20248 & ~n20258;
  assign n20275 = ~n20259 & n20274;
  assign n20276 = ~n20273 & n20275;
  assign n20277 = ~n20193 & ~n20214;
  assign n20278 = ~n20194 & ~n20277;
  assign n20279 = n20268 & n20278;
  assign n20280 = ~n20268 & ~n20278;
  assign n20281 = ~n20279 & ~n20280;
  assign n20282 = n19627 & ~n20281;
  assign n20283 = n19675 & ~n20109;
  assign n20284 = n19622 & n20272;
  assign n20285 = n19625 & ~n20281;
  assign n20286 = ~n20284 & ~n20285;
  assign n20287 = n19617 & n20272;
  assign n20288 = n19611 & n20272;
  assign n20289 = n19614 & ~n20281;
  assign n20290 = n19619 & ~n20281;
  assign n20291 = ~n20289 & ~n20290;
  assign n20292 = ~n20287 & ~n20288;
  assign n20293 = n20291 & n20292;
  assign n20294 = ~n20282 & ~n20283;
  assign n20295 = n20286 & n20294;
  assign n20296 = n20293 & n20295;
  assign n20297 = n20276 & n20296;
  assign n20298 = n19554 & ~n20297;
  assign n20299 = P4_REG0_REG_10_ & ~n19554;
  assign n2396 = n20298 | n20299;
  assign n20301 = P4_REG3_REG_11_ & n20237;
  assign n20302 = ~P4_REG3_REG_12_ & n20301;
  assign n20303 = P4_REG3_REG_12_ & ~n20301;
  assign n20304 = ~n20302 & ~n20303;
  assign n20305 = n19581 & ~n20304;
  assign n20306 = P4_REG0_REG_12_ & n19583;
  assign n20307 = P4_REG1_REG_12_ & n19585;
  assign n20308 = P4_REG2_REG_12_ & n19587;
  assign n20309 = ~n20305 & ~n20306;
  assign n20310 = ~n20307 & n20309;
  assign n20311 = ~n20308 & n20310;
  assign n20312 = n19574 & ~n20311;
  assign n20313 = n20187 & n20254;
  assign n20314 = n20181 & n20313;
  assign n20315 = P4_IR_REG_31_ & n19128;
  assign n20316 = P4_IR_REG_11_ & ~P4_IR_REG_31_;
  assign n20317 = ~n20315 & ~n20316;
  assign n20318 = n19561 & ~n20317;
  assign n20319 = P2_P3_DATAO_REG_11_ & ~n19561;
  assign n20320 = ~n20318 & ~n20319;
  assign n20321 = n20314 & n20320;
  assign n20322 = ~n20314 & ~n20320;
  assign n20323 = ~n20321 & ~n20322;
  assign n20324 = n19571 & n20323;
  assign n20325 = n19568 & ~n20320;
  assign n20326 = ~n20200 & ~n20260;
  assign n20327 = n20133 & n20262;
  assign n20328 = n20326 & ~n20327;
  assign n20329 = ~n20261 & ~n20328;
  assign n20330 = ~n20132 & n20262;
  assign n20331 = ~n20127 & n20330;
  assign n20332 = ~n20329 & ~n20331;
  assign n20333 = n20247 & ~n20320;
  assign n20334 = ~n20247 & n20320;
  assign n20335 = ~n20333 & ~n20334;
  assign n20336 = n20332 & ~n20335;
  assign n20337 = n20247 & n20320;
  assign n20338 = ~n20247 & ~n20320;
  assign n20339 = ~n20337 & ~n20338;
  assign n20340 = ~n20332 & ~n20339;
  assign n20341 = ~n20336 & ~n20340;
  assign n20342 = n19604 & ~n20341;
  assign n20343 = ~n20312 & ~n20324;
  assign n20344 = ~n20325 & n20343;
  assign n20345 = ~n20342 & n20344;
  assign n20346 = ~n20266 & ~n20335;
  assign n20347 = ~n20267 & n20278;
  assign n20348 = n20346 & ~n20347;
  assign n20349 = ~n20267 & ~n20334;
  assign n20350 = ~n20333 & n20349;
  assign n20351 = ~n20266 & ~n20278;
  assign n20352 = n20350 & ~n20351;
  assign n20353 = ~n20348 & ~n20352;
  assign n20354 = n19627 & ~n20353;
  assign n20355 = n19675 & ~n20178;
  assign n20356 = n19622 & ~n20341;
  assign n20357 = n19625 & ~n20353;
  assign n20358 = ~n20356 & ~n20357;
  assign n20359 = ~n20200 & ~n20327;
  assign n20360 = ~n20261 & ~n20359;
  assign n20361 = ~n20260 & ~n20360;
  assign n20362 = ~n20331 & n20361;
  assign n20363 = ~n20335 & n20362;
  assign n20364 = ~n20339 & ~n20362;
  assign n20365 = ~n20363 & ~n20364;
  assign n20366 = n19617 & ~n20365;
  assign n20367 = n19611 & ~n20365;
  assign n20368 = n19614 & ~n20353;
  assign n20369 = n19619 & ~n20353;
  assign n20370 = ~n20368 & ~n20369;
  assign n20371 = ~n20366 & ~n20367;
  assign n20372 = n20370 & n20371;
  assign n20373 = ~n20354 & ~n20355;
  assign n20374 = n20358 & n20373;
  assign n20375 = n20372 & n20374;
  assign n20376 = n20345 & n20375;
  assign n20377 = n19554 & ~n20376;
  assign n20378 = P4_REG0_REG_11_ & ~n19554;
  assign n2401 = n20377 | n20378;
  assign n20380 = P4_REG1_REG_13_ & n19585;
  assign n20381 = P4_REG2_REG_13_ & n19587;
  assign n20382 = P4_REG0_REG_13_ & n19583;
  assign n20383 = P4_REG3_REG_12_ & n20301;
  assign n20384 = ~P4_REG3_REG_13_ & n20383;
  assign n20385 = P4_REG3_REG_13_ & ~n20383;
  assign n20386 = ~n20384 & ~n20385;
  assign n20387 = n19581 & ~n20386;
  assign n20388 = ~n20380 & ~n20381;
  assign n20389 = ~n20382 & n20388;
  assign n20390 = ~n20387 & n20389;
  assign n20391 = n19574 & ~n20390;
  assign n20392 = P4_IR_REG_31_ & n19139;
  assign n20393 = P4_IR_REG_12_ & ~P4_IR_REG_31_;
  assign n20394 = ~n20392 & ~n20393;
  assign n20395 = n19561 & ~n20394;
  assign n20396 = P2_P3_DATAO_REG_12_ & ~n19561;
  assign n20397 = ~n20395 & ~n20396;
  assign n20398 = n20321 & n20397;
  assign n20399 = ~n20321 & ~n20397;
  assign n20400 = ~n20398 & ~n20399;
  assign n20401 = n19571 & n20400;
  assign n20402 = n19568 & ~n20397;
  assign n20403 = n20311 & ~n20397;
  assign n20404 = ~n20311 & n20397;
  assign n20405 = ~n20403 & ~n20404;
  assign n20406 = ~n20332 & ~n20337;
  assign n20407 = ~n20338 & ~n20406;
  assign n20408 = ~n20405 & n20407;
  assign n20409 = n20311 & n20397;
  assign n20410 = ~n20311 & ~n20397;
  assign n20411 = ~n20409 & ~n20410;
  assign n20412 = ~n20407 & ~n20411;
  assign n20413 = ~n20408 & ~n20412;
  assign n20414 = n19604 & ~n20413;
  assign n20415 = ~n20391 & ~n20401;
  assign n20416 = ~n20402 & n20415;
  assign n20417 = ~n20414 & n20416;
  assign n20418 = ~n20266 & ~n20333;
  assign n20419 = n20194 & n20418;
  assign n20420 = n20349 & ~n20419;
  assign n20421 = ~n20333 & ~n20420;
  assign n20422 = ~n20193 & n20418;
  assign n20423 = ~n20214 & n20422;
  assign n20424 = ~n20421 & ~n20423;
  assign n20425 = ~n20405 & ~n20424;
  assign n20426 = n20405 & n20424;
  assign n20427 = ~n20425 & ~n20426;
  assign n20428 = n19627 & ~n20427;
  assign n20429 = n19675 & ~n20247;
  assign n20430 = n19622 & ~n20413;
  assign n20431 = n19625 & ~n20427;
  assign n20432 = ~n20430 & ~n20431;
  assign n20433 = ~n20337 & ~n20362;
  assign n20434 = ~n20338 & ~n20433;
  assign n20435 = ~n20405 & n20434;
  assign n20436 = ~n20411 & ~n20434;
  assign n20437 = ~n20435 & ~n20436;
  assign n20438 = n19617 & ~n20437;
  assign n20439 = n19611 & ~n20437;
  assign n20440 = n19614 & ~n20427;
  assign n20441 = n19619 & ~n20427;
  assign n20442 = ~n20440 & ~n20441;
  assign n20443 = ~n20438 & ~n20439;
  assign n20444 = n20442 & n20443;
  assign n20445 = ~n20428 & ~n20429;
  assign n20446 = n20432 & n20445;
  assign n20447 = n20444 & n20446;
  assign n20448 = n20417 & n20447;
  assign n20449 = n19554 & ~n20448;
  assign n20450 = P4_REG0_REG_12_ & ~n19554;
  assign n2406 = n20449 | n20450;
  assign n20452 = P4_REG1_REG_14_ & n19585;
  assign n20453 = P4_REG2_REG_14_ & n19587;
  assign n20454 = P4_REG0_REG_14_ & n19583;
  assign n20455 = P4_REG3_REG_13_ & n20383;
  assign n20456 = ~P4_REG3_REG_14_ & n20455;
  assign n20457 = P4_REG3_REG_14_ & ~n20455;
  assign n20458 = ~n20456 & ~n20457;
  assign n20459 = n19581 & ~n20458;
  assign n20460 = ~n20452 & ~n20453;
  assign n20461 = ~n20454 & n20460;
  assign n20462 = ~n20459 & n20461;
  assign n20463 = n19574 & ~n20462;
  assign n20464 = n20320 & n20397;
  assign n20465 = n20314 & n20464;
  assign n20466 = P4_IR_REG_31_ & n19147;
  assign n20467 = P4_IR_REG_13_ & ~P4_IR_REG_31_;
  assign n20468 = ~n20466 & ~n20467;
  assign n20469 = n19561 & ~n20468;
  assign n20470 = P2_P3_DATAO_REG_13_ & ~n19561;
  assign n20471 = ~n20469 & ~n20470;
  assign n20472 = n20465 & n20471;
  assign n20473 = ~n20465 & ~n20471;
  assign n20474 = ~n20472 & ~n20473;
  assign n20475 = n19571 & n20474;
  assign n20476 = n19568 & ~n20471;
  assign n20477 = ~n20390 & ~n20471;
  assign n20478 = n20390 & n20471;
  assign n20479 = ~n20409 & ~n20478;
  assign n20480 = ~n20477 & n20479;
  assign n20481 = n20407 & ~n20410;
  assign n20482 = n20480 & ~n20481;
  assign n20483 = n20390 & ~n20471;
  assign n20484 = ~n20390 & n20471;
  assign n20485 = ~n20483 & ~n20484;
  assign n20486 = ~n20410 & n20485;
  assign n20487 = ~n20407 & ~n20409;
  assign n20488 = n20486 & ~n20487;
  assign n20489 = ~n20482 & ~n20488;
  assign n20490 = n19604 & n20489;
  assign n20491 = ~n20463 & ~n20475;
  assign n20492 = ~n20476 & n20491;
  assign n20493 = ~n20490 & n20492;
  assign n20494 = ~n20403 & ~n20424;
  assign n20495 = ~n20404 & ~n20494;
  assign n20496 = ~n20485 & ~n20495;
  assign n20497 = n20485 & n20495;
  assign n20498 = ~n20496 & ~n20497;
  assign n20499 = n19627 & ~n20498;
  assign n20500 = n19675 & ~n20311;
  assign n20501 = n19622 & n20489;
  assign n20502 = n19625 & ~n20498;
  assign n20503 = ~n20501 & ~n20502;
  assign n20504 = ~n20410 & n20434;
  assign n20505 = n20480 & ~n20504;
  assign n20506 = ~n20409 & ~n20434;
  assign n20507 = n20486 & ~n20506;
  assign n20508 = ~n20505 & ~n20507;
  assign n20509 = n19617 & n20508;
  assign n20510 = n19611 & n20508;
  assign n20511 = n19614 & ~n20498;
  assign n20512 = n19619 & ~n20498;
  assign n20513 = ~n20511 & ~n20512;
  assign n20514 = ~n20509 & ~n20510;
  assign n20515 = n20513 & n20514;
  assign n20516 = ~n20499 & ~n20500;
  assign n20517 = n20503 & n20516;
  assign n20518 = n20515 & n20517;
  assign n20519 = n20493 & n20518;
  assign n20520 = n19554 & ~n20519;
  assign n20521 = P4_REG0_REG_13_ & ~n19554;
  assign n2411 = n20520 | n20521;
  assign n20523 = P4_REG1_REG_15_ & n19585;
  assign n20524 = P4_REG2_REG_15_ & n19587;
  assign n20525 = P4_REG0_REG_15_ & n19583;
  assign n20526 = P4_REG3_REG_14_ & n20455;
  assign n20527 = ~P4_REG3_REG_15_ & n20526;
  assign n20528 = P4_REG3_REG_15_ & ~n20526;
  assign n20529 = ~n20527 & ~n20528;
  assign n20530 = n19581 & ~n20529;
  assign n20531 = ~n20523 & ~n20524;
  assign n20532 = ~n20525 & n20531;
  assign n20533 = ~n20530 & n20532;
  assign n20534 = n19574 & ~n20533;
  assign n20535 = P4_IR_REG_31_ & n19156;
  assign n20536 = P4_IR_REG_14_ & ~P4_IR_REG_31_;
  assign n20537 = ~n20535 & ~n20536;
  assign n20538 = n19561 & ~n20537;
  assign n20539 = P2_P3_DATAO_REG_14_ & ~n19561;
  assign n20540 = ~n20538 & ~n20539;
  assign n20541 = n20472 & n20540;
  assign n20542 = ~n20472 & ~n20540;
  assign n20543 = ~n20541 & ~n20542;
  assign n20544 = n19571 & n20543;
  assign n20545 = n19568 & ~n20540;
  assign n20546 = ~n20410 & ~n20477;
  assign n20547 = n20338 & n20479;
  assign n20548 = n20546 & ~n20547;
  assign n20549 = ~n20478 & ~n20548;
  assign n20550 = ~n20337 & n20479;
  assign n20551 = ~n20332 & n20550;
  assign n20552 = ~n20549 & ~n20551;
  assign n20553 = n20462 & ~n20540;
  assign n20554 = ~n20462 & n20540;
  assign n20555 = ~n20553 & ~n20554;
  assign n20556 = n20552 & ~n20555;
  assign n20557 = ~n20552 & n20555;
  assign n20558 = ~n20556 & ~n20557;
  assign n20559 = n19604 & ~n20558;
  assign n20560 = ~n20534 & ~n20544;
  assign n20561 = ~n20545 & n20560;
  assign n20562 = ~n20559 & n20561;
  assign n20563 = ~n20483 & ~n20495;
  assign n20564 = ~n20484 & ~n20563;
  assign n20565 = n20555 & n20564;
  assign n20566 = ~n20555 & ~n20564;
  assign n20567 = ~n20565 & ~n20566;
  assign n20568 = n19627 & ~n20567;
  assign n20569 = n19675 & ~n20390;
  assign n20570 = n19622 & ~n20558;
  assign n20571 = n19625 & ~n20567;
  assign n20572 = ~n20570 & ~n20571;
  assign n20573 = ~n20362 & n20550;
  assign n20574 = ~n20549 & ~n20573;
  assign n20575 = ~n20555 & n20574;
  assign n20576 = n20555 & ~n20574;
  assign n20577 = ~n20575 & ~n20576;
  assign n20578 = n19617 & ~n20577;
  assign n20579 = n19611 & ~n20577;
  assign n20580 = n19614 & ~n20567;
  assign n20581 = n19619 & ~n20567;
  assign n20582 = ~n20580 & ~n20581;
  assign n20583 = ~n20578 & ~n20579;
  assign n20584 = n20582 & n20583;
  assign n20585 = ~n20568 & ~n20569;
  assign n20586 = n20572 & n20585;
  assign n20587 = n20584 & n20586;
  assign n20588 = n20562 & n20587;
  assign n20589 = n19554 & ~n20588;
  assign n20590 = P4_REG0_REG_14_ & ~n19554;
  assign n2416 = n20589 | n20590;
  assign n20592 = P4_REG1_REG_16_ & n19585;
  assign n20593 = P4_REG2_REG_16_ & n19587;
  assign n20594 = P4_REG0_REG_16_ & n19583;
  assign n20595 = P4_REG3_REG_15_ & n20526;
  assign n20596 = ~P4_REG3_REG_16_ & n20595;
  assign n20597 = P4_REG3_REG_16_ & ~n20595;
  assign n20598 = ~n20596 & ~n20597;
  assign n20599 = n19581 & ~n20598;
  assign n20600 = ~n20592 & ~n20593;
  assign n20601 = ~n20594 & n20600;
  assign n20602 = ~n20599 & n20601;
  assign n20603 = n19574 & ~n20602;
  assign n20604 = n20471 & n20540;
  assign n20605 = n20465 & n20604;
  assign n20606 = P4_IR_REG_31_ & n19164;
  assign n20607 = P4_IR_REG_15_ & ~P4_IR_REG_31_;
  assign n20608 = ~n20606 & ~n20607;
  assign n20609 = n19561 & ~n20608;
  assign n20610 = P2_P3_DATAO_REG_15_ & ~n19561;
  assign n20611 = ~n20609 & ~n20610;
  assign n20612 = n20605 & n20611;
  assign n20613 = ~n20605 & ~n20611;
  assign n20614 = ~n20612 & ~n20613;
  assign n20615 = n19571 & n20614;
  assign n20616 = n19568 & ~n20611;
  assign n20617 = ~n20462 & ~n20540;
  assign n20618 = n20462 & n20540;
  assign n20619 = ~n20552 & ~n20618;
  assign n20620 = ~n20617 & ~n20619;
  assign n20621 = n20533 & ~n20611;
  assign n20622 = ~n20533 & n20611;
  assign n20623 = ~n20621 & ~n20622;
  assign n20624 = n20620 & ~n20623;
  assign n20625 = ~n20620 & n20623;
  assign n20626 = ~n20624 & ~n20625;
  assign n20627 = n19604 & ~n20626;
  assign n20628 = ~n20603 & ~n20615;
  assign n20629 = ~n20616 & n20628;
  assign n20630 = ~n20627 & n20629;
  assign n20631 = ~n20553 & ~n20564;
  assign n20632 = ~n20554 & ~n20631;
  assign n20633 = n20623 & n20632;
  assign n20634 = ~n20623 & ~n20632;
  assign n20635 = ~n20633 & ~n20634;
  assign n20636 = n19627 & ~n20635;
  assign n20637 = n19675 & ~n20462;
  assign n20638 = n19622 & ~n20626;
  assign n20639 = n19625 & ~n20635;
  assign n20640 = ~n20638 & ~n20639;
  assign n20641 = ~n20574 & ~n20618;
  assign n20642 = ~n20617 & ~n20641;
  assign n20643 = ~n20623 & n20642;
  assign n20644 = n20623 & ~n20642;
  assign n20645 = ~n20643 & ~n20644;
  assign n20646 = n19617 & ~n20645;
  assign n20647 = n19611 & ~n20645;
  assign n20648 = n19614 & ~n20635;
  assign n20649 = n19619 & ~n20635;
  assign n20650 = ~n20648 & ~n20649;
  assign n20651 = ~n20646 & ~n20647;
  assign n20652 = n20650 & n20651;
  assign n20653 = ~n20636 & ~n20637;
  assign n20654 = n20640 & n20653;
  assign n20655 = n20652 & n20654;
  assign n20656 = n20630 & n20655;
  assign n20657 = n19554 & ~n20656;
  assign n20658 = P4_REG0_REG_15_ & ~n19554;
  assign n2421 = n20657 | n20658;
  assign n20660 = P4_REG1_REG_17_ & n19585;
  assign n20661 = P4_REG2_REG_17_ & n19587;
  assign n20662 = P4_REG0_REG_17_ & n19583;
  assign n20663 = P4_REG3_REG_16_ & n20595;
  assign n20664 = ~P4_REG3_REG_17_ & n20663;
  assign n20665 = P4_REG3_REG_17_ & ~n20663;
  assign n20666 = ~n20664 & ~n20665;
  assign n20667 = n19581 & ~n20666;
  assign n20668 = ~n20660 & ~n20661;
  assign n20669 = ~n20662 & n20668;
  assign n20670 = ~n20667 & n20669;
  assign n20671 = n19574 & ~n20670;
  assign n20672 = P4_IR_REG_31_ & n19186;
  assign n20673 = P4_IR_REG_16_ & ~P4_IR_REG_31_;
  assign n20674 = ~n20672 & ~n20673;
  assign n20675 = n19561 & ~n20674;
  assign n20676 = P2_P3_DATAO_REG_16_ & ~n19561;
  assign n20677 = ~n20675 & ~n20676;
  assign n20678 = n20612 & n20677;
  assign n20679 = ~n20612 & ~n20677;
  assign n20680 = ~n20678 & ~n20679;
  assign n20681 = n19571 & n20680;
  assign n20682 = n19568 & ~n20677;
  assign n20683 = n20602 & ~n20677;
  assign n20684 = ~n20602 & n20677;
  assign n20685 = ~n20683 & ~n20684;
  assign n20686 = ~n20533 & ~n20611;
  assign n20687 = n20533 & n20611;
  assign n20688 = ~n20620 & ~n20687;
  assign n20689 = ~n20686 & ~n20688;
  assign n20690 = ~n20685 & n20689;
  assign n20691 = n20602 & n20677;
  assign n20692 = ~n20602 & ~n20677;
  assign n20693 = ~n20691 & ~n20692;
  assign n20694 = ~n20689 & ~n20693;
  assign n20695 = ~n20690 & ~n20694;
  assign n20696 = n19604 & ~n20695;
  assign n20697 = ~n20671 & ~n20681;
  assign n20698 = ~n20682 & n20697;
  assign n20699 = ~n20696 & n20698;
  assign n20700 = ~n20621 & ~n20685;
  assign n20701 = ~n20622 & n20632;
  assign n20702 = n20700 & ~n20701;
  assign n20703 = ~n20622 & ~n20684;
  assign n20704 = ~n20683 & n20703;
  assign n20705 = ~n20621 & ~n20632;
  assign n20706 = n20704 & ~n20705;
  assign n20707 = ~n20702 & ~n20706;
  assign n20708 = n19627 & ~n20707;
  assign n20709 = n19675 & ~n20533;
  assign n20710 = n19622 & ~n20695;
  assign n20711 = n19625 & ~n20707;
  assign n20712 = ~n20710 & ~n20711;
  assign n20713 = ~n20642 & ~n20687;
  assign n20714 = ~n20686 & ~n20713;
  assign n20715 = ~n20685 & n20714;
  assign n20716 = ~n20693 & ~n20714;
  assign n20717 = ~n20715 & ~n20716;
  assign n20718 = n19617 & ~n20717;
  assign n20719 = n19611 & ~n20717;
  assign n20720 = n19614 & ~n20707;
  assign n20721 = n19619 & ~n20707;
  assign n20722 = ~n20720 & ~n20721;
  assign n20723 = ~n20718 & ~n20719;
  assign n20724 = n20722 & n20723;
  assign n20725 = ~n20708 & ~n20709;
  assign n20726 = n20712 & n20725;
  assign n20727 = n20724 & n20726;
  assign n20728 = n20699 & n20727;
  assign n20729 = n19554 & ~n20728;
  assign n20730 = P4_REG0_REG_16_ & ~n19554;
  assign n2426 = n20729 | n20730;
  assign n20732 = P4_REG1_REG_18_ & n19585;
  assign n20733 = P4_REG2_REG_18_ & n19587;
  assign n20734 = P4_REG0_REG_18_ & n19583;
  assign n20735 = P4_REG3_REG_17_ & n20663;
  assign n20736 = ~P4_REG3_REG_18_ & n20735;
  assign n20737 = P4_REG3_REG_18_ & ~n20735;
  assign n20738 = ~n20736 & ~n20737;
  assign n20739 = n19581 & ~n20738;
  assign n20740 = ~n20732 & ~n20733;
  assign n20741 = ~n20734 & n20740;
  assign n20742 = ~n20739 & n20741;
  assign n20743 = n19574 & ~n20742;
  assign n20744 = n20611 & n20677;
  assign n20745 = n20605 & n20744;
  assign n20746 = P4_IR_REG_31_ & n19194;
  assign n20747 = P4_IR_REG_17_ & ~P4_IR_REG_31_;
  assign n20748 = ~n20746 & ~n20747;
  assign n20749 = n19561 & ~n20748;
  assign n20750 = P2_P3_DATAO_REG_17_ & ~n19561;
  assign n20751 = ~n20749 & ~n20750;
  assign n20752 = n20745 & n20751;
  assign n20753 = ~n20745 & ~n20751;
  assign n20754 = ~n20752 & ~n20753;
  assign n20755 = n19571 & n20754;
  assign n20756 = n19568 & ~n20751;
  assign n20757 = ~n20670 & ~n20751;
  assign n20758 = n20670 & n20751;
  assign n20759 = ~n20691 & ~n20758;
  assign n20760 = ~n20757 & n20759;
  assign n20761 = n20689 & ~n20692;
  assign n20762 = n20760 & ~n20761;
  assign n20763 = n20670 & ~n20751;
  assign n20764 = ~n20670 & n20751;
  assign n20765 = ~n20763 & ~n20764;
  assign n20766 = ~n20692 & n20765;
  assign n20767 = ~n20689 & ~n20691;
  assign n20768 = n20766 & ~n20767;
  assign n20769 = ~n20762 & ~n20768;
  assign n20770 = n19604 & n20769;
  assign n20771 = ~n20743 & ~n20755;
  assign n20772 = ~n20756 & n20771;
  assign n20773 = ~n20770 & n20772;
  assign n20774 = ~n20621 & ~n20683;
  assign n20775 = n20554 & n20774;
  assign n20776 = n20703 & ~n20775;
  assign n20777 = ~n20683 & ~n20776;
  assign n20778 = ~n20553 & n20774;
  assign n20779 = ~n20564 & n20778;
  assign n20780 = ~n20777 & ~n20779;
  assign n20781 = ~n20765 & ~n20780;
  assign n20782 = n20765 & n20780;
  assign n20783 = ~n20781 & ~n20782;
  assign n20784 = n19627 & ~n20783;
  assign n20785 = n19675 & ~n20602;
  assign n20786 = n19622 & n20769;
  assign n20787 = n19625 & ~n20783;
  assign n20788 = ~n20786 & ~n20787;
  assign n20789 = ~n20692 & n20714;
  assign n20790 = n20760 & ~n20789;
  assign n20791 = ~n20691 & ~n20714;
  assign n20792 = n20766 & ~n20791;
  assign n20793 = ~n20790 & ~n20792;
  assign n20794 = n19617 & n20793;
  assign n20795 = n19611 & n20793;
  assign n20796 = n19614 & ~n20783;
  assign n20797 = n19619 & ~n20783;
  assign n20798 = ~n20796 & ~n20797;
  assign n20799 = ~n20794 & ~n20795;
  assign n20800 = n20798 & n20799;
  assign n20801 = ~n20784 & ~n20785;
  assign n20802 = n20788 & n20801;
  assign n20803 = n20800 & n20802;
  assign n20804 = n20773 & n20803;
  assign n20805 = n19554 & ~n20804;
  assign n20806 = P4_REG0_REG_17_ & ~n19554;
  assign n2431 = n20805 | n20806;
  assign n20808 = P4_REG1_REG_19_ & n19585;
  assign n20809 = P4_REG2_REG_19_ & n19587;
  assign n20810 = P4_REG0_REG_19_ & n19583;
  assign n20811 = P4_REG3_REG_18_ & n20735;
  assign n20812 = ~P4_REG3_REG_19_ & n20811;
  assign n20813 = P4_REG3_REG_19_ & ~n20811;
  assign n20814 = ~n20812 & ~n20813;
  assign n20815 = n19581 & ~n20814;
  assign n20816 = ~n20808 & ~n20809;
  assign n20817 = ~n20810 & n20816;
  assign n20818 = ~n20815 & n20817;
  assign n20819 = n19574 & ~n20818;
  assign n20820 = P4_IR_REG_31_ & n19203;
  assign n20821 = P4_IR_REG_18_ & ~P4_IR_REG_31_;
  assign n20822 = ~n20820 & ~n20821;
  assign n20823 = n19561 & ~n20822;
  assign n20824 = P2_P3_DATAO_REG_18_ & ~n19561;
  assign n20825 = ~n20823 & ~n20824;
  assign n20826 = n20752 & n20825;
  assign n20827 = ~n20752 & ~n20825;
  assign n20828 = ~n20826 & ~n20827;
  assign n20829 = n19571 & n20828;
  assign n20830 = n19568 & ~n20825;
  assign n20831 = n20692 & ~n20751;
  assign n20832 = ~n20692 & n20751;
  assign n20833 = ~n20670 & ~n20832;
  assign n20834 = ~n20831 & ~n20833;
  assign n20835 = ~n20689 & n20759;
  assign n20836 = n20834 & ~n20835;
  assign n20837 = n20742 & ~n20825;
  assign n20838 = ~n20742 & n20825;
  assign n20839 = ~n20837 & ~n20838;
  assign n20840 = n20836 & ~n20839;
  assign n20841 = n20742 & n20825;
  assign n20842 = ~n20742 & ~n20825;
  assign n20843 = ~n20841 & ~n20842;
  assign n20844 = ~n20836 & ~n20843;
  assign n20845 = ~n20840 & ~n20844;
  assign n20846 = n19604 & ~n20845;
  assign n20847 = ~n20819 & ~n20829;
  assign n20848 = ~n20830 & n20847;
  assign n20849 = ~n20846 & n20848;
  assign n20850 = ~n20763 & ~n20780;
  assign n20851 = ~n20764 & ~n20850;
  assign n20852 = ~n20839 & ~n20851;
  assign n20853 = n20839 & n20851;
  assign n20854 = ~n20852 & ~n20853;
  assign n20855 = n19627 & ~n20854;
  assign n20856 = n19675 & ~n20670;
  assign n20857 = n19622 & ~n20845;
  assign n20858 = n19625 & ~n20854;
  assign n20859 = ~n20857 & ~n20858;
  assign n20860 = ~n20714 & n20759;
  assign n20861 = n20834 & ~n20860;
  assign n20862 = ~n20839 & n20861;
  assign n20863 = ~n20843 & ~n20861;
  assign n20864 = ~n20862 & ~n20863;
  assign n20865 = n19617 & ~n20864;
  assign n20866 = n19611 & ~n20864;
  assign n20867 = n19614 & ~n20854;
  assign n20868 = n19619 & ~n20854;
  assign n20869 = ~n20867 & ~n20868;
  assign n20870 = ~n20865 & ~n20866;
  assign n20871 = n20869 & n20870;
  assign n20872 = ~n20855 & ~n20856;
  assign n20873 = n20859 & n20872;
  assign n20874 = n20871 & n20873;
  assign n20875 = n20849 & n20874;
  assign n20876 = n19554 & ~n20875;
  assign n20877 = P4_REG0_REG_18_ & ~n19554;
  assign n2436 = n20876 | n20877;
  assign n20879 = P4_REG1_REG_20_ & n19585;
  assign n20880 = P4_REG2_REG_20_ & n19587;
  assign n20881 = P4_REG0_REG_20_ & n19583;
  assign n20882 = P4_REG3_REG_19_ & n20811;
  assign n20883 = ~P4_REG3_REG_20_ & n20882;
  assign n20884 = P4_REG3_REG_20_ & ~n20882;
  assign n20885 = ~n20883 & ~n20884;
  assign n20886 = n19581 & ~n20885;
  assign n20887 = ~n20879 & ~n20880;
  assign n20888 = ~n20881 & n20887;
  assign n20889 = ~n20886 & n20888;
  assign n20890 = n19574 & ~n20889;
  assign n20891 = n20751 & n20825;
  assign n20892 = n20745 & n20891;
  assign n20893 = ~n19479 & n19561;
  assign n20894 = P2_P3_DATAO_REG_19_ & ~n19561;
  assign n20895 = ~n20893 & ~n20894;
  assign n20896 = n20892 & n20895;
  assign n20897 = ~n20892 & ~n20895;
  assign n20898 = ~n20896 & ~n20897;
  assign n20899 = n19571 & n20898;
  assign n20900 = n19568 & ~n20895;
  assign n20901 = n20818 & ~n20895;
  assign n20902 = ~n20818 & n20895;
  assign n20903 = ~n20901 & ~n20902;
  assign n20904 = ~n20836 & ~n20841;
  assign n20905 = ~n20842 & ~n20904;
  assign n20906 = ~n20903 & n20905;
  assign n20907 = n20818 & n20895;
  assign n20908 = ~n20818 & ~n20895;
  assign n20909 = ~n20907 & ~n20908;
  assign n20910 = ~n20905 & ~n20909;
  assign n20911 = ~n20906 & ~n20910;
  assign n20912 = n19604 & ~n20911;
  assign n20913 = ~n20890 & ~n20899;
  assign n20914 = ~n20900 & n20913;
  assign n20915 = ~n20912 & n20914;
  assign n20916 = ~n20742 & ~n20851;
  assign n20917 = n20825 & ~n20851;
  assign n20918 = ~n20916 & ~n20917;
  assign n20919 = ~n20838 & n20918;
  assign n20920 = ~n20903 & ~n20919;
  assign n20921 = n20903 & n20919;
  assign n20922 = ~n20920 & ~n20921;
  assign n20923 = n19627 & ~n20922;
  assign n20924 = n19675 & ~n20742;
  assign n20925 = n19622 & ~n20911;
  assign n20926 = n19625 & ~n20922;
  assign n20927 = ~n20925 & ~n20926;
  assign n20928 = ~n20841 & ~n20861;
  assign n20929 = ~n20842 & ~n20928;
  assign n20930 = ~n20903 & n20929;
  assign n20931 = ~n20909 & ~n20929;
  assign n20932 = ~n20930 & ~n20931;
  assign n20933 = n19617 & ~n20932;
  assign n20934 = n19611 & ~n20932;
  assign n20935 = n19614 & ~n20922;
  assign n20936 = n19619 & ~n20922;
  assign n20937 = ~n20935 & ~n20936;
  assign n20938 = ~n20933 & ~n20934;
  assign n20939 = n20937 & n20938;
  assign n20940 = ~n20923 & ~n20924;
  assign n20941 = n20927 & n20940;
  assign n20942 = n20939 & n20941;
  assign n20943 = n20915 & n20942;
  assign n20944 = n19554 & ~n20943;
  assign n20945 = P4_REG0_REG_19_ & ~n19554;
  assign n2441 = n20944 | n20945;
  assign n20947 = P4_REG1_REG_21_ & n19585;
  assign n20948 = P4_REG2_REG_21_ & n19587;
  assign n20949 = P4_REG0_REG_21_ & n19583;
  assign n20950 = P4_REG3_REG_20_ & n20882;
  assign n20951 = ~P4_REG3_REG_21_ & n20950;
  assign n20952 = P4_REG3_REG_21_ & ~n20950;
  assign n20953 = ~n20951 & ~n20952;
  assign n20954 = n19581 & ~n20953;
  assign n20955 = ~n20947 & ~n20948;
  assign n20956 = ~n20949 & n20955;
  assign n20957 = ~n20954 & n20956;
  assign n20958 = n19574 & ~n20957;
  assign n20959 = P2_P3_DATAO_REG_20_ & ~n19561;
  assign n20960 = n20896 & ~n20959;
  assign n20961 = ~n20896 & n20959;
  assign n20962 = ~n20960 & ~n20961;
  assign n20963 = n19571 & n20962;
  assign n20964 = n19568 & n20959;
  assign n20965 = ~n20889 & n20959;
  assign n20966 = n20889 & ~n20959;
  assign n20967 = ~n20907 & ~n20966;
  assign n20968 = ~n20965 & n20967;
  assign n20969 = n20905 & ~n20908;
  assign n20970 = n20968 & ~n20969;
  assign n20971 = n20889 & n20959;
  assign n20972 = ~n20889 & ~n20959;
  assign n20973 = ~n20971 & ~n20972;
  assign n20974 = ~n20908 & n20973;
  assign n20975 = ~n20905 & ~n20907;
  assign n20976 = n20974 & ~n20975;
  assign n20977 = ~n20970 & ~n20976;
  assign n20978 = n19604 & n20977;
  assign n20979 = ~n20958 & ~n20963;
  assign n20980 = ~n20964 & n20979;
  assign n20981 = ~n20978 & n20980;
  assign n20982 = ~n20901 & ~n20919;
  assign n20983 = ~n20902 & ~n20982;
  assign n20984 = ~n20973 & ~n20983;
  assign n20985 = n20973 & n20983;
  assign n20986 = ~n20984 & ~n20985;
  assign n20987 = n19627 & ~n20986;
  assign n20988 = n19675 & ~n20818;
  assign n20989 = n19622 & n20977;
  assign n20990 = n19625 & ~n20986;
  assign n20991 = ~n20989 & ~n20990;
  assign n20992 = ~n20908 & n20929;
  assign n20993 = n20968 & ~n20992;
  assign n20994 = ~n20907 & ~n20929;
  assign n20995 = n20974 & ~n20994;
  assign n20996 = ~n20993 & ~n20995;
  assign n20997 = n19617 & n20996;
  assign n20998 = n19611 & n20996;
  assign n20999 = n19614 & ~n20986;
  assign n21000 = n19619 & ~n20986;
  assign n21001 = ~n20999 & ~n21000;
  assign n21002 = ~n20997 & ~n20998;
  assign n21003 = n21001 & n21002;
  assign n21004 = ~n20987 & ~n20988;
  assign n21005 = n20991 & n21004;
  assign n21006 = n21003 & n21005;
  assign n21007 = n20981 & n21006;
  assign n21008 = n19554 & ~n21007;
  assign n21009 = P4_REG0_REG_20_ & ~n19554;
  assign n2446 = n21008 | n21009;
  assign n21011 = P4_REG1_REG_22_ & n19585;
  assign n21012 = P4_REG2_REG_22_ & n19587;
  assign n21013 = P4_REG0_REG_22_ & n19583;
  assign n21014 = P4_REG3_REG_21_ & n20950;
  assign n21015 = ~P4_REG3_REG_22_ & n21014;
  assign n21016 = P4_REG3_REG_22_ & ~n21014;
  assign n21017 = ~n21015 & ~n21016;
  assign n21018 = n19581 & ~n21017;
  assign n21019 = ~n21011 & ~n21012;
  assign n21020 = ~n21013 & n21019;
  assign n21021 = ~n21018 & n21020;
  assign n21022 = n19574 & ~n21021;
  assign n21023 = n20895 & ~n20959;
  assign n21024 = n20892 & n21023;
  assign n21025 = P2_P3_DATAO_REG_21_ & ~n19561;
  assign n21026 = n21024 & ~n21025;
  assign n21027 = ~n21024 & n21025;
  assign n21028 = ~n21026 & ~n21027;
  assign n21029 = n19571 & n21028;
  assign n21030 = n19568 & n21025;
  assign n21031 = n20957 & n21025;
  assign n21032 = ~n20957 & ~n21025;
  assign n21033 = ~n21031 & ~n21032;
  assign n21034 = ~n20905 & n20967;
  assign n21035 = ~n20908 & ~n20959;
  assign n21036 = n20908 & n20959;
  assign n21037 = n20889 & ~n21036;
  assign n21038 = ~n21035 & ~n21037;
  assign n21039 = ~n21034 & ~n21038;
  assign n21040 = ~n21033 & ~n21039;
  assign n21041 = n21033 & ~n21038;
  assign n21042 = ~n21034 & n21041;
  assign n21043 = ~n21040 & ~n21042;
  assign n21044 = n19604 & n21043;
  assign n21045 = ~n21022 & ~n21029;
  assign n21046 = ~n21030 & n21045;
  assign n21047 = ~n21044 & n21046;
  assign n21048 = ~n20971 & ~n20983;
  assign n21049 = ~n20972 & ~n21048;
  assign n21050 = n21033 & n21049;
  assign n21051 = ~n21033 & ~n21049;
  assign n21052 = ~n21050 & ~n21051;
  assign n21053 = n19627 & ~n21052;
  assign n21054 = n19675 & ~n20889;
  assign n21055 = n19622 & n21043;
  assign n21056 = n19625 & ~n21052;
  assign n21057 = ~n21055 & ~n21056;
  assign n21058 = ~n20929 & n20967;
  assign n21059 = ~n21038 & ~n21058;
  assign n21060 = ~n21033 & ~n21059;
  assign n21061 = n21041 & ~n21058;
  assign n21062 = ~n21060 & ~n21061;
  assign n21063 = n19617 & n21062;
  assign n21064 = n19611 & n21062;
  assign n21065 = n19614 & ~n21052;
  assign n21066 = n19619 & ~n21052;
  assign n21067 = ~n21065 & ~n21066;
  assign n21068 = ~n21063 & ~n21064;
  assign n21069 = n21067 & n21068;
  assign n21070 = ~n21053 & ~n21054;
  assign n21071 = n21057 & n21070;
  assign n21072 = n21069 & n21071;
  assign n21073 = n21047 & n21072;
  assign n21074 = n19554 & ~n21073;
  assign n21075 = P4_REG0_REG_21_ & ~n19554;
  assign n2451 = n21074 | n21075;
  assign n21077 = P4_REG1_REG_23_ & n19585;
  assign n21078 = P4_REG2_REG_23_ & n19587;
  assign n21079 = P4_REG0_REG_23_ & n19583;
  assign n21080 = P4_REG3_REG_22_ & n21014;
  assign n21081 = ~P4_REG3_REG_23_ & n21080;
  assign n21082 = P4_REG3_REG_23_ & ~n21080;
  assign n21083 = ~n21081 & ~n21082;
  assign n21084 = n19581 & ~n21083;
  assign n21085 = ~n21077 & ~n21078;
  assign n21086 = ~n21079 & n21085;
  assign n21087 = ~n21084 & n21086;
  assign n21088 = n19574 & ~n21087;
  assign n21089 = P2_P3_DATAO_REG_22_ & ~n19561;
  assign n21090 = n21026 & ~n21089;
  assign n21091 = ~n21026 & n21089;
  assign n21092 = ~n21090 & ~n21091;
  assign n21093 = n19571 & n21092;
  assign n21094 = n19568 & n21089;
  assign n21095 = n20957 & ~n21025;
  assign n21096 = n20842 & n20967;
  assign n21097 = ~n21038 & ~n21096;
  assign n21098 = ~n21095 & ~n21097;
  assign n21099 = ~n20957 & n21025;
  assign n21100 = ~n21098 & ~n21099;
  assign n21101 = ~n20841 & n20967;
  assign n21102 = ~n21095 & n21101;
  assign n21103 = ~n20836 & n21102;
  assign n21104 = n21100 & ~n21103;
  assign n21105 = n21021 & n21089;
  assign n21106 = ~n21021 & ~n21089;
  assign n21107 = ~n21105 & ~n21106;
  assign n21108 = n21104 & ~n21107;
  assign n21109 = ~n21104 & n21107;
  assign n21110 = ~n21108 & ~n21109;
  assign n21111 = n19604 & ~n21110;
  assign n21112 = ~n21088 & ~n21093;
  assign n21113 = ~n21094 & n21112;
  assign n21114 = ~n21111 & n21113;
  assign n21115 = ~n21031 & ~n21049;
  assign n21116 = ~n21032 & ~n21115;
  assign n21117 = n21107 & n21116;
  assign n21118 = ~n21107 & ~n21116;
  assign n21119 = ~n21117 & ~n21118;
  assign n21120 = n19627 & ~n21119;
  assign n21121 = n19675 & ~n20957;
  assign n21122 = n19622 & ~n21110;
  assign n21123 = n19625 & ~n21119;
  assign n21124 = ~n21122 & ~n21123;
  assign n21125 = ~n20861 & n21102;
  assign n21126 = n21100 & ~n21125;
  assign n21127 = ~n21107 & n21126;
  assign n21128 = n21107 & ~n21126;
  assign n21129 = ~n21127 & ~n21128;
  assign n21130 = n19617 & ~n21129;
  assign n21131 = n19611 & ~n21129;
  assign n21132 = n19614 & ~n21119;
  assign n21133 = n19619 & ~n21119;
  assign n21134 = ~n21132 & ~n21133;
  assign n21135 = ~n21130 & ~n21131;
  assign n21136 = n21134 & n21135;
  assign n21137 = ~n21120 & ~n21121;
  assign n21138 = n21124 & n21137;
  assign n21139 = n21136 & n21138;
  assign n21140 = n21114 & n21139;
  assign n21141 = n19554 & ~n21140;
  assign n21142 = P4_REG0_REG_22_ & ~n19554;
  assign n2456 = n21141 | n21142;
  assign n21144 = P4_REG1_REG_24_ & n19585;
  assign n21145 = P4_REG2_REG_24_ & n19587;
  assign n21146 = P4_REG0_REG_24_ & n19583;
  assign n21147 = P4_REG3_REG_23_ & n21080;
  assign n21148 = ~P4_REG3_REG_24_ & n21147;
  assign n21149 = P4_REG3_REG_24_ & ~n21147;
  assign n21150 = ~n21148 & ~n21149;
  assign n21151 = n19581 & ~n21150;
  assign n21152 = ~n21144 & ~n21145;
  assign n21153 = ~n21146 & n21152;
  assign n21154 = ~n21151 & n21153;
  assign n21155 = n19574 & ~n21154;
  assign n21156 = ~n21025 & ~n21089;
  assign n21157 = n21024 & n21156;
  assign n21158 = P2_P3_DATAO_REG_23_ & ~n19561;
  assign n21159 = n21157 & ~n21158;
  assign n21160 = ~n21157 & n21158;
  assign n21161 = ~n21159 & ~n21160;
  assign n21162 = n19571 & n21161;
  assign n21163 = n19568 & n21158;
  assign n21164 = ~n21021 & n21089;
  assign n21165 = n21021 & ~n21089;
  assign n21166 = ~n21104 & ~n21165;
  assign n21167 = ~n21164 & ~n21166;
  assign n21168 = n21087 & n21158;
  assign n21169 = ~n21087 & ~n21158;
  assign n21170 = ~n21168 & ~n21169;
  assign n21171 = n21167 & ~n21170;
  assign n21172 = ~n21167 & n21170;
  assign n21173 = ~n21171 & ~n21172;
  assign n21174 = n19604 & ~n21173;
  assign n21175 = ~n21155 & ~n21162;
  assign n21176 = ~n21163 & n21175;
  assign n21177 = ~n21174 & n21176;
  assign n21178 = ~n21105 & ~n21170;
  assign n21179 = ~n21106 & n21116;
  assign n21180 = n21178 & ~n21179;
  assign n21181 = ~n21106 & ~n21169;
  assign n21182 = ~n21168 & n21181;
  assign n21183 = ~n21105 & ~n21116;
  assign n21184 = n21182 & ~n21183;
  assign n21185 = ~n21180 & ~n21184;
  assign n21186 = n19627 & ~n21185;
  assign n21187 = n19675 & ~n21021;
  assign n21188 = n19622 & ~n21173;
  assign n21189 = n19625 & ~n21185;
  assign n21190 = ~n21188 & ~n21189;
  assign n21191 = ~n21126 & ~n21165;
  assign n21192 = ~n21164 & ~n21191;
  assign n21193 = ~n21170 & n21192;
  assign n21194 = n21170 & ~n21192;
  assign n21195 = ~n21193 & ~n21194;
  assign n21196 = n19617 & ~n21195;
  assign n21197 = n19611 & ~n21195;
  assign n21198 = n19614 & ~n21185;
  assign n21199 = n19619 & ~n21185;
  assign n21200 = ~n21198 & ~n21199;
  assign n21201 = ~n21196 & ~n21197;
  assign n21202 = n21200 & n21201;
  assign n21203 = ~n21186 & ~n21187;
  assign n21204 = n21190 & n21203;
  assign n21205 = n21202 & n21204;
  assign n21206 = n21177 & n21205;
  assign n21207 = n19554 & ~n21206;
  assign n21208 = P4_REG0_REG_23_ & ~n19554;
  assign n2461 = n21207 | n21208;
  assign n21210 = P4_REG1_REG_25_ & n19585;
  assign n21211 = P4_REG2_REG_25_ & n19587;
  assign n21212 = P4_REG0_REG_25_ & n19583;
  assign n21213 = P4_REG3_REG_24_ & n21147;
  assign n21214 = ~P4_REG3_REG_25_ & n21213;
  assign n21215 = P4_REG3_REG_25_ & ~n21213;
  assign n21216 = ~n21214 & ~n21215;
  assign n21217 = n19581 & ~n21216;
  assign n21218 = ~n21210 & ~n21211;
  assign n21219 = ~n21212 & n21218;
  assign n21220 = ~n21217 & n21219;
  assign n21221 = n19574 & ~n21220;
  assign n21222 = P2_P3_DATAO_REG_24_ & ~n19561;
  assign n21223 = n21159 & ~n21222;
  assign n21224 = ~n21159 & n21222;
  assign n21225 = ~n21223 & ~n21224;
  assign n21226 = n19571 & n21225;
  assign n21227 = n19568 & n21222;
  assign n21228 = ~n21087 & n21158;
  assign n21229 = n21087 & ~n21158;
  assign n21230 = ~n21167 & ~n21229;
  assign n21231 = ~n21228 & ~n21230;
  assign n21232 = n21154 & n21222;
  assign n21233 = ~n21154 & ~n21222;
  assign n21234 = ~n21232 & ~n21233;
  assign n21235 = n21231 & ~n21234;
  assign n21236 = n21154 & ~n21222;
  assign n21237 = ~n21154 & n21222;
  assign n21238 = ~n21236 & ~n21237;
  assign n21239 = ~n21231 & ~n21238;
  assign n21240 = ~n21235 & ~n21239;
  assign n21241 = n19604 & ~n21240;
  assign n21242 = ~n21221 & ~n21226;
  assign n21243 = ~n21227 & n21242;
  assign n21244 = ~n21241 & n21243;
  assign n21245 = ~n21105 & ~n21168;
  assign n21246 = n21032 & n21245;
  assign n21247 = n21181 & ~n21246;
  assign n21248 = ~n21168 & ~n21247;
  assign n21249 = ~n21031 & n21245;
  assign n21250 = ~n21049 & n21249;
  assign n21251 = ~n21248 & ~n21250;
  assign n21252 = ~n21234 & ~n21251;
  assign n21253 = n21234 & n21251;
  assign n21254 = ~n21252 & ~n21253;
  assign n21255 = n19627 & ~n21254;
  assign n21256 = n19675 & ~n21087;
  assign n21257 = n19622 & ~n21240;
  assign n21258 = n19625 & ~n21254;
  assign n21259 = ~n21257 & ~n21258;
  assign n21260 = ~n21192 & ~n21229;
  assign n21261 = ~n21228 & ~n21260;
  assign n21262 = ~n21234 & n21261;
  assign n21263 = ~n21238 & ~n21261;
  assign n21264 = ~n21262 & ~n21263;
  assign n21265 = n19617 & ~n21264;
  assign n21266 = n19611 & ~n21264;
  assign n21267 = n19614 & ~n21254;
  assign n21268 = n19619 & ~n21254;
  assign n21269 = ~n21267 & ~n21268;
  assign n21270 = ~n21265 & ~n21266;
  assign n21271 = n21269 & n21270;
  assign n21272 = ~n21255 & ~n21256;
  assign n21273 = n21259 & n21272;
  assign n21274 = n21271 & n21273;
  assign n21275 = n21244 & n21274;
  assign n21276 = n19554 & ~n21275;
  assign n21277 = P4_REG0_REG_24_ & ~n19554;
  assign n2466 = n21276 | n21277;
  assign n21279 = P4_REG1_REG_26_ & n19585;
  assign n21280 = P4_REG2_REG_26_ & n19587;
  assign n21281 = P4_REG0_REG_26_ & n19583;
  assign n21282 = P4_REG3_REG_25_ & n21213;
  assign n21283 = ~P4_REG3_REG_26_ & n21282;
  assign n21284 = P4_REG3_REG_26_ & ~n21282;
  assign n21285 = ~n21283 & ~n21284;
  assign n21286 = n19581 & ~n21285;
  assign n21287 = ~n21279 & ~n21280;
  assign n21288 = ~n21281 & n21287;
  assign n21289 = ~n21286 & n21288;
  assign n21290 = n19574 & ~n21289;
  assign n21291 = ~n21158 & ~n21222;
  assign n21292 = n21157 & n21291;
  assign n21293 = P2_P3_DATAO_REG_25_ & ~n19561;
  assign n21294 = n21292 & ~n21293;
  assign n21295 = ~n21292 & n21293;
  assign n21296 = ~n21294 & ~n21295;
  assign n21297 = n19571 & n21296;
  assign n21298 = n19568 & n21293;
  assign n21299 = n21220 & n21293;
  assign n21300 = ~n21220 & ~n21293;
  assign n21301 = ~n21299 & ~n21300;
  assign n21302 = ~n21231 & ~n21236;
  assign n21303 = ~n21237 & ~n21302;
  assign n21304 = ~n21301 & n21303;
  assign n21305 = n21220 & ~n21293;
  assign n21306 = ~n21220 & n21293;
  assign n21307 = ~n21305 & ~n21306;
  assign n21308 = ~n21303 & ~n21307;
  assign n21309 = ~n21304 & ~n21308;
  assign n21310 = n19604 & ~n21309;
  assign n21311 = ~n21290 & ~n21297;
  assign n21312 = ~n21298 & n21311;
  assign n21313 = ~n21310 & n21312;
  assign n21314 = ~n21232 & ~n21251;
  assign n21315 = ~n21233 & ~n21314;
  assign n21316 = ~n21301 & ~n21315;
  assign n21317 = n21301 & n21315;
  assign n21318 = ~n21316 & ~n21317;
  assign n21319 = n19627 & ~n21318;
  assign n21320 = n19675 & ~n21154;
  assign n21321 = n19622 & ~n21309;
  assign n21322 = n19625 & ~n21318;
  assign n21323 = ~n21321 & ~n21322;
  assign n21324 = ~n21236 & ~n21261;
  assign n21325 = ~n21237 & ~n21324;
  assign n21326 = ~n21301 & n21325;
  assign n21327 = ~n21307 & ~n21325;
  assign n21328 = ~n21326 & ~n21327;
  assign n21329 = n19617 & ~n21328;
  assign n21330 = n19611 & ~n21328;
  assign n21331 = n19614 & ~n21318;
  assign n21332 = n19619 & ~n21318;
  assign n21333 = ~n21331 & ~n21332;
  assign n21334 = ~n21329 & ~n21330;
  assign n21335 = n21333 & n21334;
  assign n21336 = ~n21319 & ~n21320;
  assign n21337 = n21323 & n21336;
  assign n21338 = n21335 & n21337;
  assign n21339 = n21313 & n21338;
  assign n21340 = n19554 & ~n21339;
  assign n21341 = P4_REG0_REG_25_ & ~n19554;
  assign n2471 = n21340 | n21341;
  assign n21343 = P4_REG1_REG_27_ & n19585;
  assign n21344 = P4_REG2_REG_27_ & n19587;
  assign n21345 = P4_REG0_REG_27_ & n19583;
  assign n21346 = P4_REG3_REG_26_ & n21282;
  assign n21347 = ~P4_REG3_REG_27_ & n21346;
  assign n21348 = P4_REG3_REG_27_ & ~n21346;
  assign n21349 = ~n21347 & ~n21348;
  assign n21350 = n19581 & ~n21349;
  assign n21351 = ~n21343 & ~n21344;
  assign n21352 = ~n21345 & n21351;
  assign n21353 = ~n21350 & n21352;
  assign n21354 = n19574 & ~n21353;
  assign n21355 = P2_P3_DATAO_REG_26_ & ~n19561;
  assign n21356 = n21294 & ~n21355;
  assign n21357 = ~n21294 & n21355;
  assign n21358 = ~n21356 & ~n21357;
  assign n21359 = n19571 & n21358;
  assign n21360 = n19568 & n21355;
  assign n21361 = n21303 & ~n21306;
  assign n21362 = ~n21289 & n21355;
  assign n21363 = ~n21305 & n21355;
  assign n21364 = ~n21289 & ~n21305;
  assign n21365 = ~n21363 & ~n21364;
  assign n21366 = ~n21361 & ~n21362;
  assign n21367 = ~n21365 & n21366;
  assign n21368 = ~n21303 & ~n21305;
  assign n21369 = n21289 & n21355;
  assign n21370 = ~n21289 & ~n21355;
  assign n21371 = ~n21369 & ~n21370;
  assign n21372 = ~n21306 & ~n21368;
  assign n21373 = n21371 & n21372;
  assign n21374 = ~n21367 & ~n21373;
  assign n21375 = n19604 & n21374;
  assign n21376 = ~n21354 & ~n21359;
  assign n21377 = ~n21360 & n21376;
  assign n21378 = ~n21375 & n21377;
  assign n21379 = ~n21299 & ~n21315;
  assign n21380 = ~n21300 & ~n21379;
  assign n21381 = n21371 & n21380;
  assign n21382 = ~n21371 & ~n21380;
  assign n21383 = ~n21381 & ~n21382;
  assign n21384 = n19627 & ~n21383;
  assign n21385 = n19675 & ~n21220;
  assign n21386 = n19622 & n21374;
  assign n21387 = n19625 & ~n21383;
  assign n21388 = ~n21386 & ~n21387;
  assign n21389 = ~n21306 & n21325;
  assign n21390 = ~n21362 & ~n21389;
  assign n21391 = ~n21365 & n21390;
  assign n21392 = ~n21305 & ~n21325;
  assign n21393 = ~n21306 & ~n21392;
  assign n21394 = n21371 & n21393;
  assign n21395 = ~n21391 & ~n21394;
  assign n21396 = n19617 & n21395;
  assign n21397 = n19611 & n21395;
  assign n21398 = n19614 & ~n21383;
  assign n21399 = n19619 & ~n21383;
  assign n21400 = ~n21398 & ~n21399;
  assign n21401 = ~n21396 & ~n21397;
  assign n21402 = n21400 & n21401;
  assign n21403 = ~n21384 & ~n21385;
  assign n21404 = n21388 & n21403;
  assign n21405 = n21402 & n21404;
  assign n21406 = n21378 & n21405;
  assign n21407 = n19554 & ~n21406;
  assign n21408 = P4_REG0_REG_26_ & ~n19554;
  assign n2476 = n21407 | n21408;
  assign n21410 = P4_REG1_REG_28_ & n19585;
  assign n21411 = P4_REG2_REG_28_ & n19587;
  assign n21412 = P4_REG0_REG_28_ & n19583;
  assign n21413 = P4_REG3_REG_27_ & n21346;
  assign n21414 = ~P4_REG3_REG_28_ & n21413;
  assign n21415 = P4_REG3_REG_28_ & ~n21413;
  assign n21416 = ~n21414 & ~n21415;
  assign n21417 = n19581 & ~n21416;
  assign n21418 = ~n21410 & ~n21411;
  assign n21419 = ~n21412 & n21418;
  assign n21420 = ~n21417 & n21419;
  assign n21421 = n19574 & ~n21420;
  assign n21422 = P2_P3_DATAO_REG_27_ & ~n19561;
  assign n21423 = n21356 & ~n21422;
  assign n21424 = ~n21356 & n21422;
  assign n21425 = ~n21423 & ~n21424;
  assign n21426 = n19571 & n21425;
  assign n21427 = n19568 & n21422;
  assign n21428 = ~n21237 & ~n21306;
  assign n21429 = ~n21365 & ~n21428;
  assign n21430 = n21302 & ~n21365;
  assign n21431 = ~n21429 & ~n21430;
  assign n21432 = ~n21362 & n21431;
  assign n21433 = n21353 & n21422;
  assign n21434 = ~n21353 & ~n21422;
  assign n21435 = ~n21433 & ~n21434;
  assign n21436 = n21432 & ~n21435;
  assign n21437 = ~n21432 & n21435;
  assign n21438 = ~n21436 & ~n21437;
  assign n21439 = n19604 & ~n21438;
  assign n21440 = ~n21421 & ~n21426;
  assign n21441 = ~n21427 & n21440;
  assign n21442 = ~n21439 & n21441;
  assign n21443 = ~n21369 & ~n21435;
  assign n21444 = ~n21370 & n21380;
  assign n21445 = n21443 & ~n21444;
  assign n21446 = ~n21370 & n21435;
  assign n21447 = ~n21369 & ~n21380;
  assign n21448 = n21446 & ~n21447;
  assign n21449 = ~n21445 & ~n21448;
  assign n21450 = n19627 & ~n21449;
  assign n21451 = n19675 & ~n21289;
  assign n21452 = n19622 & ~n21438;
  assign n21453 = n19625 & ~n21449;
  assign n21454 = ~n21452 & ~n21453;
  assign n21455 = n21324 & ~n21365;
  assign n21456 = ~n21429 & ~n21455;
  assign n21457 = ~n21362 & n21456;
  assign n21458 = ~n21435 & n21457;
  assign n21459 = n21435 & ~n21457;
  assign n21460 = ~n21458 & ~n21459;
  assign n21461 = n19617 & ~n21460;
  assign n21462 = n19611 & ~n21460;
  assign n21463 = n19614 & ~n21449;
  assign n21464 = n19619 & ~n21449;
  assign n21465 = ~n21463 & ~n21464;
  assign n21466 = ~n21461 & ~n21462;
  assign n21467 = n21465 & n21466;
  assign n21468 = ~n21450 & ~n21451;
  assign n21469 = n21454 & n21468;
  assign n21470 = n21467 & n21469;
  assign n21471 = n21442 & n21470;
  assign n21472 = n19554 & ~n21471;
  assign n21473 = P4_REG0_REG_27_ & ~n19554;
  assign n2481 = n21472 | n21473;
  assign n21475 = P4_REG0_REG_29_ & n19583;
  assign n21476 = P4_REG1_REG_29_ & n19585;
  assign n21477 = P4_REG2_REG_29_ & n19587;
  assign n21478 = P4_REG3_REG_28_ & P4_REG3_REG_27_;
  assign n21479 = n21346 & n21478;
  assign n21480 = n19581 & n21479;
  assign n21481 = ~n21475 & ~n21476;
  assign n21482 = ~n21477 & n21481;
  assign n21483 = ~n21480 & n21482;
  assign n21484 = n19574 & ~n21483;
  assign n21485 = P2_P3_DATAO_REG_28_ & ~n19561;
  assign n21486 = n21423 & ~n21485;
  assign n21487 = ~n21423 & n21485;
  assign n21488 = ~n21486 & ~n21487;
  assign n21489 = n19571 & n21488;
  assign n21490 = n19568 & n21485;
  assign n21491 = n21353 & ~n21422;
  assign n21492 = n21362 & ~n21491;
  assign n21493 = ~n21236 & ~n21491;
  assign n21494 = ~n21231 & ~n21365;
  assign n21495 = n21493 & n21494;
  assign n21496 = n21429 & ~n21491;
  assign n21497 = ~n21353 & n21422;
  assign n21498 = ~n21496 & ~n21497;
  assign n21499 = ~n21492 & ~n21495;
  assign n21500 = n21498 & n21499;
  assign n21501 = n21420 & n21485;
  assign n21502 = ~n21420 & ~n21485;
  assign n21503 = ~n21501 & ~n21502;
  assign n21504 = n21500 & ~n21503;
  assign n21505 = ~n21500 & n21503;
  assign n21506 = ~n21504 & ~n21505;
  assign n21507 = n19604 & ~n21506;
  assign n21508 = ~n21484 & ~n21489;
  assign n21509 = ~n21490 & n21508;
  assign n21510 = ~n21507 & n21509;
  assign n21511 = n21353 & ~n21370;
  assign n21512 = ~n21422 & ~n21511;
  assign n21513 = ~n21353 & n21370;
  assign n21514 = ~n21512 & ~n21513;
  assign n21515 = ~n21369 & ~n21433;
  assign n21516 = ~n21380 & n21515;
  assign n21517 = n21514 & ~n21516;
  assign n21518 = ~n21503 & ~n21517;
  assign n21519 = n21503 & n21517;
  assign n21520 = ~n21518 & ~n21519;
  assign n21521 = n19627 & ~n21520;
  assign n21522 = n19675 & ~n21353;
  assign n21523 = n19622 & ~n21506;
  assign n21524 = n19625 & ~n21520;
  assign n21525 = ~n21523 & ~n21524;
  assign n21526 = ~n21261 & ~n21365;
  assign n21527 = n21493 & n21526;
  assign n21528 = ~n21492 & ~n21527;
  assign n21529 = n21498 & n21528;
  assign n21530 = ~n21503 & n21529;
  assign n21531 = n21503 & ~n21529;
  assign n21532 = ~n21530 & ~n21531;
  assign n21533 = n19617 & ~n21532;
  assign n21534 = n19611 & ~n21532;
  assign n21535 = n19614 & ~n21520;
  assign n21536 = n19619 & ~n21520;
  assign n21537 = ~n21535 & ~n21536;
  assign n21538 = ~n21533 & ~n21534;
  assign n21539 = n21537 & n21538;
  assign n21540 = ~n21521 & ~n21522;
  assign n21541 = n21525 & n21540;
  assign n21542 = n21539 & n21541;
  assign n21543 = n21510 & n21542;
  assign n21544 = n19554 & ~n21543;
  assign n21545 = P4_REG0_REG_28_ & ~n19554;
  assign n2486 = n21544 | n21545;
  assign n21547 = P2_P3_DATAO_REG_29_ & ~n19561;
  assign n21548 = n21486 & ~n21547;
  assign n21549 = ~n21486 & n21547;
  assign n21550 = ~n21548 & ~n21549;
  assign n21551 = n19571 & n21550;
  assign n21552 = n19568 & n21547;
  assign n21553 = n21485 & ~n21500;
  assign n21554 = ~n21420 & ~n21500;
  assign n21555 = ~n21420 & n21485;
  assign n21556 = ~n21553 & ~n21554;
  assign n21557 = ~n21555 & n21556;
  assign n21558 = n21483 & n21547;
  assign n21559 = ~n21483 & ~n21547;
  assign n21560 = ~n21558 & ~n21559;
  assign n21561 = n21557 & ~n21560;
  assign n21562 = ~n21557 & n21560;
  assign n21563 = ~n21561 & ~n21562;
  assign n21564 = n19604 & ~n21563;
  assign n21565 = ~n21551 & ~n21552;
  assign n21566 = ~n21564 & n21565;
  assign n21567 = n19675 & ~n21420;
  assign n21568 = ~P4_B_REG & n19560;
  assign n21569 = ~n19561 & ~n21568;
  assign n21570 = P4_REG1_REG_30_ & n19585;
  assign n21571 = P4_REG2_REG_30_ & n19587;
  assign n21572 = P4_REG0_REG_30_ & n19583;
  assign n21573 = ~n21570 & ~n21571;
  assign n21574 = ~n21572 & n21573;
  assign n21575 = ~n21569 & ~n21574;
  assign n21576 = n19573 & n21575;
  assign n21577 = n21420 & n21560;
  assign n21578 = n21485 & n21577;
  assign n21579 = ~n21420 & ~n21560;
  assign n21580 = ~n21485 & n21579;
  assign n21581 = ~n21578 & ~n21580;
  assign n21582 = ~n21501 & ~n21560;
  assign n21583 = ~n21517 & n21582;
  assign n21584 = ~n21502 & n21560;
  assign n21585 = n21517 & n21584;
  assign n21586 = n21581 & ~n21583;
  assign n21587 = ~n21585 & n21586;
  assign n21588 = n19627 & ~n21587;
  assign n21589 = n19622 & ~n21563;
  assign n21590 = n19625 & ~n21587;
  assign n21591 = ~n21589 & ~n21590;
  assign n21592 = n21485 & ~n21529;
  assign n21593 = ~n21420 & ~n21529;
  assign n21594 = ~n21592 & ~n21593;
  assign n21595 = ~n21555 & n21594;
  assign n21596 = ~n21560 & n21595;
  assign n21597 = n21560 & ~n21595;
  assign n21598 = ~n21596 & ~n21597;
  assign n21599 = n19617 & ~n21598;
  assign n21600 = n19611 & ~n21598;
  assign n21601 = n19614 & ~n21587;
  assign n21602 = n19619 & ~n21587;
  assign n21603 = ~n21601 & ~n21602;
  assign n21604 = ~n21599 & ~n21600;
  assign n21605 = n21603 & n21604;
  assign n21606 = ~n21567 & ~n21576;
  assign n21607 = ~n21588 & n21606;
  assign n21608 = n21591 & n21607;
  assign n21609 = n21605 & n21608;
  assign n21610 = n21566 & n21609;
  assign n21611 = n19554 & ~n21610;
  assign n21612 = P4_REG0_REG_29_ & ~n19554;
  assign n2491 = n21611 | n21612;
  assign n21614 = P2_P3_DATAO_REG_30_ & ~n19561;
  assign n21615 = n19568 & n21614;
  assign n21616 = P4_REG1_REG_31_ & n19585;
  assign n21617 = P4_REG2_REG_31_ & n19587;
  assign n21618 = P4_REG0_REG_31_ & n19583;
  assign n21619 = ~n21616 & ~n21617;
  assign n21620 = ~n21618 & n21619;
  assign n21621 = ~n21569 & ~n21620;
  assign n21622 = n19573 & n21621;
  assign n21623 = n21548 & ~n21614;
  assign n21624 = ~n21548 & n21614;
  assign n21625 = ~n21623 & ~n21624;
  assign n21626 = n19571 & n21625;
  assign n21627 = ~n21615 & ~n21622;
  assign n21628 = ~n21626 & n21627;
  assign n21629 = n19554 & ~n21628;
  assign n21630 = P4_REG0_REG_30_ & ~n19554;
  assign n2496 = n21629 | n21630;
  assign n21632 = P2_P3_DATAO_REG_31_ & ~n19561;
  assign n21633 = n19568 & n21632;
  assign n21634 = n21623 & ~n21632;
  assign n21635 = ~n21623 & n21632;
  assign n21636 = ~n21634 & ~n21635;
  assign n21637 = n19571 & n21636;
  assign n21638 = ~n21622 & ~n21633;
  assign n21639 = ~n21637 & n21638;
  assign n21640 = n19554 & ~n21639;
  assign n21641 = P4_REG0_REG_31_ & ~n19554;
  assign n2501 = n21640 | n21641;
  assign n21643 = n19420 & ~n19469;
  assign n21644 = n19553 & n21643;
  assign n21645 = ~n19634 & n21644;
  assign n21646 = P4_REG1_REG_0_ & ~n21644;
  assign n2506 = n21645 | n21646;
  assign n21648 = ~n19690 & n21644;
  assign n21649 = P4_REG1_REG_1_ & ~n21644;
  assign n2511 = n21648 | n21649;
  assign n21651 = ~n19750 & n21644;
  assign n21652 = P4_REG1_REG_2_ & ~n21644;
  assign n2516 = n21651 | n21652;
  assign n21654 = ~n19815 & n21644;
  assign n21655 = P4_REG1_REG_3_ & ~n21644;
  assign n2521 = n21654 | n21655;
  assign n21657 = ~n19886 & n21644;
  assign n21658 = P4_REG1_REG_4_ & ~n21644;
  assign n2526 = n21657 | n21658;
  assign n21660 = ~n19951 & n21644;
  assign n21661 = P4_REG1_REG_5_ & ~n21644;
  assign n2531 = n21660 | n21661;
  assign n21663 = ~n20025 & n21644;
  assign n21664 = P4_REG1_REG_6_ & ~n21644;
  assign n2536 = n21663 | n21664;
  assign n21666 = ~n20095 & n21644;
  assign n21667 = P4_REG1_REG_7_ & ~n21644;
  assign n2541 = n21666 | n21667;
  assign n21669 = ~n20163 & n21644;
  assign n21670 = P4_REG1_REG_8_ & ~n21644;
  assign n2546 = n21669 | n21670;
  assign n21672 = ~n20233 & n21644;
  assign n21673 = P4_REG1_REG_9_ & ~n21644;
  assign n2551 = n21672 | n21673;
  assign n21675 = ~n20297 & n21644;
  assign n21676 = P4_REG1_REG_10_ & ~n21644;
  assign n2556 = n21675 | n21676;
  assign n21678 = ~n20376 & n21644;
  assign n21679 = P4_REG1_REG_11_ & ~n21644;
  assign n2561 = n21678 | n21679;
  assign n21681 = ~n20448 & n21644;
  assign n21682 = P4_REG1_REG_12_ & ~n21644;
  assign n2566 = n21681 | n21682;
  assign n21684 = ~n20519 & n21644;
  assign n21685 = P4_REG1_REG_13_ & ~n21644;
  assign n2571 = n21684 | n21685;
  assign n21687 = ~n20588 & n21644;
  assign n21688 = P4_REG1_REG_14_ & ~n21644;
  assign n2576 = n21687 | n21688;
  assign n21690 = ~n20656 & n21644;
  assign n21691 = P4_REG1_REG_15_ & ~n21644;
  assign n2581 = n21690 | n21691;
  assign n21693 = ~n20728 & n21644;
  assign n21694 = P4_REG1_REG_16_ & ~n21644;
  assign n2586 = n21693 | n21694;
  assign n21696 = ~n20804 & n21644;
  assign n21697 = P4_REG1_REG_17_ & ~n21644;
  assign n2591 = n21696 | n21697;
  assign n21699 = ~n20875 & n21644;
  assign n21700 = P4_REG1_REG_18_ & ~n21644;
  assign n2596 = n21699 | n21700;
  assign n21702 = ~n20943 & n21644;
  assign n21703 = P4_REG1_REG_19_ & ~n21644;
  assign n2601 = n21702 | n21703;
  assign n21705 = ~n21007 & n21644;
  assign n21706 = P4_REG1_REG_20_ & ~n21644;
  assign n2606 = n21705 | n21706;
  assign n21708 = ~n21073 & n21644;
  assign n21709 = P4_REG1_REG_21_ & ~n21644;
  assign n2611 = n21708 | n21709;
  assign n21711 = ~n21140 & n21644;
  assign n21712 = P4_REG1_REG_22_ & ~n21644;
  assign n2616 = n21711 | n21712;
  assign n21714 = ~n21206 & n21644;
  assign n21715 = P4_REG1_REG_23_ & ~n21644;
  assign n2621 = n21714 | n21715;
  assign n21717 = ~n21275 & n21644;
  assign n21718 = P4_REG1_REG_24_ & ~n21644;
  assign n2626 = n21717 | n21718;
  assign n21720 = ~n21339 & n21644;
  assign n21721 = P4_REG1_REG_25_ & ~n21644;
  assign n2631 = n21720 | n21721;
  assign n21723 = ~n21406 & n21644;
  assign n21724 = P4_REG1_REG_26_ & ~n21644;
  assign n2636 = n21723 | n21724;
  assign n21726 = ~n21471 & n21644;
  assign n21727 = P4_REG1_REG_27_ & ~n21644;
  assign n2641 = n21726 | n21727;
  assign n21729 = ~n21543 & n21644;
  assign n21730 = P4_REG1_REG_28_ & ~n21644;
  assign n2646 = n21729 | n21730;
  assign n21732 = ~n21610 & n21644;
  assign n21733 = P4_REG1_REG_29_ & ~n21644;
  assign n2651 = n21732 | n21733;
  assign n21735 = ~n21628 & n21644;
  assign n21736 = P4_REG1_REG_30_ & ~n21644;
  assign n2656 = n21735 | n21736;
  assign n21738 = ~n21639 & n21644;
  assign n21739 = P4_REG1_REG_31_ & ~n21644;
  assign n2661 = n21738 | n21739;
  assign n21741 = n19479 & n19571;
  assign n21742 = n19476 & n19483;
  assign n21743 = n19603 & n21742;
  assign n21744 = ~n19480 & n19573;
  assign n21745 = n19469 & ~n21744;
  assign n21746 = ~n19473 & n21745;
  assign n21747 = n19552 & n21746;
  assign n21748 = ~n21743 & ~n21747;
  assign n21749 = n19420 & ~n21748;
  assign n21750 = n21741 & n21749;
  assign n21751 = ~n19567 & n21750;
  assign n21752 = n19568 & n21749;
  assign n21753 = ~n19567 & n21752;
  assign n21754 = ~n19633 & n21749;
  assign n21755 = P4_REG2_REG_0_ & ~n21749;
  assign n21756 = ~n21754 & ~n21755;
  assign n21757 = ~n21751 & ~n21753;
  assign n21758 = n21756 & n21757;
  assign n21759 = n21743 & n21749;
  assign n21760 = P4_REG3_REG_0_ & n21759;
  assign n21761 = n19574 & n21749;
  assign n21762 = ~n19591 & n21761;
  assign n21763 = ~n19479 & ~n19483;
  assign n21764 = n19476 & n21763;
  assign n21765 = n21749 & n21764;
  assign n21766 = ~n19602 & n21765;
  assign n21767 = ~n21760 & ~n21762;
  assign n21768 = ~n21766 & n21767;
  assign n2666 = ~n21758 | ~n21768;
  assign n21770 = ~n19663 & n21750;
  assign n21771 = ~n19643 & n21752;
  assign n21772 = ~n19689 & n21749;
  assign n21773 = P4_REG2_REG_1_ & ~n21749;
  assign n21774 = ~n21772 & ~n21773;
  assign n21775 = ~n21770 & ~n21771;
  assign n21776 = n21774 & n21775;
  assign n21777 = P4_REG3_REG_1_ & n21759;
  assign n21778 = ~n19659 & n21761;
  assign n21779 = ~n19651 & n21765;
  assign n21780 = ~n21777 & ~n21778;
  assign n21781 = ~n21779 & n21780;
  assign n2671 = ~n21776 | ~n21781;
  assign n21783 = n19725 & n21750;
  assign n21784 = ~n19699 & n21752;
  assign n21785 = ~n19749 & n21749;
  assign n21786 = P4_REG2_REG_2_ & ~n21749;
  assign n21787 = ~n21785 & ~n21786;
  assign n21788 = ~n21783 & ~n21784;
  assign n21789 = n21787 & n21788;
  assign n21790 = P4_REG3_REG_2_ & n21759;
  assign n21791 = ~n19720 & n21761;
  assign n21792 = n19712 & n21765;
  assign n21793 = ~n21790 & ~n21791;
  assign n21794 = ~n21792 & n21793;
  assign n2676 = ~n21789 | ~n21794;
  assign n21796 = n19773 & n21750;
  assign n21797 = ~n19770 & n21752;
  assign n21798 = ~n19814 & n21749;
  assign n21799 = P4_REG2_REG_3_ & ~n21749;
  assign n21800 = ~n21798 & ~n21799;
  assign n21801 = ~n21796 & ~n21797;
  assign n21802 = n21800 & n21801;
  assign n21803 = ~P4_REG3_REG_3_ & n21759;
  assign n21804 = ~n19763 & n21761;
  assign n21805 = ~n19788 & n21765;
  assign n21806 = ~n21803 & ~n21804;
  assign n21807 = ~n21805 & n21806;
  assign n2681 = ~n21802 | ~n21807;
  assign n21809 = n19856 & n21750;
  assign n21810 = ~n19824 & n21752;
  assign n21811 = ~n19885 & n21749;
  assign n21812 = P4_REG2_REG_4_ & ~n21749;
  assign n21813 = ~n21811 & ~n21812;
  assign n21814 = ~n21809 & ~n21810;
  assign n21815 = n21813 & n21814;
  assign n21816 = ~n19756 & n21759;
  assign n21817 = ~n19851 & n21761;
  assign n21818 = ~n19839 & n21765;
  assign n21819 = ~n21816 & ~n21817;
  assign n21820 = ~n21818 & n21819;
  assign n2686 = ~n21815 | ~n21820;
  assign n21822 = n19911 & n21750;
  assign n21823 = ~n19908 & n21752;
  assign n21824 = ~n19950 & n21749;
  assign n21825 = P4_REG2_REG_5_ & ~n21749;
  assign n21826 = ~n21824 & ~n21825;
  assign n21827 = ~n21822 & ~n21823;
  assign n21828 = n21826 & n21827;
  assign n21829 = ~n19844 & n21759;
  assign n21830 = ~n19901 & n21761;
  assign n21831 = n19926 & n21765;
  assign n21832 = ~n21829 & ~n21830;
  assign n21833 = ~n21831 & n21832;
  assign n2691 = ~n21828 | ~n21833;
  assign n21835 = n19976 & n21750;
  assign n21836 = ~n19972 & n21752;
  assign n21837 = ~n20024 & n21749;
  assign n21838 = P4_REG2_REG_6_ & ~n21749;
  assign n21839 = ~n21837 & ~n21838;
  assign n21840 = ~n21835 & ~n21836;
  assign n21841 = n21839 & n21840;
  assign n21842 = ~n19894 & n21759;
  assign n21843 = ~n19965 & n21761;
  assign n21844 = ~n19997 & n21765;
  assign n21845 = ~n21842 & ~n21843;
  assign n21846 = ~n21844 & n21845;
  assign n2696 = ~n21841 | ~n21846;
  assign n21848 = n20050 & n21750;
  assign n21849 = ~n20047 & n21752;
  assign n21850 = ~n20094 & n21749;
  assign n21851 = P4_REG2_REG_7_ & ~n21749;
  assign n21852 = ~n21850 & ~n21851;
  assign n21853 = ~n21848 & ~n21849;
  assign n21854 = n21852 & n21853;
  assign n21855 = ~n19958 & n21759;
  assign n21856 = ~n20040 & n21761;
  assign n21857 = n20065 & n21765;
  assign n21858 = ~n21855 & ~n21856;
  assign n21859 = ~n21857 & n21858;
  assign n2701 = ~n21854 | ~n21859;
  assign n21861 = n20119 & n21750;
  assign n21862 = ~n20116 & n21752;
  assign n21863 = ~n20162 & n21749;
  assign n21864 = P4_REG2_REG_8_ & ~n21749;
  assign n21865 = ~n21863 & ~n21864;
  assign n21866 = ~n21861 & ~n21862;
  assign n21867 = n21865 & n21866;
  assign n21868 = ~n20033 & n21759;
  assign n21869 = ~n20109 & n21761;
  assign n21870 = ~n20136 & n21765;
  assign n21871 = ~n21868 & ~n21869;
  assign n21872 = ~n21870 & n21871;
  assign n2706 = ~n21867 | ~n21872;
  assign n21874 = n20190 & n21750;
  assign n21875 = ~n20187 & n21752;
  assign n21876 = ~n20232 & n21749;
  assign n21877 = P4_REG2_REG_9_ & ~n21749;
  assign n21878 = ~n21876 & ~n21877;
  assign n21879 = ~n21874 & ~n21875;
  assign n21880 = n21878 & n21879;
  assign n21881 = ~n20102 & n21759;
  assign n21882 = ~n20178 & n21761;
  assign n21883 = ~n20203 & n21765;
  assign n21884 = ~n21881 & ~n21882;
  assign n21885 = ~n21883 & n21884;
  assign n2711 = ~n21880 | ~n21885;
  assign n21887 = n20257 & n21750;
  assign n21888 = ~n20254 & n21752;
  assign n21889 = ~n20296 & n21749;
  assign n21890 = P4_REG2_REG_10_ & ~n21749;
  assign n21891 = ~n21889 & ~n21890;
  assign n21892 = ~n21887 & ~n21888;
  assign n21893 = n21891 & n21892;
  assign n21894 = ~n20171 & n21759;
  assign n21895 = ~n20247 & n21761;
  assign n21896 = n20272 & n21765;
  assign n21897 = ~n21894 & ~n21895;
  assign n21898 = ~n21896 & n21897;
  assign n2716 = ~n21893 | ~n21898;
  assign n21900 = n20323 & n21750;
  assign n21901 = ~n20320 & n21752;
  assign n21902 = ~n20375 & n21749;
  assign n21903 = P4_REG2_REG_11_ & ~n21749;
  assign n21904 = ~n21902 & ~n21903;
  assign n21905 = ~n21900 & ~n21901;
  assign n21906 = n21904 & n21905;
  assign n21907 = ~n20240 & n21759;
  assign n21908 = ~n20311 & n21761;
  assign n21909 = ~n20341 & n21765;
  assign n21910 = ~n21907 & ~n21908;
  assign n21911 = ~n21909 & n21910;
  assign n2721 = ~n21906 | ~n21911;
  assign n21913 = n20400 & n21750;
  assign n21914 = ~n20397 & n21752;
  assign n21915 = ~n20447 & n21749;
  assign n21916 = P4_REG2_REG_12_ & ~n21749;
  assign n21917 = ~n21915 & ~n21916;
  assign n21918 = ~n21913 & ~n21914;
  assign n21919 = n21917 & n21918;
  assign n21920 = ~n20304 & n21759;
  assign n21921 = ~n20390 & n21761;
  assign n21922 = ~n20413 & n21765;
  assign n21923 = ~n21920 & ~n21921;
  assign n21924 = ~n21922 & n21923;
  assign n2726 = ~n21919 | ~n21924;
  assign n21926 = n20474 & n21750;
  assign n21927 = ~n20471 & n21752;
  assign n21928 = ~n20518 & n21749;
  assign n21929 = P4_REG2_REG_13_ & ~n21749;
  assign n21930 = ~n21928 & ~n21929;
  assign n21931 = ~n21926 & ~n21927;
  assign n21932 = n21930 & n21931;
  assign n21933 = ~n20386 & n21759;
  assign n21934 = ~n20462 & n21761;
  assign n21935 = n20489 & n21765;
  assign n21936 = ~n21933 & ~n21934;
  assign n21937 = ~n21935 & n21936;
  assign n2731 = ~n21932 | ~n21937;
  assign n21939 = n20543 & n21750;
  assign n21940 = ~n20540 & n21752;
  assign n21941 = ~n21939 & ~n21940;
  assign n21942 = ~n20458 & n21759;
  assign n21943 = ~n20533 & n21761;
  assign n21944 = ~n20558 & n21765;
  assign n21945 = ~n21942 & ~n21943;
  assign n21946 = ~n21944 & n21945;
  assign n21947 = ~n20587 & n21749;
  assign n21948 = P4_REG2_REG_14_ & ~n21749;
  assign n21949 = ~n21947 & ~n21948;
  assign n21950 = n21941 & n21946;
  assign n2736 = ~n21949 | ~n21950;
  assign n21952 = n20614 & n21750;
  assign n21953 = ~n20611 & n21752;
  assign n21954 = ~n21952 & ~n21953;
  assign n21955 = ~n20529 & n21759;
  assign n21956 = ~n20602 & n21761;
  assign n21957 = ~n20626 & n21765;
  assign n21958 = ~n21955 & ~n21956;
  assign n21959 = ~n21957 & n21958;
  assign n21960 = ~n20655 & n21749;
  assign n21961 = P4_REG2_REG_15_ & ~n21749;
  assign n21962 = ~n21960 & ~n21961;
  assign n21963 = n21954 & n21959;
  assign n2741 = ~n21962 | ~n21963;
  assign n21965 = n20680 & n21750;
  assign n21966 = ~n20677 & n21752;
  assign n21967 = ~n21965 & ~n21966;
  assign n21968 = ~n20598 & n21759;
  assign n21969 = ~n20670 & n21761;
  assign n21970 = ~n20695 & n21765;
  assign n21971 = ~n21968 & ~n21969;
  assign n21972 = ~n21970 & n21971;
  assign n21973 = ~n20727 & n21749;
  assign n21974 = P4_REG2_REG_16_ & ~n21749;
  assign n21975 = ~n21973 & ~n21974;
  assign n21976 = n21967 & n21972;
  assign n2746 = ~n21975 | ~n21976;
  assign n21978 = n20754 & n21750;
  assign n21979 = ~n20751 & n21752;
  assign n21980 = ~n21978 & ~n21979;
  assign n21981 = ~n20666 & n21759;
  assign n21982 = ~n20742 & n21761;
  assign n21983 = n20769 & n21765;
  assign n21984 = ~n21981 & ~n21982;
  assign n21985 = ~n21983 & n21984;
  assign n21986 = ~n20803 & n21749;
  assign n21987 = P4_REG2_REG_17_ & ~n21749;
  assign n21988 = ~n21986 & ~n21987;
  assign n21989 = n21980 & n21985;
  assign n2751 = ~n21988 | ~n21989;
  assign n21991 = n20828 & n21750;
  assign n21992 = ~n20825 & n21752;
  assign n21993 = ~n21991 & ~n21992;
  assign n21994 = ~n20738 & n21759;
  assign n21995 = ~n20818 & n21761;
  assign n21996 = ~n20845 & n21765;
  assign n21997 = ~n21994 & ~n21995;
  assign n21998 = ~n21996 & n21997;
  assign n21999 = ~n20874 & n21749;
  assign n22000 = P4_REG2_REG_18_ & ~n21749;
  assign n22001 = ~n21999 & ~n22000;
  assign n22002 = n21993 & n21998;
  assign n2756 = ~n22001 | ~n22002;
  assign n22004 = ~n20814 & n21759;
  assign n22005 = ~n20889 & n21761;
  assign n22006 = ~n22004 & ~n22005;
  assign n22007 = n20898 & n21750;
  assign n22008 = ~n20895 & n21752;
  assign n22009 = ~n22007 & ~n22008;
  assign n22010 = ~n20911 & n21765;
  assign n22011 = ~n20942 & n21749;
  assign n22012 = P4_REG2_REG_19_ & ~n21749;
  assign n22013 = ~n22011 & ~n22012;
  assign n22014 = n22006 & n22009;
  assign n22015 = ~n22010 & n22014;
  assign n2761 = ~n22013 | ~n22015;
  assign n22017 = ~n20885 & n21759;
  assign n22018 = ~n20957 & n21761;
  assign n22019 = ~n22017 & ~n22018;
  assign n22020 = n20962 & n21750;
  assign n22021 = n20959 & n21752;
  assign n22022 = ~n22020 & ~n22021;
  assign n22023 = n20977 & n21765;
  assign n22024 = ~n21006 & n21749;
  assign n22025 = P4_REG2_REG_20_ & ~n21749;
  assign n22026 = ~n22024 & ~n22025;
  assign n22027 = n22019 & n22022;
  assign n22028 = ~n22023 & n22027;
  assign n2766 = ~n22026 | ~n22028;
  assign n22030 = ~n20953 & n21759;
  assign n22031 = ~n21021 & n21761;
  assign n22032 = ~n22030 & ~n22031;
  assign n22033 = n21028 & n21750;
  assign n22034 = n21025 & n21752;
  assign n22035 = ~n22033 & ~n22034;
  assign n22036 = n21043 & n21765;
  assign n22037 = ~n21072 & n21749;
  assign n22038 = P4_REG2_REG_21_ & ~n21749;
  assign n22039 = ~n22037 & ~n22038;
  assign n22040 = n22032 & n22035;
  assign n22041 = ~n22036 & n22040;
  assign n2771 = ~n22039 | ~n22041;
  assign n22043 = ~n21017 & n21759;
  assign n22044 = ~n21087 & n21761;
  assign n22045 = ~n22043 & ~n22044;
  assign n22046 = n21092 & n21750;
  assign n22047 = n21089 & n21752;
  assign n22048 = ~n22046 & ~n22047;
  assign n22049 = ~n21110 & n21765;
  assign n22050 = ~n21139 & n21749;
  assign n22051 = P4_REG2_REG_22_ & ~n21749;
  assign n22052 = ~n22050 & ~n22051;
  assign n22053 = n22045 & n22048;
  assign n22054 = ~n22049 & n22053;
  assign n2776 = ~n22052 | ~n22054;
  assign n22056 = ~n21083 & n21759;
  assign n22057 = ~n21154 & n21761;
  assign n22058 = ~n22056 & ~n22057;
  assign n22059 = n21161 & n21750;
  assign n22060 = n21158 & n21752;
  assign n22061 = ~n22059 & ~n22060;
  assign n22062 = ~n21173 & n21765;
  assign n22063 = ~n21205 & n21749;
  assign n22064 = P4_REG2_REG_23_ & ~n21749;
  assign n22065 = ~n22063 & ~n22064;
  assign n22066 = n22058 & n22061;
  assign n22067 = ~n22062 & n22066;
  assign n2781 = ~n22065 | ~n22067;
  assign n22069 = ~n21150 & n21759;
  assign n22070 = ~n21220 & n21761;
  assign n22071 = ~n22069 & ~n22070;
  assign n22072 = n21225 & n21750;
  assign n22073 = n21222 & n21752;
  assign n22074 = ~n22072 & ~n22073;
  assign n22075 = ~n21240 & n21765;
  assign n22076 = ~n21274 & n21749;
  assign n22077 = P4_REG2_REG_24_ & ~n21749;
  assign n22078 = ~n22076 & ~n22077;
  assign n22079 = n22071 & n22074;
  assign n22080 = ~n22075 & n22079;
  assign n2786 = ~n22078 | ~n22080;
  assign n22082 = ~n21216 & n21759;
  assign n22083 = ~n21289 & n21761;
  assign n22084 = ~n22082 & ~n22083;
  assign n22085 = n21296 & n21750;
  assign n22086 = n21293 & n21752;
  assign n22087 = ~n22085 & ~n22086;
  assign n22088 = ~n21309 & n21765;
  assign n22089 = ~n21338 & n21749;
  assign n22090 = P4_REG2_REG_25_ & ~n21749;
  assign n22091 = ~n22089 & ~n22090;
  assign n22092 = n22084 & n22087;
  assign n22093 = ~n22088 & n22092;
  assign n2791 = ~n22091 | ~n22093;
  assign n22095 = ~n21285 & n21759;
  assign n22096 = ~n21353 & n21761;
  assign n22097 = ~n22095 & ~n22096;
  assign n22098 = n21358 & n21750;
  assign n22099 = n21355 & n21752;
  assign n22100 = ~n22098 & ~n22099;
  assign n22101 = n21374 & n21765;
  assign n22102 = ~n21405 & n21749;
  assign n22103 = P4_REG2_REG_26_ & ~n21749;
  assign n22104 = ~n22102 & ~n22103;
  assign n22105 = n22097 & n22100;
  assign n22106 = ~n22101 & n22105;
  assign n2796 = ~n22104 | ~n22106;
  assign n22108 = ~n21349 & n21759;
  assign n22109 = ~n21420 & n21761;
  assign n22110 = ~n22108 & ~n22109;
  assign n22111 = n21425 & n21750;
  assign n22112 = n21422 & n21752;
  assign n22113 = ~n22111 & ~n22112;
  assign n22114 = ~n21438 & n21765;
  assign n22115 = ~n21470 & n21749;
  assign n22116 = P4_REG2_REG_27_ & ~n21749;
  assign n22117 = ~n22115 & ~n22116;
  assign n22118 = n22110 & n22113;
  assign n22119 = ~n22114 & n22118;
  assign n2801 = ~n22117 | ~n22119;
  assign n22121 = ~n21416 & n21759;
  assign n22122 = ~n21483 & n21761;
  assign n22123 = ~n22121 & ~n22122;
  assign n22124 = n21488 & n21750;
  assign n22125 = n21485 & n21752;
  assign n22126 = ~n22124 & ~n22125;
  assign n22127 = ~n21506 & n21765;
  assign n22128 = ~n21542 & n21749;
  assign n22129 = P4_REG2_REG_28_ & ~n21749;
  assign n22130 = ~n22128 & ~n22129;
  assign n22131 = n22123 & n22126;
  assign n22132 = ~n22127 & n22131;
  assign n2806 = ~n22130 | ~n22132;
  assign n22134 = n21547 & n21752;
  assign n22135 = n21479 & n21759;
  assign n22136 = n21550 & n21750;
  assign n22137 = ~n21563 & n21765;
  assign n22138 = ~n21609 & n21749;
  assign n22139 = P4_REG2_REG_29_ & ~n21749;
  assign n22140 = ~n22138 & ~n22139;
  assign n22141 = ~n22134 & ~n22135;
  assign n22142 = ~n22136 & n22141;
  assign n22143 = ~n22137 & n22142;
  assign n2811 = ~n22140 | ~n22143;
  assign n22145 = n21625 & n21750;
  assign n22146 = n21614 & n21752;
  assign n22147 = n21622 & n21749;
  assign n22148 = P4_REG2_REG_30_ & ~n21749;
  assign n22149 = ~n22147 & ~n22148;
  assign n22150 = ~n22145 & ~n22146;
  assign n2816 = ~n22149 | ~n22150;
  assign n22152 = n21636 & n21750;
  assign n22153 = n21632 & n21752;
  assign n22154 = P4_REG2_REG_31_ & ~n21749;
  assign n22155 = ~n22147 & ~n22154;
  assign n22156 = ~n22152 & ~n22153;
  assign n2821 = ~n22155 | ~n22156;
  assign n22158 = n19407 & n19418;
  assign n22159 = n19419 & ~n19573;
  assign n22160 = n19407 & ~n22159;
  assign n22161 = ~n19561 & ~n22160;
  assign n3241 = ~P4_STATE_REG | n22161;
  assign n22163 = ~n22158 & ~n3241;
  assign n22164 = P4_ADDR_REG_19_ & n22163;
  assign n22165 = P4_STATE_REG & ~n19407;
  assign n22166 = ~n22163 & n22165;
  assign n22167 = n19557 & n22166;
  assign n22168 = ~P4_REG1_REG_18_ & n20822;
  assign n22169 = P4_REG1_REG_19_ & n19479;
  assign n22170 = ~P4_REG1_REG_19_ & ~n19479;
  assign n22171 = ~n22169 & ~n22170;
  assign n22172 = ~n22168 & ~n22171;
  assign n22173 = P4_REG1_REG_17_ & ~n20748;
  assign n22174 = ~P4_REG1_REG_17_ & n20748;
  assign n22175 = P4_REG1_REG_16_ & ~n20674;
  assign n22176 = ~P4_REG1_REG_16_ & n20674;
  assign n22177 = P4_REG1_REG_12_ & ~n20394;
  assign n22178 = ~P4_REG1_REG_12_ & n20394;
  assign n22179 = P4_REG1_REG_11_ & ~n20317;
  assign n22180 = ~P4_REG1_REG_11_ & n20317;
  assign n22181 = P4_REG1_REG_9_ & ~n20184;
  assign n22182 = ~P4_REG1_REG_9_ & n20184;
  assign n22183 = P4_REG1_REG_7_ & ~n20044;
  assign n22184 = ~P4_REG1_REG_7_ & n20044;
  assign n22185 = P4_REG1_REG_6_ & ~n19969;
  assign n22186 = ~P4_REG1_REG_6_ & n19969;
  assign n22187 = P4_REG1_REG_4_ & ~n19821;
  assign n22188 = ~P4_REG1_REG_4_ & n19821;
  assign n22189 = P4_REG1_REG_2_ & ~n19696;
  assign n22190 = ~P4_REG1_REG_2_ & n19696;
  assign n22191 = P4_REG1_REG_0_ & ~n19564;
  assign n22192 = P4_REG1_REG_1_ & n22191;
  assign n22193 = ~P4_REG1_REG_1_ & ~n22191;
  assign n22194 = ~n19640 & ~n22193;
  assign n22195 = ~n22192 & ~n22194;
  assign n22196 = ~n22190 & ~n22195;
  assign n22197 = ~n22189 & ~n22196;
  assign n22198 = P4_REG1_REG_3_ & ~n22197;
  assign n22199 = ~n19767 & ~n22197;
  assign n22200 = P4_REG1_REG_3_ & ~n19767;
  assign n22201 = ~n22198 & ~n22199;
  assign n22202 = ~n22200 & n22201;
  assign n22203 = ~n22188 & ~n22202;
  assign n22204 = ~n22187 & ~n22203;
  assign n22205 = P4_REG1_REG_5_ & ~n22204;
  assign n22206 = ~P4_REG1_REG_5_ & n22204;
  assign n22207 = ~n19905 & ~n22206;
  assign n22208 = ~n22205 & ~n22207;
  assign n22209 = ~n22186 & ~n22208;
  assign n22210 = ~n22185 & ~n22209;
  assign n22211 = ~n22184 & ~n22210;
  assign n22212 = ~n22183 & ~n22211;
  assign n22213 = P4_REG1_REG_8_ & ~n22212;
  assign n22214 = ~P4_REG1_REG_8_ & n22212;
  assign n22215 = ~n20113 & ~n22214;
  assign n22216 = ~n22213 & ~n22215;
  assign n22217 = ~n22182 & ~n22216;
  assign n22218 = ~n22181 & ~n22217;
  assign n22219 = P4_REG1_REG_10_ & ~n22218;
  assign n22220 = ~P4_REG1_REG_10_ & n22218;
  assign n22221 = ~n20251 & ~n22220;
  assign n22222 = ~n22219 & ~n22221;
  assign n22223 = ~n22180 & ~n22222;
  assign n22224 = ~n22179 & ~n22223;
  assign n22225 = ~n22178 & ~n22224;
  assign n22226 = ~n22177 & ~n22225;
  assign n22227 = P4_REG1_REG_13_ & ~n22226;
  assign n22228 = ~P4_REG1_REG_13_ & n22226;
  assign n22229 = ~n20468 & ~n22228;
  assign n22230 = ~n22227 & ~n22229;
  assign n22231 = P4_REG1_REG_14_ & ~n22230;
  assign n22232 = ~P4_REG1_REG_14_ & n22230;
  assign n22233 = ~n20537 & ~n22232;
  assign n22234 = ~n22231 & ~n22233;
  assign n22235 = P4_REG1_REG_15_ & ~n22234;
  assign n22236 = ~P4_REG1_REG_15_ & n22234;
  assign n22237 = ~n20608 & ~n22236;
  assign n22238 = ~n22235 & ~n22237;
  assign n22239 = ~n22176 & ~n22238;
  assign n22240 = ~n22175 & ~n22239;
  assign n22241 = ~n22174 & ~n22240;
  assign n22242 = ~n22173 & ~n22241;
  assign n22243 = P4_REG1_REG_18_ & ~n20822;
  assign n22244 = n22242 & ~n22243;
  assign n22245 = n22172 & ~n22244;
  assign n22246 = n22171 & ~n22243;
  assign n22247 = ~n22168 & ~n22242;
  assign n22248 = n22246 & ~n22247;
  assign n22249 = ~n22245 & ~n22248;
  assign n22250 = n22167 & n22249;
  assign n22251 = ~n22164 & ~n22250;
  assign n22252 = ~n19568 & ~n21743;
  assign n22253 = ~n19622 & ~n19625;
  assign n22254 = ~n21741 & n22253;
  assign n22255 = ~n19610 & ~n19627;
  assign n22256 = ~n19619 & n22255;
  assign n22257 = ~n19616 & ~n21764;
  assign n22258 = ~n19614 & n22257;
  assign n22259 = n22252 & n22254;
  assign n22260 = n22256 & n22259;
  assign n22261 = n22258 & n22260;
  assign n22262 = n19560 & ~n22261;
  assign n22263 = ~n19479 & n22262;
  assign n22264 = n19420 & ~n22163;
  assign n22265 = n22263 & n22264;
  assign n22266 = P4_REG3_REG_19_ & ~P4_STATE_REG;
  assign n22267 = ~n22265 & ~n22266;
  assign n22268 = n19560 & n22166;
  assign n22269 = ~n19479 & n22268;
  assign n22270 = n19557 & ~n22261;
  assign n22271 = n22264 & n22270;
  assign n22272 = n22249 & n22271;
  assign n22273 = n22267 & ~n22269;
  assign n22274 = ~n22272 & n22273;
  assign n22275 = ~P4_REG2_REG_18_ & n20822;
  assign n22276 = P4_REG2_REG_19_ & n19479;
  assign n22277 = ~P4_REG2_REG_19_ & ~n19479;
  assign n22278 = ~n22276 & ~n22277;
  assign n22279 = ~n22275 & ~n22278;
  assign n22280 = P4_REG2_REG_17_ & ~n20748;
  assign n22281 = ~P4_REG2_REG_17_ & n20748;
  assign n22282 = P4_REG2_REG_16_ & ~n20674;
  assign n22283 = ~P4_REG2_REG_16_ & n20674;
  assign n22284 = P4_REG2_REG_15_ & ~n20608;
  assign n22285 = ~P4_REG2_REG_15_ & n20608;
  assign n22286 = P4_REG2_REG_14_ & ~n20537;
  assign n22287 = ~P4_REG2_REG_14_ & n20537;
  assign n22288 = P4_REG2_REG_13_ & ~n20468;
  assign n22289 = ~P4_REG2_REG_13_ & n20468;
  assign n22290 = P4_REG2_REG_12_ & ~n20394;
  assign n22291 = ~P4_REG2_REG_12_ & n20394;
  assign n22292 = P4_REG2_REG_11_ & ~n20317;
  assign n22293 = ~P4_REG2_REG_11_ & n20317;
  assign n22294 = P4_REG2_REG_10_ & ~n20251;
  assign n22295 = ~P4_REG2_REG_10_ & n20251;
  assign n22296 = P4_REG2_REG_9_ & ~n20184;
  assign n22297 = ~P4_REG2_REG_9_ & n20184;
  assign n22298 = P4_REG2_REG_8_ & ~n20113;
  assign n22299 = ~P4_REG2_REG_8_ & n20113;
  assign n22300 = P4_REG2_REG_7_ & ~n20044;
  assign n22301 = ~P4_REG2_REG_7_ & n20044;
  assign n22302 = P4_REG2_REG_6_ & ~n19969;
  assign n22303 = ~P4_REG2_REG_6_ & n19969;
  assign n22304 = P4_REG2_REG_5_ & ~n19905;
  assign n22305 = ~P4_REG2_REG_5_ & n19905;
  assign n22306 = P4_REG2_REG_4_ & ~n19821;
  assign n22307 = ~P4_REG2_REG_4_ & n19821;
  assign n22308 = P4_REG2_REG_3_ & ~n19767;
  assign n22309 = ~P4_REG2_REG_3_ & n19767;
  assign n22310 = P4_REG2_REG_2_ & ~n19696;
  assign n22311 = ~P4_REG2_REG_2_ & n19696;
  assign n22312 = P4_REG2_REG_0_ & ~n19564;
  assign n22313 = ~n19640 & n22312;
  assign n22314 = n19640 & ~n22312;
  assign n22315 = P4_REG2_REG_1_ & ~n22314;
  assign n22316 = ~n22313 & ~n22315;
  assign n22317 = ~n22311 & ~n22316;
  assign n22318 = ~n22310 & ~n22317;
  assign n22319 = ~n22309 & ~n22318;
  assign n22320 = ~n22308 & ~n22319;
  assign n22321 = ~n22307 & ~n22320;
  assign n22322 = ~n22306 & ~n22321;
  assign n22323 = ~n22305 & ~n22322;
  assign n22324 = ~n22304 & ~n22323;
  assign n22325 = ~n22303 & ~n22324;
  assign n22326 = ~n22302 & ~n22325;
  assign n22327 = ~n22301 & ~n22326;
  assign n22328 = ~n22300 & ~n22327;
  assign n22329 = ~n22299 & ~n22328;
  assign n22330 = ~n22298 & ~n22329;
  assign n22331 = ~n22297 & ~n22330;
  assign n22332 = ~n22296 & ~n22331;
  assign n22333 = ~n22295 & ~n22332;
  assign n22334 = ~n22294 & ~n22333;
  assign n22335 = ~n22293 & ~n22334;
  assign n22336 = ~n22292 & ~n22335;
  assign n22337 = ~n22291 & ~n22336;
  assign n22338 = ~n22290 & ~n22337;
  assign n22339 = ~n22289 & ~n22338;
  assign n22340 = ~n22288 & ~n22339;
  assign n22341 = ~n22287 & ~n22340;
  assign n22342 = ~n22286 & ~n22341;
  assign n22343 = ~n22285 & ~n22342;
  assign n22344 = ~n22284 & ~n22343;
  assign n22345 = ~n22283 & ~n22344;
  assign n22346 = ~n22282 & ~n22345;
  assign n22347 = ~n22281 & ~n22346;
  assign n22348 = ~n22280 & ~n22347;
  assign n22349 = P4_REG2_REG_18_ & ~n20822;
  assign n22350 = n22348 & ~n22349;
  assign n22351 = n22279 & ~n22350;
  assign n22352 = n22278 & ~n22349;
  assign n22353 = ~n22275 & ~n22348;
  assign n22354 = n22352 & ~n22353;
  assign n22355 = ~n22351 & ~n22354;
  assign n22356 = ~n19557 & ~n19560;
  assign n22357 = n22166 & n22356;
  assign n22358 = ~n22261 & n22356;
  assign n22359 = n22264 & n22358;
  assign n22360 = ~n22357 & ~n22359;
  assign n22361 = n22355 & ~n22360;
  assign n22362 = n22251 & n22274;
  assign n2826 = n22361 | ~n22362;
  assign n22364 = ~n20822 & n22262;
  assign n22365 = P4_REG1_REG_18_ & n20822;
  assign n22366 = ~P4_REG1_REG_18_ & ~n20822;
  assign n22367 = ~n22365 & ~n22366;
  assign n22368 = n22242 & ~n22367;
  assign n22369 = ~n22242 & n22367;
  assign n22370 = ~n22368 & ~n22369;
  assign n22371 = n22270 & ~n22370;
  assign n22372 = P4_REG2_REG_18_ & n20822;
  assign n22373 = ~P4_REG2_REG_18_ & ~n20822;
  assign n22374 = ~n22372 & ~n22373;
  assign n22375 = n22348 & ~n22374;
  assign n22376 = ~n22348 & n22374;
  assign n22377 = ~n22375 & ~n22376;
  assign n22378 = n22358 & ~n22377;
  assign n22379 = ~n22364 & ~n22371;
  assign n22380 = ~n22378 & n22379;
  assign n22381 = n22264 & ~n22380;
  assign n22382 = P4_ADDR_REG_18_ & n22163;
  assign n22383 = ~n20822 & n22268;
  assign n22384 = n22167 & ~n22370;
  assign n22385 = P4_REG3_REG_18_ & ~P4_STATE_REG;
  assign n22386 = n22357 & ~n22377;
  assign n22387 = ~n22382 & ~n22383;
  assign n22388 = ~n22384 & n22387;
  assign n22389 = ~n22385 & n22388;
  assign n22390 = ~n22386 & n22389;
  assign n2831 = n22381 | ~n22390;
  assign n22392 = ~n20748 & n22262;
  assign n22393 = P4_REG1_REG_17_ & n20748;
  assign n22394 = ~P4_REG1_REG_17_ & ~n20748;
  assign n22395 = ~n22393 & ~n22394;
  assign n22396 = n22240 & ~n22395;
  assign n22397 = ~n22240 & n22395;
  assign n22398 = ~n22396 & ~n22397;
  assign n22399 = n22270 & ~n22398;
  assign n22400 = P4_REG2_REG_17_ & n20748;
  assign n22401 = ~P4_REG2_REG_17_ & ~n20748;
  assign n22402 = ~n22400 & ~n22401;
  assign n22403 = n22346 & ~n22402;
  assign n22404 = ~n22346 & n22402;
  assign n22405 = ~n22403 & ~n22404;
  assign n22406 = n22358 & ~n22405;
  assign n22407 = ~n22392 & ~n22399;
  assign n22408 = ~n22406 & n22407;
  assign n22409 = n22264 & ~n22408;
  assign n22410 = P4_ADDR_REG_17_ & n22163;
  assign n22411 = ~n20748 & n22268;
  assign n22412 = n22167 & ~n22398;
  assign n22413 = P4_REG3_REG_17_ & ~P4_STATE_REG;
  assign n22414 = n22357 & ~n22405;
  assign n22415 = ~n22410 & ~n22411;
  assign n22416 = ~n22412 & n22415;
  assign n22417 = ~n22413 & n22416;
  assign n22418 = ~n22414 & n22417;
  assign n2836 = n22409 | ~n22418;
  assign n22420 = ~n20674 & n22262;
  assign n22421 = P4_REG1_REG_16_ & n20674;
  assign n22422 = ~P4_REG1_REG_16_ & ~n20674;
  assign n22423 = ~n22421 & ~n22422;
  assign n22424 = n22238 & ~n22423;
  assign n22425 = ~n22238 & n22423;
  assign n22426 = ~n22424 & ~n22425;
  assign n22427 = n22270 & ~n22426;
  assign n22428 = P4_REG2_REG_16_ & n20674;
  assign n22429 = ~P4_REG2_REG_16_ & ~n20674;
  assign n22430 = ~n22428 & ~n22429;
  assign n22431 = n22344 & ~n22430;
  assign n22432 = ~n22344 & n22430;
  assign n22433 = ~n22431 & ~n22432;
  assign n22434 = n22358 & ~n22433;
  assign n22435 = ~n22420 & ~n22427;
  assign n22436 = ~n22434 & n22435;
  assign n22437 = n22264 & ~n22436;
  assign n22438 = P4_ADDR_REG_16_ & n22163;
  assign n22439 = ~n20674 & n22268;
  assign n22440 = n22167 & ~n22426;
  assign n22441 = P4_REG3_REG_16_ & ~P4_STATE_REG;
  assign n22442 = n22357 & ~n22433;
  assign n22443 = ~n22438 & ~n22439;
  assign n22444 = ~n22440 & n22443;
  assign n22445 = ~n22441 & n22444;
  assign n22446 = ~n22442 & n22445;
  assign n2841 = n22437 | ~n22446;
  assign n22448 = P4_ADDR_REG_15_ & n22163;
  assign n22449 = ~n20608 & n22268;
  assign n22450 = ~n22448 & ~n22449;
  assign n22451 = P4_REG2_REG_15_ & n20608;
  assign n22452 = ~P4_REG2_REG_15_ & ~n20608;
  assign n22453 = ~n22451 & ~n22452;
  assign n22454 = n22342 & ~n22453;
  assign n22455 = ~n22342 & n22453;
  assign n22456 = ~n22454 & ~n22455;
  assign n22457 = n22357 & ~n22456;
  assign n22458 = P4_REG3_REG_15_ & ~P4_STATE_REG;
  assign n22459 = ~n22457 & ~n22458;
  assign n22460 = ~n22235 & ~n22236;
  assign n22461 = ~n20608 & ~n22460;
  assign n22462 = n20608 & n22460;
  assign n22463 = ~n22461 & ~n22462;
  assign n22464 = n22167 & ~n22463;
  assign n22465 = ~n20608 & n22262;
  assign n22466 = n22358 & ~n22456;
  assign n22467 = n22270 & ~n22463;
  assign n22468 = ~n22465 & ~n22466;
  assign n22469 = ~n22467 & n22468;
  assign n22470 = n22264 & ~n22469;
  assign n22471 = n22450 & n22459;
  assign n22472 = ~n22464 & n22471;
  assign n2846 = n22470 | ~n22472;
  assign n22474 = P4_ADDR_REG_14_ & n22163;
  assign n22475 = ~n20537 & n22268;
  assign n22476 = ~n22474 & ~n22475;
  assign n22477 = P4_REG2_REG_14_ & n20537;
  assign n22478 = ~P4_REG2_REG_14_ & ~n20537;
  assign n22479 = ~n22477 & ~n22478;
  assign n22480 = n22340 & ~n22479;
  assign n22481 = ~n22340 & n22479;
  assign n22482 = ~n22480 & ~n22481;
  assign n22483 = n22357 & ~n22482;
  assign n22484 = P4_REG3_REG_14_ & ~P4_STATE_REG;
  assign n22485 = ~n22483 & ~n22484;
  assign n22486 = ~n22231 & ~n22232;
  assign n22487 = ~n20537 & ~n22486;
  assign n22488 = n20537 & n22486;
  assign n22489 = ~n22487 & ~n22488;
  assign n22490 = n22167 & ~n22489;
  assign n22491 = ~n20537 & n22262;
  assign n22492 = n22358 & ~n22482;
  assign n22493 = n22270 & ~n22489;
  assign n22494 = ~n22491 & ~n22492;
  assign n22495 = ~n22493 & n22494;
  assign n22496 = n22264 & ~n22495;
  assign n22497 = n22476 & n22485;
  assign n22498 = ~n22490 & n22497;
  assign n2851 = n22496 | ~n22498;
  assign n22500 = P4_ADDR_REG_13_ & n22163;
  assign n22501 = ~n20468 & n22268;
  assign n22502 = ~n22500 & ~n22501;
  assign n22503 = P4_REG2_REG_13_ & n20468;
  assign n22504 = ~P4_REG2_REG_13_ & ~n20468;
  assign n22505 = ~n22503 & ~n22504;
  assign n22506 = n22338 & ~n22505;
  assign n22507 = ~n22338 & n22505;
  assign n22508 = ~n22506 & ~n22507;
  assign n22509 = n22357 & ~n22508;
  assign n22510 = P4_REG3_REG_13_ & ~P4_STATE_REG;
  assign n22511 = ~n22509 & ~n22510;
  assign n22512 = ~n22227 & ~n22228;
  assign n22513 = ~n20468 & ~n22512;
  assign n22514 = n20468 & n22512;
  assign n22515 = ~n22513 & ~n22514;
  assign n22516 = n22167 & ~n22515;
  assign n22517 = ~n20468 & n22262;
  assign n22518 = n22358 & ~n22508;
  assign n22519 = n22270 & ~n22515;
  assign n22520 = ~n22517 & ~n22518;
  assign n22521 = ~n22519 & n22520;
  assign n22522 = n22264 & ~n22521;
  assign n22523 = n22502 & n22511;
  assign n22524 = ~n22516 & n22523;
  assign n2856 = n22522 | ~n22524;
  assign n22526 = P4_REG2_REG_12_ & n20394;
  assign n22527 = ~P4_REG2_REG_12_ & ~n20394;
  assign n22528 = ~n22526 & ~n22527;
  assign n22529 = n22336 & ~n22528;
  assign n22530 = ~n22336 & n22528;
  assign n22531 = ~n22529 & ~n22530;
  assign n22532 = n22357 & ~n22531;
  assign n22533 = P4_REG3_REG_12_ & ~P4_STATE_REG;
  assign n22534 = ~n22532 & ~n22533;
  assign n22535 = P4_ADDR_REG_12_ & n22163;
  assign n22536 = ~n20394 & n22268;
  assign n22537 = P4_REG1_REG_12_ & n20394;
  assign n22538 = ~P4_REG1_REG_12_ & ~n20394;
  assign n22539 = ~n22537 & ~n22538;
  assign n22540 = n22224 & ~n22539;
  assign n22541 = ~n22224 & n22539;
  assign n22542 = ~n22540 & ~n22541;
  assign n22543 = n22167 & ~n22542;
  assign n22544 = ~n22535 & ~n22536;
  assign n22545 = ~n22543 & n22544;
  assign n22546 = ~n20394 & n22262;
  assign n22547 = n22358 & ~n22531;
  assign n22548 = n22270 & ~n22542;
  assign n22549 = ~n22546 & ~n22547;
  assign n22550 = ~n22548 & n22549;
  assign n22551 = n22264 & ~n22550;
  assign n22552 = n22534 & n22545;
  assign n2861 = n22551 | ~n22552;
  assign n22554 = P4_REG2_REG_11_ & n20317;
  assign n22555 = ~P4_REG2_REG_11_ & ~n20317;
  assign n22556 = ~n22554 & ~n22555;
  assign n22557 = n22334 & ~n22556;
  assign n22558 = ~n22334 & n22556;
  assign n22559 = ~n22557 & ~n22558;
  assign n22560 = n22357 & ~n22559;
  assign n22561 = P4_REG3_REG_11_ & ~P4_STATE_REG;
  assign n22562 = ~n22560 & ~n22561;
  assign n22563 = P4_ADDR_REG_11_ & n22163;
  assign n22564 = ~n20317 & n22268;
  assign n22565 = P4_REG1_REG_11_ & n20317;
  assign n22566 = ~P4_REG1_REG_11_ & ~n20317;
  assign n22567 = ~n22565 & ~n22566;
  assign n22568 = n22222 & ~n22567;
  assign n22569 = ~n22222 & n22567;
  assign n22570 = ~n22568 & ~n22569;
  assign n22571 = n22167 & ~n22570;
  assign n22572 = ~n22563 & ~n22564;
  assign n22573 = ~n22571 & n22572;
  assign n22574 = ~n20317 & n22262;
  assign n22575 = n22358 & ~n22559;
  assign n22576 = n22270 & ~n22570;
  assign n22577 = ~n22574 & ~n22575;
  assign n22578 = ~n22576 & n22577;
  assign n22579 = n22264 & ~n22578;
  assign n22580 = n22562 & n22573;
  assign n2866 = n22579 | ~n22580;
  assign n22582 = P4_ADDR_REG_10_ & n22163;
  assign n22583 = ~n20251 & n22268;
  assign n22584 = ~n22582 & ~n22583;
  assign n22585 = P4_REG2_REG_10_ & n20251;
  assign n22586 = ~P4_REG2_REG_10_ & ~n20251;
  assign n22587 = ~n22585 & ~n22586;
  assign n22588 = n22332 & ~n22587;
  assign n22589 = ~n22332 & n22587;
  assign n22590 = ~n22588 & ~n22589;
  assign n22591 = n22357 & ~n22590;
  assign n22592 = P4_REG3_REG_10_ & ~P4_STATE_REG;
  assign n22593 = ~n22591 & ~n22592;
  assign n22594 = ~n22219 & ~n22220;
  assign n22595 = ~n20251 & ~n22594;
  assign n22596 = n20251 & n22594;
  assign n22597 = ~n22595 & ~n22596;
  assign n22598 = n22167 & ~n22597;
  assign n22599 = ~n20251 & n22262;
  assign n22600 = n22358 & ~n22590;
  assign n22601 = n22270 & ~n22597;
  assign n22602 = ~n22599 & ~n22600;
  assign n22603 = ~n22601 & n22602;
  assign n22604 = n22264 & ~n22603;
  assign n22605 = n22584 & n22593;
  assign n22606 = ~n22598 & n22605;
  assign n2871 = n22604 | ~n22606;
  assign n22608 = P4_REG2_REG_9_ & n20184;
  assign n22609 = ~P4_REG2_REG_9_ & ~n20184;
  assign n22610 = ~n22608 & ~n22609;
  assign n22611 = n22330 & ~n22610;
  assign n22612 = ~n22330 & n22610;
  assign n22613 = ~n22611 & ~n22612;
  assign n22614 = n22357 & ~n22613;
  assign n22615 = P4_REG3_REG_9_ & ~P4_STATE_REG;
  assign n22616 = ~n22614 & ~n22615;
  assign n22617 = P4_ADDR_REG_9_ & n22163;
  assign n22618 = ~n20184 & n22268;
  assign n22619 = P4_REG1_REG_9_ & n20184;
  assign n22620 = ~P4_REG1_REG_9_ & ~n20184;
  assign n22621 = ~n22619 & ~n22620;
  assign n22622 = n22216 & ~n22621;
  assign n22623 = ~n22216 & n22621;
  assign n22624 = ~n22622 & ~n22623;
  assign n22625 = n22167 & ~n22624;
  assign n22626 = ~n22617 & ~n22618;
  assign n22627 = ~n22625 & n22626;
  assign n22628 = ~n20184 & n22262;
  assign n22629 = n22358 & ~n22613;
  assign n22630 = n22270 & ~n22624;
  assign n22631 = ~n22628 & ~n22629;
  assign n22632 = ~n22630 & n22631;
  assign n22633 = n22264 & ~n22632;
  assign n22634 = n22616 & n22627;
  assign n2876 = n22633 | ~n22634;
  assign n22636 = P4_ADDR_REG_8_ & n22163;
  assign n22637 = ~n20113 & n22268;
  assign n22638 = ~n22636 & ~n22637;
  assign n22639 = P4_REG2_REG_8_ & n20113;
  assign n22640 = ~P4_REG2_REG_8_ & ~n20113;
  assign n22641 = ~n22639 & ~n22640;
  assign n22642 = n22328 & ~n22641;
  assign n22643 = ~n22328 & n22641;
  assign n22644 = ~n22642 & ~n22643;
  assign n22645 = n22357 & ~n22644;
  assign n22646 = P4_REG3_REG_8_ & ~P4_STATE_REG;
  assign n22647 = ~n22645 & ~n22646;
  assign n22648 = ~n22213 & ~n22214;
  assign n22649 = ~n20113 & ~n22648;
  assign n22650 = n20113 & n22648;
  assign n22651 = ~n22649 & ~n22650;
  assign n22652 = n22167 & ~n22651;
  assign n22653 = ~n20113 & n22262;
  assign n22654 = n22358 & ~n22644;
  assign n22655 = n22270 & ~n22651;
  assign n22656 = ~n22653 & ~n22654;
  assign n22657 = ~n22655 & n22656;
  assign n22658 = n22264 & ~n22657;
  assign n22659 = n22638 & n22647;
  assign n22660 = ~n22652 & n22659;
  assign n2881 = n22658 | ~n22660;
  assign n22662 = P4_REG2_REG_7_ & n20044;
  assign n22663 = ~P4_REG2_REG_7_ & ~n20044;
  assign n22664 = ~n22662 & ~n22663;
  assign n22665 = n22326 & ~n22664;
  assign n22666 = ~n22326 & n22664;
  assign n22667 = ~n22665 & ~n22666;
  assign n22668 = n22357 & ~n22667;
  assign n22669 = P4_REG3_REG_7_ & ~P4_STATE_REG;
  assign n22670 = ~n22668 & ~n22669;
  assign n22671 = P4_ADDR_REG_7_ & n22163;
  assign n22672 = ~n20044 & n22268;
  assign n22673 = P4_REG1_REG_7_ & n20044;
  assign n22674 = ~P4_REG1_REG_7_ & ~n20044;
  assign n22675 = ~n22673 & ~n22674;
  assign n22676 = n22210 & ~n22675;
  assign n22677 = ~n22210 & n22675;
  assign n22678 = ~n22676 & ~n22677;
  assign n22679 = n22167 & ~n22678;
  assign n22680 = ~n22671 & ~n22672;
  assign n22681 = ~n22679 & n22680;
  assign n22682 = ~n20044 & n22262;
  assign n22683 = n22358 & ~n22667;
  assign n22684 = n22270 & ~n22678;
  assign n22685 = ~n22682 & ~n22683;
  assign n22686 = ~n22684 & n22685;
  assign n22687 = n22264 & ~n22686;
  assign n22688 = n22670 & n22681;
  assign n2886 = n22687 | ~n22688;
  assign n22690 = P4_REG1_REG_6_ & n19969;
  assign n22691 = ~P4_REG1_REG_6_ & ~n19969;
  assign n22692 = ~n22690 & ~n22691;
  assign n22693 = n22208 & ~n22692;
  assign n22694 = ~n22208 & n22692;
  assign n22695 = ~n22693 & ~n22694;
  assign n22696 = n22167 & ~n22695;
  assign n22697 = ~n19969 & n22268;
  assign n22698 = P4_ADDR_REG_6_ & n22163;
  assign n22699 = P4_REG3_REG_6_ & ~P4_STATE_REG;
  assign n22700 = ~n19969 & n22262;
  assign n22701 = P4_REG2_REG_6_ & n19969;
  assign n22702 = ~P4_REG2_REG_6_ & ~n19969;
  assign n22703 = ~n22701 & ~n22702;
  assign n22704 = n22324 & ~n22703;
  assign n22705 = ~n22324 & n22703;
  assign n22706 = ~n22704 & ~n22705;
  assign n22707 = n22358 & ~n22706;
  assign n22708 = n22270 & ~n22695;
  assign n22709 = ~n22700 & ~n22707;
  assign n22710 = ~n22708 & n22709;
  assign n22711 = n22264 & ~n22710;
  assign n22712 = ~n22699 & ~n22711;
  assign n22713 = n22357 & ~n22706;
  assign n22714 = ~n22696 & ~n22697;
  assign n22715 = ~n22698 & n22714;
  assign n22716 = n22712 & n22715;
  assign n2891 = n22713 | ~n22716;
  assign n22718 = ~n22205 & ~n22206;
  assign n22719 = ~n19905 & ~n22718;
  assign n22720 = n19905 & n22718;
  assign n22721 = ~n22719 & ~n22720;
  assign n22722 = n22167 & ~n22721;
  assign n22723 = ~n19905 & n22268;
  assign n22724 = P4_ADDR_REG_5_ & n22163;
  assign n22725 = P4_REG3_REG_5_ & ~P4_STATE_REG;
  assign n22726 = ~n19905 & n22262;
  assign n22727 = P4_REG2_REG_5_ & n19905;
  assign n22728 = ~P4_REG2_REG_5_ & ~n19905;
  assign n22729 = ~n22727 & ~n22728;
  assign n22730 = n22322 & ~n22729;
  assign n22731 = ~n22322 & n22729;
  assign n22732 = ~n22730 & ~n22731;
  assign n22733 = n22358 & ~n22732;
  assign n22734 = n22270 & ~n22721;
  assign n22735 = ~n22726 & ~n22733;
  assign n22736 = ~n22734 & n22735;
  assign n22737 = n22264 & ~n22736;
  assign n22738 = ~n22725 & ~n22737;
  assign n22739 = n22357 & ~n22732;
  assign n22740 = ~n22722 & ~n22723;
  assign n22741 = ~n22724 & n22740;
  assign n22742 = n22738 & n22741;
  assign n2896 = n22739 | ~n22742;
  assign n22744 = P4_REG1_REG_4_ & n19821;
  assign n22745 = ~P4_REG1_REG_4_ & ~n19821;
  assign n22746 = ~n22744 & ~n22745;
  assign n22747 = n22202 & ~n22746;
  assign n22748 = ~n22202 & n22746;
  assign n22749 = ~n22747 & ~n22748;
  assign n22750 = n22167 & ~n22749;
  assign n22751 = ~n19821 & n22268;
  assign n22752 = P4_ADDR_REG_4_ & n22163;
  assign n22753 = ~n22750 & ~n22751;
  assign n22754 = ~n22752 & n22753;
  assign n22755 = P4_REG3_REG_4_ & ~P4_STATE_REG;
  assign n22756 = P4_REG2_REG_4_ & n19821;
  assign n22757 = ~P4_REG2_REG_4_ & ~n19821;
  assign n22758 = ~n22756 & ~n22757;
  assign n22759 = n22320 & ~n22758;
  assign n22760 = ~n22320 & n22758;
  assign n22761 = ~n22759 & ~n22760;
  assign n22762 = n22357 & ~n22761;
  assign n22763 = ~n19821 & n22262;
  assign n22764 = n22358 & ~n22761;
  assign n22765 = n22270 & ~n22749;
  assign n22766 = ~n22763 & ~n22764;
  assign n22767 = ~n22765 & n22766;
  assign n22768 = n22264 & ~n22767;
  assign n3246 = P4_STATE_REG & n22158;
  assign n22770 = P4_REG2_REG_0_ & n22356;
  assign n22771 = n19564 & n22770;
  assign n22772 = ~P4_REG2_REG_0_ & ~n19557;
  assign n22773 = ~n19560 & ~n22772;
  assign n22774 = ~n19564 & ~n22773;
  assign n22775 = ~n19418 & ~n22257;
  assign n22776 = ~n19599 & n22775;
  assign n22777 = P4_REG1_REG_0_ & n19418;
  assign n22778 = ~n22776 & ~n22777;
  assign n22779 = ~n19479 & n19483;
  assign n22780 = ~n19418 & n22779;
  assign n22781 = ~n19484 & ~n19610;
  assign n22782 = ~n19619 & n22781;
  assign n22783 = ~n19614 & n22782;
  assign n22784 = ~n19418 & ~n22783;
  assign n22785 = ~n22780 & ~n22784;
  assign n22786 = n19483 & n19487;
  assign n22787 = ~n19418 & n22786;
  assign n22788 = n22785 & ~n22787;
  assign n22789 = ~n19567 & ~n22788;
  assign n22790 = n22778 & ~n22789;
  assign n22791 = ~n19613 & ~n22779;
  assign n22792 = ~n22787 & n22791;
  assign n22793 = ~n19418 & ~n22792;
  assign n22794 = ~n22790 & ~n22793;
  assign n22795 = n22790 & n22793;
  assign n22796 = ~n22794 & ~n22795;
  assign n22797 = n22793 & n22796;
  assign n22798 = ~n22793 & ~n22796;
  assign n22799 = ~n22797 & ~n22798;
  assign n22800 = n19418 & ~n19564;
  assign n22801 = ~n19567 & n22775;
  assign n22802 = ~n22800 & ~n22801;
  assign n22803 = ~n19599 & ~n22785;
  assign n22804 = n22802 & ~n22803;
  assign n22805 = ~n22799 & n22804;
  assign n22806 = n22799 & ~n22804;
  assign n22807 = ~n22805 & ~n22806;
  assign n22808 = n19557 & ~n19560;
  assign n22809 = ~n22807 & n22808;
  assign n22810 = ~n22771 & ~n22774;
  assign n22811 = ~n22809 & n22810;
  assign n22812 = n3246 & ~n22811;
  assign n22813 = ~n22768 & ~n22812;
  assign n22814 = ~n22755 & ~n22762;
  assign n22815 = n22813 & n22814;
  assign n2901 = ~n22754 | ~n22815;
  assign n22817 = ~P4_REG1_REG_3_ & n22197;
  assign n22818 = ~n22198 & ~n22817;
  assign n22819 = ~n19767 & ~n22818;
  assign n22820 = n19767 & n22818;
  assign n22821 = ~n22819 & ~n22820;
  assign n22822 = n22167 & ~n22821;
  assign n22823 = ~n19767 & n22268;
  assign n22824 = P4_ADDR_REG_3_ & n22163;
  assign n22825 = P4_REG3_REG_3_ & ~P4_STATE_REG;
  assign n22826 = ~n19767 & n22262;
  assign n22827 = P4_REG2_REG_3_ & n19767;
  assign n22828 = ~P4_REG2_REG_3_ & ~n19767;
  assign n22829 = ~n22827 & ~n22828;
  assign n22830 = n22318 & ~n22829;
  assign n22831 = ~n22318 & n22829;
  assign n22832 = ~n22830 & ~n22831;
  assign n22833 = n22358 & ~n22832;
  assign n22834 = n22270 & ~n22821;
  assign n22835 = ~n22826 & ~n22833;
  assign n22836 = ~n22834 & n22835;
  assign n22837 = n22264 & ~n22836;
  assign n22838 = ~n22825 & ~n22837;
  assign n22839 = n22357 & ~n22832;
  assign n22840 = ~n22822 & ~n22823;
  assign n22841 = ~n22824 & n22840;
  assign n22842 = n22838 & n22841;
  assign n2906 = n22839 | ~n22842;
  assign n22844 = P4_REG1_REG_2_ & n19696;
  assign n22845 = ~P4_REG1_REG_2_ & ~n19696;
  assign n22846 = ~n22844 & ~n22845;
  assign n22847 = n22195 & ~n22846;
  assign n22848 = ~n22195 & n22846;
  assign n22849 = ~n22847 & ~n22848;
  assign n22850 = n22167 & ~n22849;
  assign n22851 = ~n19696 & n22268;
  assign n22852 = P4_ADDR_REG_2_ & n22163;
  assign n22853 = ~n22850 & ~n22851;
  assign n22854 = ~n22852 & n22853;
  assign n22855 = P4_REG3_REG_2_ & ~P4_STATE_REG;
  assign n22856 = P4_REG2_REG_2_ & n19696;
  assign n22857 = ~P4_REG2_REG_2_ & ~n19696;
  assign n22858 = ~n22856 & ~n22857;
  assign n22859 = n22316 & ~n22858;
  assign n22860 = ~n22316 & n22858;
  assign n22861 = ~n22859 & ~n22860;
  assign n22862 = n22357 & ~n22861;
  assign n22863 = ~n19696 & n22262;
  assign n22864 = n22358 & ~n22861;
  assign n22865 = n22270 & ~n22849;
  assign n22866 = ~n22863 & ~n22864;
  assign n22867 = ~n22865 & n22866;
  assign n22868 = n22264 & ~n22867;
  assign n22869 = ~n22812 & ~n22868;
  assign n22870 = ~n22855 & ~n22862;
  assign n22871 = n22869 & n22870;
  assign n2911 = ~n22854 | ~n22871;
  assign n22873 = n19640 & n22191;
  assign n22874 = ~n19640 & ~n22191;
  assign n22875 = ~n22873 & ~n22874;
  assign n22876 = ~P4_REG1_REG_1_ & ~n22875;
  assign n22877 = n19640 & ~n22191;
  assign n22878 = P4_REG1_REG_1_ & n22877;
  assign n22879 = ~n19640 & n22192;
  assign n22880 = ~n22876 & ~n22878;
  assign n22881 = ~n22879 & n22880;
  assign n22882 = n22167 & ~n22881;
  assign n22883 = ~n19640 & n22268;
  assign n22884 = P4_ADDR_REG_1_ & n22163;
  assign n22885 = P4_REG3_REG_1_ & ~P4_STATE_REG;
  assign n22886 = ~n19640 & n22262;
  assign n22887 = P4_REG2_REG_1_ & n22313;
  assign n22888 = ~n19640 & ~n22312;
  assign n22889 = ~P4_REG2_REG_1_ & n22888;
  assign n22890 = ~n22887 & ~n22889;
  assign n22891 = ~P4_REG2_REG_1_ & n22312;
  assign n22892 = P4_REG2_REG_1_ & ~n22312;
  assign n22893 = ~n22891 & ~n22892;
  assign n22894 = n19640 & ~n22893;
  assign n22895 = n22890 & ~n22894;
  assign n22896 = n22358 & ~n22895;
  assign n22897 = n22270 & ~n22881;
  assign n22898 = ~n22886 & ~n22896;
  assign n22899 = ~n22897 & n22898;
  assign n22900 = n22264 & ~n22899;
  assign n22901 = ~n22885 & ~n22900;
  assign n22902 = n22357 & ~n22895;
  assign n22903 = ~n22882 & ~n22883;
  assign n22904 = ~n22884 & n22903;
  assign n22905 = n22901 & n22904;
  assign n2916 = n22902 | ~n22905;
  assign n22907 = P4_REG1_REG_0_ & n19564;
  assign n22908 = ~P4_REG1_REG_0_ & ~n19564;
  assign n22909 = ~n22907 & ~n22908;
  assign n22910 = n22167 & ~n22909;
  assign n22911 = ~n19564 & n22268;
  assign n22912 = P4_ADDR_REG_0_ & n22163;
  assign n22913 = P4_REG3_REG_0_ & ~P4_STATE_REG;
  assign n22914 = ~n19564 & n22262;
  assign n22915 = P4_REG2_REG_0_ & n19564;
  assign n22916 = ~P4_REG2_REG_0_ & ~n19564;
  assign n22917 = ~n22915 & ~n22916;
  assign n22918 = n22358 & ~n22917;
  assign n22919 = n22270 & ~n22909;
  assign n22920 = ~n22914 & ~n22918;
  assign n22921 = ~n22919 & n22920;
  assign n22922 = n22264 & ~n22921;
  assign n22923 = ~n22913 & ~n22922;
  assign n22924 = n22357 & ~n22917;
  assign n22925 = ~n22910 & ~n22911;
  assign n22926 = ~n22912 & n22925;
  assign n22927 = n22923 & n22926;
  assign n2921 = n22924 | ~n22927;
  assign n22929 = ~n19599 & n3246;
  assign n22930 = P4_DATAO_REG_0_ & ~n3246;
  assign n2926 = n22929 | n22930;
  assign n22932 = ~n19591 & n3246;
  assign n22933 = P4_DATAO_REG_1_ & ~n3246;
  assign n2931 = n22932 | n22933;
  assign n22935 = ~n19659 & n3246;
  assign n22936 = P4_DATAO_REG_2_ & ~n3246;
  assign n2936 = n22935 | n22936;
  assign n22938 = ~n19720 & n3246;
  assign n22939 = P4_DATAO_REG_3_ & ~n3246;
  assign n2941 = n22938 | n22939;
  assign n22941 = ~n19763 & n3246;
  assign n22942 = P4_DATAO_REG_4_ & ~n3246;
  assign n2946 = n22941 | n22942;
  assign n22944 = ~n19851 & n3246;
  assign n22945 = P4_DATAO_REG_5_ & ~n3246;
  assign n2951 = n22944 | n22945;
  assign n22947 = ~n19901 & n3246;
  assign n22948 = P4_DATAO_REG_6_ & ~n3246;
  assign n2956 = n22947 | n22948;
  assign n22950 = ~n19965 & n3246;
  assign n22951 = P4_DATAO_REG_7_ & ~n3246;
  assign n2961 = n22950 | n22951;
  assign n22953 = ~n20040 & n3246;
  assign n22954 = P4_DATAO_REG_8_ & ~n3246;
  assign n2966 = n22953 | n22954;
  assign n22956 = ~n20109 & n3246;
  assign n22957 = P4_DATAO_REG_9_ & ~n3246;
  assign n2971 = n22956 | n22957;
  assign n22959 = ~n20178 & n3246;
  assign n22960 = P4_DATAO_REG_10_ & ~n3246;
  assign n2976 = n22959 | n22960;
  assign n22962 = ~n20247 & n3246;
  assign n22963 = P4_DATAO_REG_11_ & ~n3246;
  assign n2981 = n22962 | n22963;
  assign n22965 = ~n20311 & n3246;
  assign n22966 = P4_DATAO_REG_12_ & ~n3246;
  assign n2986 = n22965 | n22966;
  assign n22968 = ~n20390 & n3246;
  assign n22969 = P4_DATAO_REG_13_ & ~n3246;
  assign n2991 = n22968 | n22969;
  assign n22971 = ~n20462 & n3246;
  assign n22972 = P4_DATAO_REG_14_ & ~n3246;
  assign n2996 = n22971 | n22972;
  assign n22974 = ~n20533 & n3246;
  assign n22975 = P4_DATAO_REG_15_ & ~n3246;
  assign n3001 = n22974 | n22975;
  assign n22977 = ~n20602 & n3246;
  assign n22978 = P4_DATAO_REG_16_ & ~n3246;
  assign n3006 = n22977 | n22978;
  assign n22980 = ~n20670 & n3246;
  assign n22981 = P4_DATAO_REG_17_ & ~n3246;
  assign n3011 = n22980 | n22981;
  assign n22983 = ~n20742 & n3246;
  assign n22984 = P4_DATAO_REG_18_ & ~n3246;
  assign n3016 = n22983 | n22984;
  assign n22986 = ~n20818 & n3246;
  assign n22987 = P4_DATAO_REG_19_ & ~n3246;
  assign n3021 = n22986 | n22987;
  assign n22989 = ~n20889 & n3246;
  assign n22990 = P4_DATAO_REG_20_ & ~n3246;
  assign n3026 = n22989 | n22990;
  assign n22992 = ~n20957 & n3246;
  assign n22993 = P4_DATAO_REG_21_ & ~n3246;
  assign n3031 = n22992 | n22993;
  assign n22995 = ~n21021 & n3246;
  assign n22996 = P4_DATAO_REG_22_ & ~n3246;
  assign n3036 = n22995 | n22996;
  assign n22998 = ~n21087 & n3246;
  assign n22999 = P4_DATAO_REG_23_ & ~n3246;
  assign n3041 = n22998 | n22999;
  assign n23001 = ~n21154 & n3246;
  assign n23002 = P4_DATAO_REG_24_ & ~n3246;
  assign n3046 = n23001 | n23002;
  assign n23004 = ~n21220 & n3246;
  assign n23005 = P4_DATAO_REG_25_ & ~n3246;
  assign n3051 = n23004 | n23005;
  assign n23007 = ~n21289 & n3246;
  assign n23008 = P4_DATAO_REG_26_ & ~n3246;
  assign n3056 = n23007 | n23008;
  assign n23010 = ~n21353 & n3246;
  assign n23011 = P4_DATAO_REG_27_ & ~n3246;
  assign n3061 = n23010 | n23011;
  assign n23013 = ~n21420 & n3246;
  assign n23014 = P4_DATAO_REG_28_ & ~n3246;
  assign n3066 = n23013 | n23014;
  assign n23016 = ~n21483 & n3246;
  assign n23017 = P4_DATAO_REG_29_ & ~n3246;
  assign n3071 = n23016 | n23017;
  assign n23019 = ~n21574 & n3246;
  assign n23020 = P4_DATAO_REG_30_ & ~n3246;
  assign n3076 = n23019 | n23020;
  assign n23022 = ~n21620 & n3246;
  assign n23023 = P4_DATAO_REG_31_ & ~n3246;
  assign n3081 = n23022 | n23023;
  assign n23025 = ~n19407 & ~n19487;
  assign n23026 = ~n19487 & n19616;
  assign n23027 = n22356 & n23026;
  assign n23028 = n19407 & ~n23027;
  assign n23029 = P4_STATE_REG & ~n22158;
  assign n23030 = ~n23025 & ~n23028;
  assign n23031 = n23029 & n23030;
  assign n23032 = P4_B_REG & ~n23031;
  assign n23033 = n19407 & n19609;
  assign n23034 = ~n19407 & n19609;
  assign n23035 = n21632 & n23034;
  assign n23036 = n19487 & ~n21620;
  assign n23037 = ~n23035 & ~n23036;
  assign n23038 = ~n21574 & n21620;
  assign n23039 = ~n21620 & ~n23038;
  assign n23040 = n21574 & ~n21620;
  assign n23041 = ~n23038 & ~n23040;
  assign n23042 = n23038 & n23041;
  assign n23043 = ~n23039 & ~n23042;
  assign n23044 = ~n19476 & ~n23043;
  assign n23045 = n23037 & ~n23044;
  assign n23046 = ~n21620 & n23034;
  assign n23047 = ~n19609 & n21632;
  assign n23048 = ~n23046 & ~n23047;
  assign n23049 = n23033 & n23045;
  assign n23050 = ~n23048 & n23049;
  assign n23051 = ~n23033 & ~n23045;
  assign n23052 = n23048 & n23051;
  assign n23053 = ~n23050 & ~n23052;
  assign n23054 = n23045 & ~n23048;
  assign n23055 = ~n23045 & n23048;
  assign n23056 = ~n23054 & ~n23055;
  assign n23057 = n23053 & ~n23056;
  assign n23058 = n21614 & n23034;
  assign n23059 = n19487 & ~n21574;
  assign n23060 = ~n23058 & ~n23059;
  assign n23061 = ~n21574 & ~n23038;
  assign n23062 = n21574 & n23038;
  assign n23063 = ~n23061 & ~n23062;
  assign n23064 = ~n19476 & ~n23063;
  assign n23065 = n23060 & ~n23064;
  assign n23066 = ~n21574 & n23034;
  assign n23067 = ~n19609 & n21614;
  assign n23068 = ~n23066 & ~n23067;
  assign n23069 = ~n23065 & n23068;
  assign n23070 = n23053 & n23069;
  assign n23071 = ~n23057 & ~n23070;
  assign n23072 = n23065 & ~n23068;
  assign n23073 = ~n21483 & n23034;
  assign n23074 = ~n19609 & n21547;
  assign n23075 = n19407 & ~n21420;
  assign n23076 = ~n23073 & ~n23074;
  assign n23077 = ~n23075 & n23076;
  assign n23078 = ~n21483 & ~n23038;
  assign n23079 = ~n21483 & n23038;
  assign n23080 = ~n23078 & ~n23079;
  assign n23081 = ~n19476 & ~n23080;
  assign n23082 = n19487 & ~n21483;
  assign n23083 = n21547 & n23034;
  assign n23084 = ~n19407 & ~n23083;
  assign n23085 = ~n23082 & n23084;
  assign n23086 = ~n23081 & n23085;
  assign n23087 = ~n23077 & n23086;
  assign n23088 = n23053 & ~n23072;
  assign n23089 = ~n23087 & n23088;
  assign n23090 = ~n21289 & ~n23038;
  assign n23091 = ~n21289 & n23038;
  assign n23092 = ~n23090 & ~n23091;
  assign n23093 = ~n19476 & ~n23092;
  assign n23094 = n19487 & ~n21289;
  assign n23095 = n21355 & n23034;
  assign n23096 = ~n19407 & ~n23095;
  assign n23097 = ~n23094 & n23096;
  assign n23098 = ~n23093 & n23097;
  assign n23099 = ~n21289 & n23034;
  assign n23100 = ~n19609 & n21355;
  assign n23101 = n19407 & ~n21220;
  assign n23102 = ~n23099 & ~n23100;
  assign n23103 = ~n23101 & n23102;
  assign n23104 = ~n23098 & n23103;
  assign n23105 = n19407 & ~n21154;
  assign n23106 = ~n19609 & n21293;
  assign n23107 = ~n21220 & n23034;
  assign n23108 = ~n23105 & ~n23106;
  assign n23109 = ~n23107 & n23108;
  assign n23110 = ~n21220 & ~n23038;
  assign n23111 = ~n21220 & n23038;
  assign n23112 = ~n23110 & ~n23111;
  assign n23113 = ~n19476 & ~n23112;
  assign n23114 = n19487 & ~n21220;
  assign n23115 = n21293 & n23034;
  assign n23116 = ~n19407 & ~n23115;
  assign n23117 = ~n23114 & n23116;
  assign n23118 = ~n23113 & n23117;
  assign n23119 = ~n23109 & n23118;
  assign n23120 = n23098 & ~n23103;
  assign n23121 = ~n23119 & ~n23120;
  assign n23122 = ~n21154 & ~n23038;
  assign n23123 = ~n21154 & n23038;
  assign n23124 = ~n23122 & ~n23123;
  assign n23125 = ~n19476 & ~n23124;
  assign n23126 = n19487 & ~n21154;
  assign n23127 = n21222 & n23034;
  assign n23128 = ~n19407 & ~n23127;
  assign n23129 = ~n23126 & n23128;
  assign n23130 = ~n23125 & n23129;
  assign n23131 = ~n21154 & n23034;
  assign n23132 = ~n19609 & n21222;
  assign n23133 = n19407 & ~n21087;
  assign n23134 = ~n23131 & ~n23132;
  assign n23135 = ~n23133 & n23134;
  assign n23136 = ~n23130 & n23135;
  assign n23137 = n19407 & ~n21021;
  assign n23138 = ~n19609 & n21158;
  assign n23139 = ~n21087 & n23034;
  assign n23140 = ~n23137 & ~n23138;
  assign n23141 = ~n23139 & n23140;
  assign n23142 = ~n21087 & ~n23038;
  assign n23143 = ~n21087 & n23038;
  assign n23144 = ~n23142 & ~n23143;
  assign n23145 = ~n19476 & ~n23144;
  assign n23146 = n19487 & ~n21087;
  assign n23147 = n21158 & n23034;
  assign n23148 = ~n19407 & ~n23147;
  assign n23149 = ~n23146 & n23148;
  assign n23150 = ~n23145 & n23149;
  assign n23151 = ~n23141 & n23150;
  assign n23152 = n23130 & ~n23135;
  assign n23153 = ~n23151 & ~n23152;
  assign n23154 = ~n21021 & ~n23038;
  assign n23155 = ~n21021 & n23038;
  assign n23156 = ~n23154 & ~n23155;
  assign n23157 = ~n19476 & ~n23156;
  assign n23158 = n19487 & ~n21021;
  assign n23159 = n21089 & n23034;
  assign n23160 = ~n19407 & ~n23159;
  assign n23161 = ~n23158 & n23160;
  assign n23162 = ~n23157 & n23161;
  assign n23163 = ~n21021 & n23034;
  assign n23164 = ~n19609 & n21089;
  assign n23165 = n19407 & ~n20957;
  assign n23166 = ~n23163 & ~n23164;
  assign n23167 = ~n23165 & n23166;
  assign n23168 = ~n23162 & n23167;
  assign n23169 = n19407 & ~n20889;
  assign n23170 = ~n19609 & n21025;
  assign n23171 = ~n20957 & n23034;
  assign n23172 = ~n23169 & ~n23170;
  assign n23173 = ~n23171 & n23172;
  assign n23174 = ~n20957 & ~n23038;
  assign n23175 = ~n20957 & n23038;
  assign n23176 = ~n23174 & ~n23175;
  assign n23177 = ~n19476 & ~n23176;
  assign n23178 = n19487 & ~n20957;
  assign n23179 = n21025 & n23034;
  assign n23180 = ~n19407 & ~n23179;
  assign n23181 = ~n23178 & n23180;
  assign n23182 = ~n23177 & n23181;
  assign n23183 = ~n23173 & n23182;
  assign n23184 = n23162 & ~n23167;
  assign n23185 = ~n23183 & ~n23184;
  assign n23186 = ~n20889 & ~n23038;
  assign n23187 = ~n20889 & n23038;
  assign n23188 = ~n23186 & ~n23187;
  assign n23189 = ~n19476 & ~n23188;
  assign n23190 = n19487 & ~n20889;
  assign n23191 = n20959 & n23034;
  assign n23192 = ~n19407 & ~n23191;
  assign n23193 = ~n23190 & n23192;
  assign n23194 = ~n23189 & n23193;
  assign n23195 = ~n20889 & n23034;
  assign n23196 = ~n19609 & n20959;
  assign n23197 = n19407 & ~n20818;
  assign n23198 = ~n23195 & ~n23196;
  assign n23199 = ~n23197 & n23198;
  assign n23200 = ~n23194 & n23199;
  assign n23201 = n23173 & ~n23182;
  assign n23202 = ~n23200 & ~n23201;
  assign n23203 = n19407 & ~n20742;
  assign n23204 = ~n19609 & ~n20895;
  assign n23205 = ~n20818 & n23034;
  assign n23206 = ~n23203 & ~n23204;
  assign n23207 = ~n23205 & n23206;
  assign n23208 = ~n20818 & ~n23038;
  assign n23209 = ~n20818 & n23038;
  assign n23210 = ~n23208 & ~n23209;
  assign n23211 = ~n19476 & ~n23210;
  assign n23212 = ~n20895 & n23034;
  assign n23213 = n19487 & ~n20818;
  assign n23214 = ~n19407 & ~n23212;
  assign n23215 = ~n23213 & n23214;
  assign n23216 = ~n23211 & n23215;
  assign n23217 = ~n23207 & n23216;
  assign n23218 = n23194 & ~n23199;
  assign n23219 = ~n23217 & ~n23218;
  assign n23220 = ~n20742 & ~n23038;
  assign n23221 = ~n20742 & n23038;
  assign n23222 = ~n23220 & ~n23221;
  assign n23223 = ~n19476 & ~n23222;
  assign n23224 = ~n20825 & n23034;
  assign n23225 = n19487 & ~n20742;
  assign n23226 = ~n19407 & ~n23224;
  assign n23227 = ~n23225 & n23226;
  assign n23228 = ~n23223 & n23227;
  assign n23229 = ~n20742 & n23034;
  assign n23230 = ~n19609 & ~n20825;
  assign n23231 = n19407 & ~n20670;
  assign n23232 = ~n23229 & ~n23230;
  assign n23233 = ~n23231 & n23232;
  assign n23234 = ~n23228 & n23233;
  assign n23235 = n23207 & ~n23216;
  assign n23236 = ~n23234 & ~n23235;
  assign n23237 = n19407 & ~n20602;
  assign n23238 = ~n19609 & ~n20751;
  assign n23239 = ~n20670 & n23034;
  assign n23240 = ~n23237 & ~n23238;
  assign n23241 = ~n23239 & n23240;
  assign n23242 = ~n20670 & ~n23038;
  assign n23243 = ~n20670 & n23038;
  assign n23244 = ~n23242 & ~n23243;
  assign n23245 = ~n19476 & ~n23244;
  assign n23246 = ~n20751 & n23034;
  assign n23247 = n19487 & ~n20670;
  assign n23248 = ~n19407 & ~n23246;
  assign n23249 = ~n23247 & n23248;
  assign n23250 = ~n23245 & n23249;
  assign n23251 = ~n23241 & n23250;
  assign n23252 = n23228 & ~n23233;
  assign n23253 = ~n23251 & ~n23252;
  assign n23254 = ~n20602 & ~n23038;
  assign n23255 = ~n20602 & n23038;
  assign n23256 = ~n23254 & ~n23255;
  assign n23257 = ~n19476 & ~n23256;
  assign n23258 = ~n20677 & n23034;
  assign n23259 = n19487 & ~n20602;
  assign n23260 = ~n19407 & ~n23258;
  assign n23261 = ~n23259 & n23260;
  assign n23262 = ~n23257 & n23261;
  assign n23263 = ~n20602 & n23034;
  assign n23264 = ~n19609 & ~n20677;
  assign n23265 = n19407 & ~n20533;
  assign n23266 = ~n23263 & ~n23264;
  assign n23267 = ~n23265 & n23266;
  assign n23268 = ~n23262 & n23267;
  assign n23269 = n23241 & ~n23250;
  assign n23270 = ~n23268 & ~n23269;
  assign n23271 = n19407 & ~n20462;
  assign n23272 = ~n19609 & ~n20611;
  assign n23273 = ~n20533 & n23034;
  assign n23274 = ~n23271 & ~n23272;
  assign n23275 = ~n23273 & n23274;
  assign n23276 = ~n20533 & ~n23038;
  assign n23277 = ~n20533 & n23038;
  assign n23278 = ~n23276 & ~n23277;
  assign n23279 = ~n19476 & ~n23278;
  assign n23280 = ~n20611 & n23034;
  assign n23281 = n19487 & ~n20533;
  assign n23282 = ~n19407 & ~n23280;
  assign n23283 = ~n23281 & n23282;
  assign n23284 = ~n23279 & n23283;
  assign n23285 = ~n23275 & n23284;
  assign n23286 = n23262 & ~n23267;
  assign n23287 = ~n23285 & ~n23286;
  assign n23288 = ~n20462 & ~n23038;
  assign n23289 = ~n20462 & n23038;
  assign n23290 = ~n23288 & ~n23289;
  assign n23291 = ~n19476 & ~n23290;
  assign n23292 = ~n20540 & n23034;
  assign n23293 = n19487 & ~n20462;
  assign n23294 = ~n19407 & ~n23292;
  assign n23295 = ~n23293 & n23294;
  assign n23296 = ~n23291 & n23295;
  assign n23297 = ~n20462 & n23034;
  assign n23298 = ~n19609 & ~n20540;
  assign n23299 = n19407 & ~n20390;
  assign n23300 = ~n23297 & ~n23298;
  assign n23301 = ~n23299 & n23300;
  assign n23302 = ~n23296 & n23301;
  assign n23303 = n23275 & ~n23284;
  assign n23304 = ~n23302 & ~n23303;
  assign n23305 = n19407 & ~n20311;
  assign n23306 = ~n19609 & ~n20471;
  assign n23307 = ~n20390 & n23034;
  assign n23308 = ~n23305 & ~n23306;
  assign n23309 = ~n23307 & n23308;
  assign n23310 = ~n20390 & ~n23038;
  assign n23311 = ~n20390 & n23038;
  assign n23312 = ~n23310 & ~n23311;
  assign n23313 = ~n19476 & ~n23312;
  assign n23314 = ~n20471 & n23034;
  assign n23315 = n19487 & ~n20390;
  assign n23316 = ~n19407 & ~n23314;
  assign n23317 = ~n23315 & n23316;
  assign n23318 = ~n23313 & n23317;
  assign n23319 = ~n23309 & n23318;
  assign n23320 = n23296 & ~n23301;
  assign n23321 = ~n23319 & ~n23320;
  assign n23322 = ~n20311 & ~n23038;
  assign n23323 = ~n20311 & n23038;
  assign n23324 = ~n23322 & ~n23323;
  assign n23325 = ~n19476 & ~n23324;
  assign n23326 = ~n20397 & n23034;
  assign n23327 = n19487 & ~n20311;
  assign n23328 = ~n19407 & ~n23326;
  assign n23329 = ~n23327 & n23328;
  assign n23330 = ~n23325 & n23329;
  assign n23331 = ~n20311 & n23034;
  assign n23332 = ~n19609 & ~n20397;
  assign n23333 = n19407 & ~n20247;
  assign n23334 = ~n23331 & ~n23332;
  assign n23335 = ~n23333 & n23334;
  assign n23336 = ~n23330 & n23335;
  assign n23337 = n23309 & ~n23318;
  assign n23338 = ~n23336 & ~n23337;
  assign n23339 = n19407 & ~n20178;
  assign n23340 = ~n19609 & ~n20320;
  assign n23341 = ~n20247 & n23034;
  assign n23342 = ~n23339 & ~n23340;
  assign n23343 = ~n23341 & n23342;
  assign n23344 = ~n20247 & ~n23038;
  assign n23345 = ~n20247 & n23038;
  assign n23346 = ~n23344 & ~n23345;
  assign n23347 = ~n19476 & ~n23346;
  assign n23348 = ~n20320 & n23034;
  assign n23349 = n19487 & ~n20247;
  assign n23350 = ~n19407 & ~n23348;
  assign n23351 = ~n23349 & n23350;
  assign n23352 = ~n23347 & n23351;
  assign n23353 = ~n23343 & n23352;
  assign n23354 = n23330 & ~n23335;
  assign n23355 = ~n23353 & ~n23354;
  assign n23356 = ~n20178 & ~n23038;
  assign n23357 = ~n20178 & n23038;
  assign n23358 = ~n23356 & ~n23357;
  assign n23359 = ~n19476 & ~n23358;
  assign n23360 = ~n20254 & n23034;
  assign n23361 = n19487 & ~n20178;
  assign n23362 = ~n19407 & ~n23360;
  assign n23363 = ~n23361 & n23362;
  assign n23364 = ~n23359 & n23363;
  assign n23365 = ~n20178 & n23034;
  assign n23366 = ~n19609 & ~n20254;
  assign n23367 = n19407 & ~n20109;
  assign n23368 = ~n23365 & ~n23366;
  assign n23369 = ~n23367 & n23368;
  assign n23370 = ~n23364 & n23369;
  assign n23371 = n23343 & ~n23352;
  assign n23372 = ~n23370 & ~n23371;
  assign n23373 = ~n20109 & n23034;
  assign n23374 = ~n19609 & ~n20187;
  assign n23375 = n19407 & ~n20040;
  assign n23376 = ~n23373 & ~n23374;
  assign n23377 = ~n23375 & n23376;
  assign n23378 = ~n20109 & ~n23038;
  assign n23379 = ~n20109 & n23038;
  assign n23380 = ~n23378 & ~n23379;
  assign n23381 = ~n19476 & ~n23380;
  assign n23382 = ~n20187 & n23034;
  assign n23383 = n19487 & ~n20109;
  assign n23384 = ~n19407 & ~n23382;
  assign n23385 = ~n23383 & n23384;
  assign n23386 = ~n23381 & n23385;
  assign n23387 = ~n23377 & n23386;
  assign n23388 = n23364 & ~n23369;
  assign n23389 = ~n23387 & ~n23388;
  assign n23390 = ~n20040 & ~n23038;
  assign n23391 = ~n20040 & n23038;
  assign n23392 = ~n23390 & ~n23391;
  assign n23393 = ~n19476 & ~n23392;
  assign n23394 = ~n20116 & n23034;
  assign n23395 = n19487 & ~n20040;
  assign n23396 = ~n19407 & ~n23394;
  assign n23397 = ~n23395 & n23396;
  assign n23398 = ~n23393 & n23397;
  assign n23399 = ~n20040 & n23034;
  assign n23400 = ~n19609 & ~n20116;
  assign n23401 = n19407 & ~n19965;
  assign n23402 = ~n23399 & ~n23400;
  assign n23403 = ~n23401 & n23402;
  assign n23404 = ~n23398 & n23403;
  assign n23405 = n23377 & ~n23386;
  assign n23406 = ~n23404 & ~n23405;
  assign n23407 = ~n19965 & n23034;
  assign n23408 = ~n19609 & ~n20047;
  assign n23409 = n19407 & ~n19901;
  assign n23410 = ~n23407 & ~n23408;
  assign n23411 = ~n23409 & n23410;
  assign n23412 = ~n19965 & ~n23038;
  assign n23413 = ~n19965 & n23038;
  assign n23414 = ~n23412 & ~n23413;
  assign n23415 = ~n19476 & ~n23414;
  assign n23416 = ~n20047 & n23034;
  assign n23417 = n19487 & ~n19965;
  assign n23418 = ~n19407 & ~n23416;
  assign n23419 = ~n23417 & n23418;
  assign n23420 = ~n23415 & n23419;
  assign n23421 = ~n23411 & n23420;
  assign n23422 = n23398 & ~n23403;
  assign n23423 = ~n23421 & ~n23422;
  assign n23424 = ~n19901 & ~n23038;
  assign n23425 = ~n19901 & n23038;
  assign n23426 = ~n23424 & ~n23425;
  assign n23427 = ~n19476 & ~n23426;
  assign n23428 = ~n19972 & n23034;
  assign n23429 = n19487 & ~n19901;
  assign n23430 = ~n19407 & ~n23428;
  assign n23431 = ~n23429 & n23430;
  assign n23432 = ~n23427 & n23431;
  assign n23433 = ~n19901 & n23034;
  assign n23434 = ~n19609 & ~n19972;
  assign n23435 = n19407 & ~n19851;
  assign n23436 = ~n23433 & ~n23434;
  assign n23437 = ~n23435 & n23436;
  assign n23438 = ~n23432 & n23437;
  assign n23439 = n23411 & ~n23420;
  assign n23440 = ~n23438 & ~n23439;
  assign n23441 = ~n19851 & n23034;
  assign n23442 = ~n19609 & ~n19908;
  assign n23443 = n19407 & ~n19763;
  assign n23444 = ~n23441 & ~n23442;
  assign n23445 = ~n23443 & n23444;
  assign n23446 = ~n19851 & ~n23038;
  assign n23447 = ~n19851 & n23038;
  assign n23448 = ~n23446 & ~n23447;
  assign n23449 = ~n19476 & ~n23448;
  assign n23450 = ~n19908 & n23034;
  assign n23451 = n19487 & ~n19851;
  assign n23452 = ~n19407 & ~n23450;
  assign n23453 = ~n23451 & n23452;
  assign n23454 = ~n23449 & n23453;
  assign n23455 = ~n23445 & n23454;
  assign n23456 = n23432 & ~n23437;
  assign n23457 = ~n23455 & ~n23456;
  assign n23458 = ~n19763 & ~n23038;
  assign n23459 = ~n19763 & n23038;
  assign n23460 = ~n23458 & ~n23459;
  assign n23461 = ~n19476 & ~n23460;
  assign n23462 = ~n19824 & n23034;
  assign n23463 = n19487 & ~n19763;
  assign n23464 = ~n19407 & ~n23462;
  assign n23465 = ~n23463 & n23464;
  assign n23466 = ~n23461 & n23465;
  assign n23467 = ~n19763 & n23034;
  assign n23468 = ~n19609 & ~n19824;
  assign n23469 = n19407 & ~n19720;
  assign n23470 = ~n23467 & ~n23468;
  assign n23471 = ~n23469 & n23470;
  assign n23472 = ~n23466 & n23471;
  assign n23473 = n23445 & ~n23454;
  assign n23474 = ~n23472 & ~n23473;
  assign n23475 = ~n19720 & n23034;
  assign n23476 = ~n19609 & ~n19770;
  assign n23477 = n19407 & ~n19659;
  assign n23478 = ~n23475 & ~n23476;
  assign n23479 = ~n23477 & n23478;
  assign n23480 = ~n19720 & ~n23038;
  assign n23481 = ~n19720 & n23038;
  assign n23482 = ~n23480 & ~n23481;
  assign n23483 = ~n19476 & ~n23482;
  assign n23484 = ~n19770 & n23034;
  assign n23485 = n19487 & ~n19720;
  assign n23486 = ~n19407 & ~n23484;
  assign n23487 = ~n23485 & n23486;
  assign n23488 = ~n23483 & n23487;
  assign n23489 = ~n23479 & n23488;
  assign n23490 = n23466 & ~n23471;
  assign n23491 = ~n23489 & ~n23490;
  assign n23492 = ~n19659 & ~n23038;
  assign n23493 = ~n19659 & n23038;
  assign n23494 = ~n23492 & ~n23493;
  assign n23495 = ~n19476 & ~n23494;
  assign n23496 = ~n19699 & n23034;
  assign n23497 = n19487 & ~n19659;
  assign n23498 = ~n19407 & ~n23496;
  assign n23499 = ~n23497 & n23498;
  assign n23500 = ~n23495 & n23499;
  assign n23501 = ~n19659 & n23034;
  assign n23502 = ~n19609 & ~n19699;
  assign n23503 = n19407 & ~n19591;
  assign n23504 = ~n23501 & ~n23502;
  assign n23505 = ~n23503 & n23504;
  assign n23506 = ~n23500 & n23505;
  assign n23507 = n23479 & ~n23488;
  assign n23508 = ~n23506 & ~n23507;
  assign n23509 = ~n19591 & n23034;
  assign n23510 = ~n19609 & ~n19643;
  assign n23511 = n19407 & ~n19599;
  assign n23512 = ~n23509 & ~n23510;
  assign n23513 = ~n23511 & n23512;
  assign n23514 = ~n19591 & ~n23038;
  assign n23515 = ~n19591 & n23038;
  assign n23516 = ~n23514 & ~n23515;
  assign n23517 = ~n19476 & ~n23516;
  assign n23518 = ~n19643 & n23034;
  assign n23519 = n19487 & ~n19591;
  assign n23520 = ~n19407 & ~n23518;
  assign n23521 = ~n23519 & n23520;
  assign n23522 = ~n23517 & n23521;
  assign n23523 = ~n23513 & n23522;
  assign n23524 = n23500 & ~n23505;
  assign n23525 = ~n23523 & ~n23524;
  assign n23526 = ~n19599 & n23034;
  assign n23527 = ~n19567 & ~n19609;
  assign n23528 = ~n23526 & ~n23527;
  assign n23529 = ~n19599 & ~n23038;
  assign n23530 = ~n19599 & n23038;
  assign n23531 = ~n23529 & ~n23530;
  assign n23532 = ~n19476 & ~n23531;
  assign n23533 = ~n19567 & n23034;
  assign n23534 = n19487 & ~n19599;
  assign n23535 = ~n19407 & ~n23533;
  assign n23536 = ~n23534 & n23535;
  assign n23537 = ~n23532 & n23536;
  assign n23538 = ~n23528 & n23537;
  assign n23539 = n23513 & ~n23522;
  assign n23540 = n23538 & ~n23539;
  assign n23541 = n23525 & ~n23540;
  assign n23542 = n23508 & ~n23541;
  assign n23543 = n23491 & ~n23542;
  assign n23544 = n23474 & ~n23543;
  assign n23545 = n23457 & ~n23544;
  assign n23546 = n23440 & ~n23545;
  assign n23547 = n23423 & ~n23546;
  assign n23548 = n23406 & ~n23547;
  assign n23549 = n23389 & ~n23548;
  assign n23550 = n23372 & ~n23549;
  assign n23551 = n23355 & ~n23550;
  assign n23552 = n23338 & ~n23551;
  assign n23553 = n23321 & ~n23552;
  assign n23554 = n23304 & ~n23553;
  assign n23555 = n23287 & ~n23554;
  assign n23556 = n23270 & ~n23555;
  assign n23557 = n23253 & ~n23556;
  assign n23558 = n23236 & ~n23557;
  assign n23559 = n23219 & ~n23558;
  assign n23560 = n23202 & ~n23559;
  assign n23561 = n23185 & ~n23560;
  assign n23562 = n23141 & ~n23150;
  assign n23563 = ~n23168 & ~n23561;
  assign n23564 = ~n23562 & n23563;
  assign n23565 = n23153 & ~n23564;
  assign n23566 = n23109 & ~n23118;
  assign n23567 = ~n23136 & ~n23565;
  assign n23568 = ~n23566 & n23567;
  assign n23569 = n23121 & ~n23568;
  assign n23570 = ~n21353 & ~n23038;
  assign n23571 = ~n21353 & n23038;
  assign n23572 = ~n23570 & ~n23571;
  assign n23573 = ~n19476 & ~n23572;
  assign n23574 = n19487 & ~n21353;
  assign n23575 = n21422 & n23034;
  assign n23576 = ~n19407 & ~n23575;
  assign n23577 = ~n23574 & n23576;
  assign n23578 = ~n23573 & n23577;
  assign n23579 = n19407 & ~n21289;
  assign n23580 = ~n19609 & n21422;
  assign n23581 = ~n21353 & n23034;
  assign n23582 = ~n23579 & ~n23580;
  assign n23583 = ~n23581 & n23582;
  assign n23584 = ~n23578 & n23583;
  assign n23585 = ~n23104 & ~n23569;
  assign n23586 = ~n23584 & n23585;
  assign n23587 = n23578 & ~n23583;
  assign n23588 = ~n21420 & n23034;
  assign n23589 = ~n19609 & n21485;
  assign n23590 = n19407 & ~n21353;
  assign n23591 = ~n23588 & ~n23589;
  assign n23592 = ~n23590 & n23591;
  assign n23593 = ~n21420 & ~n23038;
  assign n23594 = ~n21420 & n23038;
  assign n23595 = ~n23593 & ~n23594;
  assign n23596 = ~n19476 & ~n23595;
  assign n23597 = n19487 & ~n21420;
  assign n23598 = n21485 & n23034;
  assign n23599 = ~n19407 & ~n23598;
  assign n23600 = ~n23597 & n23599;
  assign n23601 = ~n23596 & n23600;
  assign n23602 = ~n23592 & n23601;
  assign n23603 = ~n23587 & ~n23602;
  assign n23604 = n23089 & ~n23586;
  assign n23605 = n23603 & n23604;
  assign n23606 = ~n23072 & n23592;
  assign n23607 = ~n23087 & n23606;
  assign n23608 = n23053 & ~n23601;
  assign n23609 = n23607 & n23608;
  assign n23610 = ~n23072 & n23077;
  assign n23611 = n23053 & ~n23086;
  assign n23612 = n23610 & n23611;
  assign n23613 = ~n23609 & ~n23612;
  assign n23614 = n23071 & ~n23605;
  assign n23615 = n23613 & n23614;
  assign n23616 = n19420 & n23027;
  assign n23617 = n23615 & n23616;
  assign n23618 = ~n23032 & ~n23617;
  assign n23619 = ~n19914 & ~n19915;
  assign n23620 = ~n19786 & ~n23619;
  assign n23621 = ~n19703 & n23620;
  assign n23622 = ~n20053 & ~n20054;
  assign n23623 = ~n19995 & ~n23622;
  assign n23624 = ~n20411 & n23623;
  assign n23625 = ~n20757 & ~n20758;
  assign n23626 = n23621 & n23624;
  assign n23627 = ~n20693 & n23626;
  assign n23628 = ~n23625 & n23627;
  assign n23629 = n19567 & n19599;
  assign n23630 = ~n19648 & ~n23629;
  assign n23631 = ~n20617 & ~n20618;
  assign n23632 = ~n19647 & ~n23630;
  assign n23633 = ~n23631 & n23632;
  assign n23634 = ~n20477 & ~n20478;
  assign n23635 = ~n20134 & ~n20201;
  assign n23636 = ~n23634 & n23635;
  assign n23637 = ~n20686 & ~n20687;
  assign n23638 = n23633 & n23636;
  assign n23639 = ~n23637 & n23638;
  assign n23640 = ~n20843 & n23639;
  assign n23641 = n21420 & ~n21485;
  assign n23642 = ~n21555 & ~n23641;
  assign n23643 = ~n21491 & ~n21497;
  assign n23644 = ~n23642 & ~n23643;
  assign n23645 = ~n21228 & ~n21229;
  assign n23646 = ~n21238 & ~n23645;
  assign n23647 = ~n21164 & ~n21165;
  assign n23648 = ~n21095 & ~n21099;
  assign n23649 = ~n23647 & ~n23648;
  assign n23650 = n21289 & ~n21355;
  assign n23651 = ~n21362 & ~n23650;
  assign n23652 = ~n21307 & ~n23651;
  assign n23653 = n23646 & n23649;
  assign n23654 = n23652 & n23653;
  assign n23655 = ~n20260 & ~n20261;
  assign n23656 = ~n19837 & ~n23655;
  assign n23657 = ~n20339 & n23656;
  assign n23658 = ~n20909 & n23657;
  assign n23659 = n21574 & ~n21614;
  assign n23660 = ~n21574 & n21614;
  assign n23661 = ~n23659 & ~n23660;
  assign n23662 = n21620 & ~n21632;
  assign n23663 = ~n21620 & n21632;
  assign n23664 = ~n23662 & ~n23663;
  assign n23665 = ~n20965 & ~n20966;
  assign n23666 = ~n23661 & ~n23664;
  assign n23667 = ~n23665 & n23666;
  assign n23668 = n21483 & ~n21547;
  assign n23669 = ~n21483 & n21547;
  assign n23670 = ~n23668 & ~n23669;
  assign n23671 = n23658 & n23667;
  assign n23672 = ~n23670 & n23671;
  assign n23673 = n23628 & n23640;
  assign n23674 = n23644 & n23673;
  assign n23675 = n23654 & n23674;
  assign n23676 = n23672 & n23675;
  assign n23677 = n19484 & ~n23676;
  assign n23678 = ~n19479 & n23677;
  assign n23679 = n19573 & n23615;
  assign n23680 = ~n19476 & n23679;
  assign n23681 = n21169 & ~n21232;
  assign n23682 = ~n21233 & ~n23681;
  assign n23683 = ~n21300 & n23682;
  assign n23684 = n19921 & ~n19979;
  assign n23685 = ~n20129 & ~n20194;
  assign n23686 = n20334 & ~n20403;
  assign n23687 = ~n20060 & n23685;
  assign n23688 = ~n20267 & n23687;
  assign n23689 = ~n23686 & n23688;
  assign n23690 = ~n19980 & n23689;
  assign n23691 = ~n23684 & n23690;
  assign n23692 = ~n20404 & ~n20484;
  assign n23693 = ~n20554 & ~n20622;
  assign n23694 = n20764 & ~n20837;
  assign n23695 = ~n20838 & ~n20902;
  assign n23696 = ~n20972 & ~n23694;
  assign n23697 = n23695 & n23696;
  assign n23698 = ~n20684 & n23697;
  assign n23699 = ~n21032 & n23698;
  assign n23700 = n23693 & n23699;
  assign n23701 = n23692 & n23700;
  assign n23702 = ~n21168 & ~n21232;
  assign n23703 = n21106 & n23702;
  assign n23704 = n23691 & n23701;
  assign n23705 = ~n23703 & n23704;
  assign n23706 = n23683 & n23705;
  assign n23707 = ~n21370 & n23706;
  assign n23708 = ~n21574 & ~n21614;
  assign n23709 = n21620 & n21632;
  assign n23710 = ~n23708 & ~n23709;
  assign n23711 = ~n21559 & n23710;
  assign n23712 = ~n21434 & n23711;
  assign n23713 = n19763 & n23712;
  assign n23714 = ~n19824 & n23707;
  assign n23715 = ~n21502 & n23714;
  assign n23716 = n23713 & n23715;
  assign n23717 = ~n23686 & ~n23703;
  assign n23718 = ~n21370 & n23717;
  assign n23719 = ~n20267 & n23701;
  assign n23720 = n23683 & n23719;
  assign n23721 = n23718 & n23720;
  assign n23722 = n20040 & ~n20194;
  assign n23723 = ~n21502 & n23722;
  assign n23724 = ~n20116 & n23721;
  assign n23725 = n23712 & n23724;
  assign n23726 = n23723 & n23725;
  assign n23727 = ~n21370 & n23683;
  assign n23728 = ~n19781 & ~n19827;
  assign n23729 = n19659 & n23728;
  assign n23730 = ~n21502 & n23729;
  assign n23731 = ~n19699 & n23705;
  assign n23732 = n23727 & n23731;
  assign n23733 = n23712 & n23732;
  assign n23734 = n23730 & n23733;
  assign n23735 = ~n23716 & ~n23726;
  assign n23736 = ~n23734 & n23735;
  assign n23737 = n20178 & ~n21502;
  assign n23738 = n23701 & ~n23703;
  assign n23739 = ~n20254 & n23738;
  assign n23740 = n23727 & n23739;
  assign n23741 = ~n23686 & n23740;
  assign n23742 = n23712 & n23741;
  assign n23743 = n23737 & n23742;
  assign n23744 = ~n20540 & n23699;
  assign n23745 = ~n23703 & n23727;
  assign n23746 = ~n20622 & n23712;
  assign n23747 = n20462 & ~n21502;
  assign n23748 = n23744 & n23745;
  assign n23749 = n23746 & n23748;
  assign n23750 = n23747 & n23749;
  assign n23751 = ~n20677 & n23695;
  assign n23752 = ~n20972 & ~n23703;
  assign n23753 = ~n21370 & n23752;
  assign n23754 = n23683 & n23753;
  assign n23755 = ~n21032 & n23754;
  assign n23756 = ~n23694 & n23712;
  assign n23757 = n20602 & ~n21502;
  assign n23758 = n23751 & n23755;
  assign n23759 = n23756 & n23758;
  assign n23760 = n23757 & n23759;
  assign n23761 = n20889 & ~n21032;
  assign n23762 = ~n21502 & n23761;
  assign n23763 = n20959 & n23745;
  assign n23764 = n23712 & n23763;
  assign n23765 = n23762 & n23764;
  assign n23766 = ~n23760 & ~n23765;
  assign n23767 = ~n23743 & ~n23750;
  assign n23768 = n23766 & n23767;
  assign n23769 = n20742 & ~n20902;
  assign n23770 = ~n21502 & n23769;
  assign n23771 = ~n20825 & n23755;
  assign n23772 = n23712 & n23771;
  assign n23773 = n23770 & n23772;
  assign n23774 = ~n21031 & ~n21105;
  assign n23775 = n23702 & n23774;
  assign n23776 = ~n21502 & ~n23775;
  assign n23777 = n23712 & n23745;
  assign n23778 = n23776 & n23777;
  assign n23779 = ~n20751 & n23695;
  assign n23780 = n20670 & n23712;
  assign n23781 = n23755 & n23779;
  assign n23782 = ~n21502 & n23781;
  assign n23783 = n23780 & n23782;
  assign n23784 = n21485 & ~n23708;
  assign n23785 = ~n21559 & n23784;
  assign n23786 = n21420 & n23785;
  assign n23787 = ~n23709 & n23786;
  assign n23788 = n21574 & n21614;
  assign n23789 = n21547 & ~n23708;
  assign n23790 = n21483 & n23789;
  assign n23791 = ~n23788 & ~n23790;
  assign n23792 = ~n23709 & ~n23791;
  assign n23793 = n21422 & ~n21559;
  assign n23794 = ~n23708 & n23793;
  assign n23795 = n21353 & n23794;
  assign n23796 = ~n23709 & n23795;
  assign n23797 = ~n21502 & n23796;
  assign n23798 = ~n23787 & ~n23792;
  assign n23799 = ~n23797 & n23798;
  assign n23800 = ~n23773 & ~n23778;
  assign n23801 = ~n23783 & n23800;
  assign n23802 = n23799 & n23801;
  assign n23803 = n19720 & ~n19827;
  assign n23804 = ~n21502 & n23803;
  assign n23805 = ~n19770 & n23707;
  assign n23806 = n23712 & n23805;
  assign n23807 = n23804 & n23806;
  assign n23808 = n19851 & ~n21502;
  assign n23809 = ~n19908 & n23738;
  assign n23810 = n23727 & n23809;
  assign n23811 = n23690 & n23810;
  assign n23812 = n23712 & n23811;
  assign n23813 = n23808 & n23812;
  assign n23814 = ~n19972 & n23712;
  assign n23815 = n19901 & ~n21502;
  assign n23816 = n23689 & n23701;
  assign n23817 = n23745 & n23816;
  assign n23818 = n23814 & n23817;
  assign n23819 = n23815 & n23818;
  assign n23820 = ~n20611 & n23699;
  assign n23821 = n20533 & n23712;
  assign n23822 = n23745 & n23820;
  assign n23823 = ~n21502 & n23822;
  assign n23824 = n23821 & n23823;
  assign n23825 = ~n23819 & ~n23824;
  assign n23826 = n20390 & n23712;
  assign n23827 = ~n20471 & n23700;
  assign n23828 = n23745 & n23827;
  assign n23829 = ~n21502 & n23828;
  assign n23830 = n23826 & n23829;
  assign n23831 = n20818 & n23712;
  assign n23832 = ~n20895 & n23755;
  assign n23833 = ~n21502 & n23832;
  assign n23834 = n23831 & n23833;
  assign n23835 = ~n23830 & ~n23834;
  assign n23836 = ~n20047 & n23685;
  assign n23837 = n19965 & n23712;
  assign n23838 = n23721 & n23836;
  assign n23839 = ~n21502 & n23838;
  assign n23840 = n23837 & n23839;
  assign n23841 = n23835 & ~n23840;
  assign n23842 = ~n23807 & ~n23813;
  assign n23843 = n23825 & n23842;
  assign n23844 = n23841 & n23843;
  assign n23845 = ~n19708 & n23728;
  assign n23846 = ~n19643 & n23845;
  assign n23847 = n19591 & n23712;
  assign n23848 = n23707 & n23846;
  assign n23849 = ~n21502 & n23848;
  assign n23850 = n23847 & n23849;
  assign n23851 = n21299 & ~n21370;
  assign n23852 = ~n21369 & ~n23851;
  assign n23853 = n23712 & ~n23852;
  assign n23854 = ~n21502 & n23853;
  assign n23855 = ~n21620 & ~n21632;
  assign n23856 = ~n21106 & ~n21502;
  assign n23857 = n19483 & ~n19603;
  assign n23858 = ~n19567 & ~n23857;
  assign n23859 = ~n19599 & ~n23858;
  assign n23860 = n19567 & n23857;
  assign n23861 = ~n23684 & ~n23859;
  assign n23862 = ~n19668 & n23861;
  assign n23863 = n23845 & n23862;
  assign n23864 = ~n23860 & n23863;
  assign n23865 = n23701 & n23864;
  assign n23866 = n23727 & n23865;
  assign n23867 = n23690 & n23866;
  assign n23868 = n23712 & n23867;
  assign n23869 = n23856 & n23868;
  assign n23870 = ~n23855 & ~n23869;
  assign n23871 = n20247 & n23712;
  assign n23872 = ~n20320 & n23738;
  assign n23873 = n23727 & n23872;
  assign n23874 = ~n21502 & n23873;
  assign n23875 = n23871 & n23874;
  assign n23876 = n20109 & n23712;
  assign n23877 = ~n20187 & n23721;
  assign n23878 = ~n21502 & n23877;
  assign n23879 = n23876 & n23878;
  assign n23880 = ~n20484 & n23712;
  assign n23881 = n20311 & ~n21502;
  assign n23882 = ~n20397 & n23700;
  assign n23883 = n23745 & n23882;
  assign n23884 = n23880 & n23883;
  assign n23885 = n23881 & n23884;
  assign n23886 = ~n23875 & ~n23879;
  assign n23887 = ~n23885 & n23886;
  assign n23888 = ~n23850 & ~n23854;
  assign n23889 = n23870 & n23888;
  assign n23890 = n23887 & n23889;
  assign n23891 = n23736 & n23768;
  assign n23892 = n23802 & n23891;
  assign n23893 = n23844 & n23892;
  assign n23894 = n23890 & n23893;
  assign n23895 = ~n19573 & ~n23894;
  assign n23896 = n19573 & ~n23615;
  assign n23897 = ~n23895 & ~n23896;
  assign n23898 = n19476 & ~n23897;
  assign n23899 = ~n23680 & ~n23898;
  assign n23900 = n19484 & n23676;
  assign n23901 = n23899 & ~n23900;
  assign n23902 = n19479 & ~n23901;
  assign n23903 = n21764 & n23894;
  assign n23904 = ~n19479 & n23034;
  assign n23905 = n23894 & n23904;
  assign n23906 = n19487 & n19614;
  assign n23907 = n21614 & n23063;
  assign n23908 = ~n21632 & ~n23043;
  assign n23909 = n21547 & n23080;
  assign n23910 = ~n23907 & ~n23908;
  assign n23911 = ~n23909 & n23910;
  assign n23912 = ~n21485 & n23911;
  assign n23913 = ~n23595 & n23912;
  assign n23914 = n21632 & n23043;
  assign n23915 = ~n23913 & ~n23914;
  assign n23916 = n21422 & n23572;
  assign n23917 = ~n21355 & ~n23092;
  assign n23918 = n21222 & n23124;
  assign n23919 = ~n21158 & ~n23144;
  assign n23920 = n21158 & n23144;
  assign n23921 = n21089 & n23156;
  assign n23922 = ~n23920 & ~n23921;
  assign n23923 = ~n20959 & ~n23188;
  assign n23924 = n21025 & n23176;
  assign n23925 = n23923 & ~n23924;
  assign n23926 = ~n20825 & n23222;
  assign n23927 = n20895 & ~n23210;
  assign n23928 = n23926 & ~n23927;
  assign n23929 = n20677 & ~n23256;
  assign n23930 = n20611 & ~n23278;
  assign n23931 = n20540 & ~n23290;
  assign n23932 = ~n20116 & n23392;
  assign n23933 = ~n20047 & n23414;
  assign n23934 = ~n20187 & n23380;
  assign n23935 = ~n20254 & n23358;
  assign n23936 = ~n23932 & ~n23933;
  assign n23937 = ~n23934 & n23936;
  assign n23938 = ~n23935 & n23937;
  assign n23939 = n19972 & ~n23426;
  assign n23940 = n20047 & ~n23414;
  assign n23941 = ~n23939 & ~n23940;
  assign n23942 = ~n19908 & n23448;
  assign n23943 = ~n19972 & n23426;
  assign n23944 = ~n23942 & ~n23943;
  assign n23945 = n19908 & ~n23448;
  assign n23946 = n19824 & ~n23460;
  assign n23947 = ~n23945 & ~n23946;
  assign n23948 = n23944 & ~n23947;
  assign n23949 = n23941 & ~n23948;
  assign n23950 = n23938 & ~n23949;
  assign n23951 = n19770 & ~n23482;
  assign n23952 = ~n19824 & n23460;
  assign n23953 = n23944 & ~n23952;
  assign n23954 = n23938 & n23953;
  assign n23955 = n23951 & n23954;
  assign n23956 = n20254 & ~n23358;
  assign n23957 = ~n23934 & ~n23935;
  assign n23958 = n20187 & ~n23380;
  assign n23959 = n20116 & ~n23392;
  assign n23960 = ~n23958 & ~n23959;
  assign n23961 = n23957 & ~n23960;
  assign n23962 = n20471 & ~n23312;
  assign n23963 = n20397 & ~n23324;
  assign n23964 = ~n23962 & ~n23963;
  assign n23965 = n20320 & ~n23346;
  assign n23966 = n23964 & ~n23965;
  assign n23967 = ~n23956 & ~n23961;
  assign n23968 = n23966 & n23967;
  assign n23969 = n19699 & ~n23494;
  assign n23970 = ~n19770 & n23482;
  assign n23971 = n23954 & ~n23970;
  assign n23972 = n23969 & n23971;
  assign n23973 = ~n19699 & n23494;
  assign n23974 = ~n19643 & n23516;
  assign n23975 = ~n23973 & ~n23974;
  assign n23976 = ~n19567 & n23531;
  assign n23977 = n19643 & ~n23516;
  assign n23978 = n23976 & ~n23977;
  assign n23979 = n23975 & ~n23978;
  assign n23980 = n23971 & n23979;
  assign n23981 = ~n23950 & ~n23955;
  assign n23982 = n23968 & n23981;
  assign n23983 = ~n23972 & n23982;
  assign n23984 = ~n23980 & n23983;
  assign n23985 = ~n20397 & n23324;
  assign n23986 = ~n23962 & n23985;
  assign n23987 = ~n20320 & n23346;
  assign n23988 = n23964 & n23987;
  assign n23989 = ~n20540 & n23290;
  assign n23990 = ~n20471 & n23312;
  assign n23991 = ~n23989 & ~n23990;
  assign n23992 = ~n23986 & ~n23988;
  assign n23993 = n23991 & n23992;
  assign n23994 = ~n23984 & n23993;
  assign n23995 = ~n23931 & ~n23994;
  assign n23996 = ~n20611 & n23278;
  assign n23997 = ~n23995 & ~n23996;
  assign n23998 = ~n23930 & ~n23997;
  assign n23999 = ~n20677 & n23256;
  assign n24000 = ~n23998 & ~n23999;
  assign n24001 = n20825 & ~n23222;
  assign n24002 = ~n23927 & ~n24001;
  assign n24003 = n20751 & ~n23244;
  assign n24004 = n24002 & ~n24003;
  assign n24005 = ~n23929 & ~n24000;
  assign n24006 = n24004 & n24005;
  assign n24007 = ~n20895 & n23210;
  assign n24008 = n20959 & n23188;
  assign n24009 = ~n24007 & ~n24008;
  assign n24010 = ~n20751 & n23244;
  assign n24011 = n24002 & n24010;
  assign n24012 = n24009 & ~n24011;
  assign n24013 = ~n23924 & n24012;
  assign n24014 = ~n23928 & ~n24006;
  assign n24015 = n24013 & n24014;
  assign n24016 = ~n21089 & ~n23156;
  assign n24017 = ~n21025 & ~n23176;
  assign n24018 = ~n24016 & ~n24017;
  assign n24019 = ~n23925 & ~n24015;
  assign n24020 = n24018 & n24019;
  assign n24021 = n23922 & ~n24020;
  assign n24022 = ~n21222 & ~n23124;
  assign n24023 = ~n23919 & ~n24021;
  assign n24024 = ~n24022 & n24023;
  assign n24025 = ~n23918 & ~n24024;
  assign n24026 = n23112 & ~n24025;
  assign n24027 = n21355 & n23092;
  assign n24028 = ~n24026 & ~n24027;
  assign n24029 = ~n23112 & n24025;
  assign n24030 = n21293 & ~n24029;
  assign n24031 = n24028 & ~n24030;
  assign n24032 = ~n21422 & ~n23572;
  assign n24033 = ~n23917 & ~n24031;
  assign n24034 = ~n24032 & n24033;
  assign n24035 = ~n23595 & n23911;
  assign n24036 = ~n23916 & ~n24034;
  assign n24037 = n24035 & n24036;
  assign n24038 = ~n21614 & ~n23063;
  assign n24039 = ~n23908 & n24038;
  assign n24040 = ~n21547 & ~n23907;
  assign n24041 = ~n23908 & n24040;
  assign n24042 = ~n23080 & n24041;
  assign n24043 = ~n24039 & ~n24042;
  assign n24044 = ~n21485 & ~n23916;
  assign n24045 = n23911 & n24044;
  assign n24046 = ~n24034 & n24045;
  assign n24047 = n23915 & ~n24037;
  assign n24048 = n24043 & n24047;
  assign n24049 = ~n24046 & n24048;
  assign n24050 = n23906 & n24049;
  assign n24051 = n19619 & ~n24049;
  assign n24052 = n21743 & ~n23615;
  assign n24053 = ~n23903 & ~n23905;
  assign n24054 = ~n24050 & n24053;
  assign n24055 = ~n24051 & n24054;
  assign n24056 = ~n24052 & n24055;
  assign n24057 = ~n23678 & ~n23902;
  assign n24058 = n24056 & n24057;
  assign n24059 = n22165 & ~n24058;
  assign n3086 = ~n23618 | n24059;
  assign n24061 = n19420 & n19568;
  assign n24062 = ~n19469 & ~n19473;
  assign n24063 = n19552 & n24062;
  assign n24064 = n24061 & ~n24063;
  assign n24065 = n19407 & ~n21744;
  assign n24066 = ~n22158 & n24065;
  assign n24067 = ~n19619 & ~n21764;
  assign n24068 = n19487 & ~n24067;
  assign n24069 = ~n19622 & ~n19627;
  assign n24070 = ~n19625 & n24069;
  assign n24071 = n19483 & ~n24070;
  assign n24072 = ~n19617 & ~n21741;
  assign n24073 = ~n23906 & n24072;
  assign n24074 = ~n19611 & ~n24068;
  assign n24075 = ~n24071 & n24074;
  assign n24076 = n24073 & n24075;
  assign n24077 = ~n24063 & ~n24076;
  assign n24078 = n24066 & ~n24077;
  assign n24079 = P4_STATE_REG & ~n24078;
  assign n24080 = ~n24064 & ~n24079;
  assign n24081 = ~n20529 & ~n24080;
  assign n24082 = n24061 & n24063;
  assign n24083 = n19420 & n21743;
  assign n24084 = ~n24082 & ~n24083;
  assign n24085 = ~n20611 & ~n24084;
  assign n24086 = n19420 & n23026;
  assign n24087 = n19560 & n24063;
  assign n24088 = ~n20602 & n24087;
  assign n24089 = ~n19560 & n24063;
  assign n24090 = ~n20462 & n24089;
  assign n24091 = ~n20529 & ~n24063;
  assign n24092 = ~n24088 & ~n24090;
  assign n24093 = ~n24091 & n24092;
  assign n24094 = n24086 & ~n24093;
  assign n24095 = ~n20462 & ~n22785;
  assign n24096 = ~n20540 & n22775;
  assign n24097 = ~n24095 & ~n24096;
  assign n24098 = ~n20462 & n22775;
  assign n24099 = ~n20540 & ~n22788;
  assign n24100 = ~n24098 & ~n24099;
  assign n24101 = ~n22793 & ~n24100;
  assign n24102 = n22793 & n24100;
  assign n24103 = ~n24101 & ~n24102;
  assign n24104 = ~n24097 & ~n24103;
  assign n24105 = n24097 & n24103;
  assign n24106 = ~n20247 & n22775;
  assign n24107 = ~n20320 & ~n22788;
  assign n24108 = ~n24106 & ~n24107;
  assign n24109 = ~n22793 & ~n24108;
  assign n24110 = n22793 & n24108;
  assign n24111 = ~n24109 & ~n24110;
  assign n24112 = ~n20247 & ~n22785;
  assign n24113 = ~n20320 & n22775;
  assign n24114 = ~n24112 & ~n24113;
  assign n24115 = n24111 & n24114;
  assign n24116 = ~n20311 & n22775;
  assign n24117 = ~n20397 & ~n22788;
  assign n24118 = ~n24116 & ~n24117;
  assign n24119 = ~n22793 & ~n24118;
  assign n24120 = n22793 & n24118;
  assign n24121 = ~n24119 & ~n24120;
  assign n24122 = ~n20311 & ~n22785;
  assign n24123 = ~n20397 & n22775;
  assign n24124 = ~n24122 & ~n24123;
  assign n24125 = n24121 & n24124;
  assign n24126 = ~n20390 & n22775;
  assign n24127 = ~n20471 & ~n22788;
  assign n24128 = ~n24126 & ~n24127;
  assign n24129 = ~n22793 & ~n24128;
  assign n24130 = n22793 & n24128;
  assign n24131 = ~n24129 & ~n24130;
  assign n24132 = ~n20390 & ~n22785;
  assign n24133 = ~n20471 & n22775;
  assign n24134 = ~n24132 & ~n24133;
  assign n24135 = n24131 & n24134;
  assign n24136 = ~n24125 & ~n24135;
  assign n24137 = ~n24115 & n24136;
  assign n24138 = ~n20178 & ~n22785;
  assign n24139 = ~n20254 & n22775;
  assign n24140 = ~n24138 & ~n24139;
  assign n24141 = ~n20178 & n22775;
  assign n24142 = ~n20254 & ~n22788;
  assign n24143 = ~n24141 & ~n24142;
  assign n24144 = ~n22793 & ~n24143;
  assign n24145 = n22793 & n24143;
  assign n24146 = ~n24144 & ~n24145;
  assign n24147 = ~n24140 & ~n24146;
  assign n24148 = n24140 & n24146;
  assign n24149 = ~n20109 & n22775;
  assign n24150 = ~n20187 & ~n22788;
  assign n24151 = ~n24149 & ~n24150;
  assign n24152 = ~n22793 & ~n24151;
  assign n24153 = n22793 & n24151;
  assign n24154 = ~n24152 & ~n24153;
  assign n24155 = ~n20109 & ~n22785;
  assign n24156 = ~n20187 & n22775;
  assign n24157 = ~n24155 & ~n24156;
  assign n24158 = n24154 & n24157;
  assign n24159 = ~n20040 & ~n22785;
  assign n24160 = ~n20116 & n22775;
  assign n24161 = ~n24159 & ~n24160;
  assign n24162 = ~n20040 & n22775;
  assign n24163 = ~n20116 & ~n22788;
  assign n24164 = ~n24162 & ~n24163;
  assign n24165 = ~n22793 & ~n24164;
  assign n24166 = n22793 & n24164;
  assign n24167 = ~n24165 & ~n24166;
  assign n24168 = ~n24161 & ~n24167;
  assign n24169 = n24161 & n24167;
  assign n24170 = ~n19851 & ~n22785;
  assign n24171 = ~n19908 & n22775;
  assign n24172 = ~n24170 & ~n24171;
  assign n24173 = ~n19851 & n22775;
  assign n24174 = ~n19908 & ~n22788;
  assign n24175 = ~n24173 & ~n24174;
  assign n24176 = ~n22793 & ~n24175;
  assign n24177 = n22793 & n24175;
  assign n24178 = ~n24176 & ~n24177;
  assign n24179 = ~n24172 & ~n24178;
  assign n24180 = ~n19901 & n22775;
  assign n24181 = ~n19972 & ~n22788;
  assign n24182 = ~n24180 & ~n24181;
  assign n24183 = ~n22793 & ~n24182;
  assign n24184 = n22793 & n24182;
  assign n24185 = ~n24183 & ~n24184;
  assign n24186 = ~n19901 & ~n22785;
  assign n24187 = ~n19972 & n22775;
  assign n24188 = ~n24186 & ~n24187;
  assign n24189 = n24185 & n24188;
  assign n24190 = ~n19965 & n22775;
  assign n24191 = ~n20047 & ~n22788;
  assign n24192 = ~n24190 & ~n24191;
  assign n24193 = ~n22793 & ~n24192;
  assign n24194 = n22793 & n24192;
  assign n24195 = ~n24193 & ~n24194;
  assign n24196 = ~n19965 & ~n22785;
  assign n24197 = ~n20047 & n22775;
  assign n24198 = ~n24196 & ~n24197;
  assign n24199 = n24195 & n24198;
  assign n24200 = ~n24189 & ~n24199;
  assign n24201 = n24179 & n24200;
  assign n24202 = ~n24185 & ~n24188;
  assign n24203 = ~n24198 & n24202;
  assign n24204 = n24195 & ~n24203;
  assign n24205 = n24198 & ~n24202;
  assign n24206 = ~n24204 & ~n24205;
  assign n24207 = ~n24201 & ~n24206;
  assign n24208 = n24172 & n24178;
  assign n24209 = n24200 & ~n24208;
  assign n24210 = ~n19763 & n22775;
  assign n24211 = ~n19824 & ~n22788;
  assign n24212 = ~n24210 & ~n24211;
  assign n24213 = ~n22793 & ~n24212;
  assign n24214 = n22793 & n24212;
  assign n24215 = ~n24213 & ~n24214;
  assign n24216 = ~n19763 & ~n22785;
  assign n24217 = ~n19824 & n22775;
  assign n24218 = ~n24216 & ~n24217;
  assign n24219 = n24215 & n24218;
  assign n24220 = ~n19720 & ~n22785;
  assign n24221 = ~n19770 & n22775;
  assign n24222 = ~n24220 & ~n24221;
  assign n24223 = ~n19659 & ~n22785;
  assign n24224 = ~n19699 & n22775;
  assign n24225 = ~n24223 & ~n24224;
  assign n24226 = ~n19659 & n22775;
  assign n24227 = n22788 & ~n24226;
  assign n24228 = n19699 & ~n24226;
  assign n24229 = ~n24227 & ~n24228;
  assign n24230 = ~n22793 & n24229;
  assign n24231 = n22793 & ~n24229;
  assign n24232 = ~n24230 & ~n24231;
  assign n24233 = ~n24225 & ~n24232;
  assign n24234 = ~n24222 & n24233;
  assign n24235 = ~n19720 & n22775;
  assign n24236 = n22788 & ~n24235;
  assign n24237 = n19770 & ~n24235;
  assign n24238 = ~n24236 & ~n24237;
  assign n24239 = ~n22793 & n24238;
  assign n24240 = n22793 & ~n24238;
  assign n24241 = ~n24239 & ~n24240;
  assign n24242 = n24222 & ~n24233;
  assign n24243 = ~n24241 & ~n24242;
  assign n24244 = ~n24234 & ~n24243;
  assign n24245 = n24225 & n24232;
  assign n24246 = n24222 & n24241;
  assign n24247 = ~n24245 & ~n24246;
  assign n24248 = n22793 & ~n22804;
  assign n24249 = ~n19591 & n22775;
  assign n24250 = ~n19643 & ~n22788;
  assign n24251 = ~n24249 & ~n24250;
  assign n24252 = ~n22793 & ~n24251;
  assign n24253 = n22793 & n24251;
  assign n24254 = ~n24252 & ~n24253;
  assign n24255 = ~n19591 & ~n22785;
  assign n24256 = ~n19643 & n22775;
  assign n24257 = ~n24255 & ~n24256;
  assign n24258 = n24254 & n24257;
  assign n24259 = n24248 & ~n24258;
  assign n24260 = ~n24254 & ~n24257;
  assign n24261 = ~n22793 & n22804;
  assign n24262 = ~n22796 & ~n24258;
  assign n24263 = ~n24261 & n24262;
  assign n24264 = ~n24259 & ~n24260;
  assign n24265 = ~n24263 & n24264;
  assign n24266 = n24247 & ~n24265;
  assign n24267 = n24244 & ~n24266;
  assign n24268 = ~n24219 & ~n24267;
  assign n24269 = ~n24215 & ~n24218;
  assign n24270 = ~n24268 & ~n24269;
  assign n24271 = n24209 & ~n24270;
  assign n24272 = n24207 & ~n24271;
  assign n24273 = ~n24169 & ~n24272;
  assign n24274 = ~n24168 & ~n24273;
  assign n24275 = ~n24158 & ~n24274;
  assign n24276 = ~n24154 & ~n24157;
  assign n24277 = ~n24275 & ~n24276;
  assign n24278 = ~n24148 & ~n24277;
  assign n24279 = ~n24147 & ~n24278;
  assign n24280 = n24137 & ~n24279;
  assign n24281 = ~n24131 & ~n24134;
  assign n24282 = ~n24121 & ~n24124;
  assign n24283 = ~n24281 & ~n24282;
  assign n24284 = ~n24111 & ~n24114;
  assign n24285 = n24136 & n24284;
  assign n24286 = n24283 & ~n24285;
  assign n24287 = ~n24135 & ~n24286;
  assign n24288 = ~n24280 & ~n24287;
  assign n24289 = ~n24105 & ~n24288;
  assign n24290 = ~n24104 & ~n24289;
  assign n24291 = ~n20533 & n22775;
  assign n24292 = ~n20611 & ~n22788;
  assign n24293 = ~n24291 & ~n24292;
  assign n24294 = ~n22793 & ~n24293;
  assign n24295 = n22793 & n24293;
  assign n24296 = ~n24294 & ~n24295;
  assign n24297 = ~n20533 & ~n22785;
  assign n24298 = ~n20611 & n22775;
  assign n24299 = ~n24297 & ~n24298;
  assign n24300 = ~n24296 & n24299;
  assign n24301 = n24296 & ~n24299;
  assign n24302 = ~n24300 & ~n24301;
  assign n24303 = n24290 & ~n24302;
  assign n24304 = ~n24290 & n24302;
  assign n24305 = ~n24303 & ~n24304;
  assign n24306 = n19420 & ~n24076;
  assign n24307 = n24063 & n24306;
  assign n24308 = ~n24305 & n24307;
  assign n24309 = ~n24081 & ~n24085;
  assign n24310 = ~n22458 & n24309;
  assign n24311 = ~n24094 & n24310;
  assign n3091 = n24308 | ~n24311;
  assign n24313 = n19568 & ~n24063;
  assign n24314 = n24078 & ~n24313;
  assign n24315 = P4_STATE_REG & ~n24314;
  assign n24316 = ~n21285 & n24315;
  assign n24317 = n19568 & n24063;
  assign n24318 = ~n21743 & ~n24317;
  assign n24319 = n19420 & ~n24318;
  assign n24320 = n21355 & n24319;
  assign n24321 = P4_REG3_REG_26_ & ~P4_STATE_REG;
  assign n24322 = ~n21285 & ~n24063;
  assign n24323 = ~n21220 & n24089;
  assign n24324 = ~n21353 & n24087;
  assign n24325 = ~n24322 & ~n24323;
  assign n24326 = ~n24324 & n24325;
  assign n24327 = n24086 & ~n24326;
  assign n24328 = ~n21220 & n22775;
  assign n24329 = n21293 & ~n22788;
  assign n24330 = ~n24328 & ~n24329;
  assign n24331 = ~n22793 & ~n24330;
  assign n24332 = n22793 & n24330;
  assign n24333 = ~n24331 & ~n24332;
  assign n24334 = ~n21220 & ~n22785;
  assign n24335 = n21293 & n22775;
  assign n24336 = ~n24334 & ~n24335;
  assign n24337 = n24333 & n24336;
  assign n24338 = ~n21289 & n22775;
  assign n24339 = n21355 & ~n22788;
  assign n24340 = ~n24338 & ~n24339;
  assign n24341 = ~n22793 & ~n24340;
  assign n24342 = n22793 & n24340;
  assign n24343 = ~n24341 & ~n24342;
  assign n24344 = ~n21289 & ~n22785;
  assign n24345 = n21355 & n22775;
  assign n24346 = ~n24344 & ~n24345;
  assign n24347 = n24343 & n24346;
  assign n24348 = ~n24343 & ~n24346;
  assign n24349 = ~n24337 & ~n24347;
  assign n24350 = ~n24348 & n24349;
  assign n24351 = ~n21154 & n22775;
  assign n24352 = n21222 & ~n22788;
  assign n24353 = ~n24351 & ~n24352;
  assign n24354 = ~n22793 & ~n24353;
  assign n24355 = n22793 & n24353;
  assign n24356 = ~n24354 & ~n24355;
  assign n24357 = ~n21154 & ~n22785;
  assign n24358 = n21222 & n22775;
  assign n24359 = ~n24357 & ~n24358;
  assign n24360 = n24356 & n24359;
  assign n24361 = ~n21087 & ~n22785;
  assign n24362 = n21158 & n22775;
  assign n24363 = ~n24361 & ~n24362;
  assign n24364 = ~n21087 & n22775;
  assign n24365 = n21158 & ~n22788;
  assign n24366 = ~n24364 & ~n24365;
  assign n24367 = ~n22793 & ~n24366;
  assign n24368 = n22793 & n24366;
  assign n24369 = ~n24367 & ~n24368;
  assign n24370 = ~n24363 & ~n24369;
  assign n24371 = n24363 & n24369;
  assign n24372 = ~n21021 & ~n22785;
  assign n24373 = n21089 & n22775;
  assign n24374 = ~n24372 & ~n24373;
  assign n24375 = ~n21021 & n22775;
  assign n24376 = n21089 & ~n22788;
  assign n24377 = ~n24375 & ~n24376;
  assign n24378 = ~n22793 & ~n24377;
  assign n24379 = n22793 & n24377;
  assign n24380 = ~n24378 & ~n24379;
  assign n24381 = ~n24374 & ~n24380;
  assign n24382 = n24374 & n24380;
  assign n24383 = ~n20818 & n22775;
  assign n24384 = ~n20895 & ~n22788;
  assign n24385 = ~n24383 & ~n24384;
  assign n24386 = ~n22793 & ~n24385;
  assign n24387 = n22793 & n24385;
  assign n24388 = ~n24386 & ~n24387;
  assign n24389 = ~n20818 & ~n22785;
  assign n24390 = ~n20895 & n22775;
  assign n24391 = ~n24389 & ~n24390;
  assign n24392 = n24388 & n24391;
  assign n24393 = ~n20889 & n22775;
  assign n24394 = n20959 & ~n22788;
  assign n24395 = ~n24393 & ~n24394;
  assign n24396 = ~n22793 & ~n24395;
  assign n24397 = n22793 & n24395;
  assign n24398 = ~n24396 & ~n24397;
  assign n24399 = ~n20889 & ~n22785;
  assign n24400 = n20959 & n22775;
  assign n24401 = ~n24399 & ~n24400;
  assign n24402 = n24398 & n24401;
  assign n24403 = ~n20957 & n22775;
  assign n24404 = n21025 & ~n22788;
  assign n24405 = ~n24403 & ~n24404;
  assign n24406 = ~n22793 & ~n24405;
  assign n24407 = n22793 & n24405;
  assign n24408 = ~n24406 & ~n24407;
  assign n24409 = ~n20957 & ~n22785;
  assign n24410 = n21025 & n22775;
  assign n24411 = ~n24409 & ~n24410;
  assign n24412 = n24408 & n24411;
  assign n24413 = ~n24402 & ~n24412;
  assign n24414 = ~n24392 & n24413;
  assign n24415 = ~n20742 & ~n22785;
  assign n24416 = ~n20825 & n22775;
  assign n24417 = ~n24415 & ~n24416;
  assign n24418 = ~n20742 & n22775;
  assign n24419 = ~n20825 & ~n22788;
  assign n24420 = ~n24418 & ~n24419;
  assign n24421 = ~n22793 & ~n24420;
  assign n24422 = n22793 & n24420;
  assign n24423 = ~n24421 & ~n24422;
  assign n24424 = ~n24417 & ~n24423;
  assign n24425 = n24417 & n24423;
  assign n24426 = ~n20670 & ~n22785;
  assign n24427 = ~n20751 & n22775;
  assign n24428 = ~n24426 & ~n24427;
  assign n24429 = ~n20602 & ~n22785;
  assign n24430 = ~n20677 & n22775;
  assign n24431 = ~n24429 & ~n24430;
  assign n24432 = ~n20602 & n22775;
  assign n24433 = ~n20677 & ~n22788;
  assign n24434 = ~n24432 & ~n24433;
  assign n24435 = ~n22793 & ~n24434;
  assign n24436 = n22793 & n24434;
  assign n24437 = ~n24435 & ~n24436;
  assign n24438 = ~n24431 & ~n24437;
  assign n24439 = ~n24428 & n24438;
  assign n24440 = ~n20670 & n22775;
  assign n24441 = ~n20751 & ~n22788;
  assign n24442 = ~n24440 & ~n24441;
  assign n24443 = ~n22793 & ~n24442;
  assign n24444 = n22793 & n24442;
  assign n24445 = ~n24443 & ~n24444;
  assign n24446 = n24428 & ~n24438;
  assign n24447 = ~n24445 & ~n24446;
  assign n24448 = ~n24439 & ~n24447;
  assign n24449 = n24431 & n24437;
  assign n24450 = n24428 & n24445;
  assign n24451 = ~n24449 & ~n24450;
  assign n24452 = ~n24296 & ~n24299;
  assign n24453 = n24296 & n24299;
  assign n24454 = ~n24290 & ~n24453;
  assign n24455 = ~n24452 & ~n24454;
  assign n24456 = n24451 & ~n24455;
  assign n24457 = n24448 & ~n24456;
  assign n24458 = ~n24425 & ~n24457;
  assign n24459 = ~n24424 & ~n24458;
  assign n24460 = n24414 & ~n24459;
  assign n24461 = ~n24408 & ~n24411;
  assign n24462 = ~n24398 & ~n24401;
  assign n24463 = ~n24461 & ~n24462;
  assign n24464 = ~n24388 & ~n24391;
  assign n24465 = n24413 & n24464;
  assign n24466 = n24463 & ~n24465;
  assign n24467 = ~n24412 & ~n24466;
  assign n24468 = ~n24460 & ~n24467;
  assign n24469 = ~n24382 & ~n24468;
  assign n24470 = ~n24381 & ~n24469;
  assign n24471 = ~n24371 & ~n24470;
  assign n24472 = ~n24370 & ~n24471;
  assign n24473 = ~n24360 & ~n24472;
  assign n24474 = n24350 & n24473;
  assign n24475 = ~n24356 & ~n24359;
  assign n24476 = ~n24333 & ~n24336;
  assign n24477 = ~n24475 & ~n24476;
  assign n24478 = ~n24343 & n24346;
  assign n24479 = n24343 & ~n24346;
  assign n24480 = ~n24478 & ~n24479;
  assign n24481 = n24477 & n24480;
  assign n24482 = ~n24473 & n24481;
  assign n24483 = ~n24347 & n24476;
  assign n24484 = ~n24348 & n24483;
  assign n24485 = n24337 & n24480;
  assign n24486 = ~n24348 & n24475;
  assign n24487 = ~n24337 & n24486;
  assign n24488 = ~n24347 & n24487;
  assign n24489 = ~n24484 & ~n24485;
  assign n24490 = ~n24488 & n24489;
  assign n24491 = ~n24474 & ~n24482;
  assign n24492 = n24490 & n24491;
  assign n24493 = n24307 & n24492;
  assign n24494 = ~n24316 & ~n24320;
  assign n24495 = ~n24321 & n24494;
  assign n24496 = ~n24327 & n24495;
  assign n3096 = n24493 | ~n24496;
  assign n24498 = ~n19894 & ~n24080;
  assign n24499 = ~n19972 & ~n24084;
  assign n24500 = ~n24185 & n24188;
  assign n24501 = n24185 & ~n24188;
  assign n24502 = ~n24500 & ~n24501;
  assign n24503 = ~n24208 & ~n24270;
  assign n24504 = ~n24179 & ~n24503;
  assign n24505 = ~n24502 & n24504;
  assign n24506 = ~n24189 & ~n24202;
  assign n24507 = ~n24504 & ~n24506;
  assign n24508 = ~n24505 & ~n24507;
  assign n24509 = n24307 & ~n24508;
  assign n24510 = ~n22699 & ~n24509;
  assign n24511 = ~n19965 & n24087;
  assign n24512 = ~n19851 & n24089;
  assign n24513 = ~n19894 & ~n24063;
  assign n24514 = ~n24511 & ~n24512;
  assign n24515 = ~n24513 & n24514;
  assign n24516 = n24086 & ~n24515;
  assign n24517 = ~n24498 & ~n24499;
  assign n24518 = n24510 & n24517;
  assign n3101 = n24516 | ~n24518;
  assign n24520 = ~n20738 & ~n24080;
  assign n24521 = ~n20825 & ~n24084;
  assign n24522 = ~n20818 & n24087;
  assign n24523 = ~n20670 & n24089;
  assign n24524 = ~n20738 & ~n24063;
  assign n24525 = ~n24522 & ~n24523;
  assign n24526 = ~n24524 & n24525;
  assign n24527 = n24086 & ~n24526;
  assign n24528 = n24417 & ~n24423;
  assign n24529 = ~n24417 & n24423;
  assign n24530 = ~n24528 & ~n24529;
  assign n24531 = n24457 & ~n24530;
  assign n24532 = ~n24457 & n24530;
  assign n24533 = ~n24531 & ~n24532;
  assign n24534 = n24307 & ~n24533;
  assign n24535 = ~n24520 & ~n24521;
  assign n24536 = ~n22385 & n24535;
  assign n24537 = ~n24527 & n24536;
  assign n3106 = n24534 | ~n24537;
  assign n24539 = n24225 & ~n24232;
  assign n24540 = ~n24225 & n24232;
  assign n24541 = ~n24539 & ~n24540;
  assign n24542 = n24265 & ~n24541;
  assign n24543 = ~n24233 & ~n24245;
  assign n24544 = ~n24265 & ~n24543;
  assign n24545 = ~n24542 & ~n24544;
  assign n24546 = n24307 & ~n24545;
  assign n24547 = ~n22855 & ~n24546;
  assign n24548 = ~n19699 & ~n24084;
  assign n24549 = n24547 & ~n24548;
  assign n24550 = P4_REG3_REG_2_ & ~n24080;
  assign n24551 = ~n19720 & n24087;
  assign n24552 = ~n19591 & n24089;
  assign n24553 = P4_REG3_REG_2_ & ~n24063;
  assign n24554 = ~n24551 & ~n24552;
  assign n24555 = ~n24553 & n24554;
  assign n24556 = n24086 & ~n24555;
  assign n24557 = n24549 & ~n24550;
  assign n3111 = n24556 | ~n24557;
  assign n24559 = ~n20240 & ~n24080;
  assign n24560 = ~n20320 & ~n24084;
  assign n24561 = ~n20311 & n24087;
  assign n24562 = ~n20178 & n24089;
  assign n24563 = ~n20240 & ~n24063;
  assign n24564 = ~n24561 & ~n24562;
  assign n24565 = ~n24563 & n24564;
  assign n24566 = n24086 & ~n24565;
  assign n24567 = ~n24111 & n24114;
  assign n24568 = n24111 & ~n24114;
  assign n24569 = ~n24567 & ~n24568;
  assign n24570 = n24279 & ~n24569;
  assign n24571 = ~n24115 & ~n24284;
  assign n24572 = ~n24279 & ~n24571;
  assign n24573 = ~n24570 & ~n24572;
  assign n24574 = n24307 & ~n24573;
  assign n24575 = ~n24559 & ~n24560;
  assign n24576 = ~n22561 & n24575;
  assign n24577 = ~n24566 & n24576;
  assign n3116 = n24574 | ~n24577;
  assign n24579 = ~n21017 & n24315;
  assign n24580 = n21089 & n24319;
  assign n24581 = P4_REG3_REG_22_ & ~P4_STATE_REG;
  assign n24582 = ~n21087 & n24087;
  assign n24583 = ~n20957 & n24089;
  assign n24584 = ~n21017 & ~n24063;
  assign n24585 = ~n24582 & ~n24583;
  assign n24586 = ~n24584 & n24585;
  assign n24587 = n24086 & ~n24586;
  assign n24588 = n24374 & ~n24380;
  assign n24589 = ~n24374 & n24380;
  assign n24590 = ~n24588 & ~n24589;
  assign n24591 = n24468 & ~n24590;
  assign n24592 = ~n24468 & n24590;
  assign n24593 = ~n24591 & ~n24592;
  assign n24594 = n24307 & ~n24593;
  assign n24595 = ~n24579 & ~n24580;
  assign n24596 = ~n24581 & n24595;
  assign n24597 = ~n24587 & n24596;
  assign n3121 = n24594 | ~n24597;
  assign n24599 = ~n20386 & ~n24080;
  assign n24600 = ~n20471 & ~n24084;
  assign n24601 = ~n20462 & n24087;
  assign n24602 = ~n20311 & n24089;
  assign n24603 = ~n20386 & ~n24063;
  assign n24604 = ~n24601 & ~n24602;
  assign n24605 = ~n24603 & n24604;
  assign n24606 = n24086 & ~n24605;
  assign n24607 = n24136 & ~n24281;
  assign n24608 = ~n24115 & ~n24279;
  assign n24609 = ~n24284 & ~n24608;
  assign n24610 = ~n24282 & n24609;
  assign n24611 = n24607 & ~n24610;
  assign n24612 = ~n24131 & n24134;
  assign n24613 = n24131 & ~n24134;
  assign n24614 = ~n24612 & ~n24613;
  assign n24615 = ~n24282 & n24614;
  assign n24616 = ~n24125 & ~n24609;
  assign n24617 = n24615 & ~n24616;
  assign n24618 = ~n24611 & ~n24617;
  assign n24619 = n24307 & n24618;
  assign n24620 = ~n24599 & ~n24600;
  assign n24621 = ~n22510 & n24620;
  assign n24622 = ~n24606 & n24621;
  assign n3126 = n24619 | ~n24622;
  assign n24624 = ~n20885 & n24315;
  assign n24625 = n20959 & n24319;
  assign n24626 = P4_REG3_REG_20_ & ~P4_STATE_REG;
  assign n24627 = ~n20957 & n24087;
  assign n24628 = ~n20818 & n24089;
  assign n24629 = ~n20885 & ~n24063;
  assign n24630 = ~n24627 & ~n24628;
  assign n24631 = ~n24629 & n24630;
  assign n24632 = n24086 & ~n24631;
  assign n24633 = ~n24398 & n24401;
  assign n24634 = n24398 & ~n24401;
  assign n24635 = ~n24633 & ~n24634;
  assign n24636 = ~n24392 & ~n24459;
  assign n24637 = ~n24464 & ~n24636;
  assign n24638 = ~n24635 & n24637;
  assign n24639 = ~n24402 & ~n24462;
  assign n24640 = ~n24637 & ~n24639;
  assign n24641 = ~n24638 & ~n24640;
  assign n24642 = n24307 & ~n24641;
  assign n24643 = ~n24624 & ~n24625;
  assign n24644 = ~n24626 & n24643;
  assign n24645 = ~n24632 & n24644;
  assign n3131 = n24642 | ~n24645;
  assign n24647 = ~n22807 & n24307;
  assign n24648 = ~n22913 & ~n24647;
  assign n24649 = ~n24061 & ~n24086;
  assign n24650 = ~n24063 & ~n24649;
  assign n24651 = ~n24079 & ~n24650;
  assign n24652 = P4_REG3_REG_0_ & ~n24651;
  assign n24653 = ~n19567 & ~n24084;
  assign n24654 = ~n19591 & n24086;
  assign n24655 = n24087 & n24654;
  assign n24656 = ~n24653 & ~n24655;
  assign n24657 = n24648 & ~n24652;
  assign n3136 = ~n24656 | ~n24657;
  assign n24659 = ~n20102 & ~n24080;
  assign n24660 = ~n20187 & ~n24084;
  assign n24661 = ~n20178 & n24087;
  assign n24662 = ~n20040 & n24089;
  assign n24663 = ~n20102 & ~n24063;
  assign n24664 = ~n24661 & ~n24662;
  assign n24665 = ~n24663 & n24664;
  assign n24666 = n24086 & ~n24665;
  assign n24667 = ~n24154 & n24157;
  assign n24668 = n24154 & ~n24157;
  assign n24669 = ~n24667 & ~n24668;
  assign n24670 = n24274 & ~n24669;
  assign n24671 = ~n24274 & n24669;
  assign n24672 = ~n24670 & ~n24671;
  assign n24673 = n24307 & ~n24672;
  assign n24674 = ~n24659 & ~n24660;
  assign n24675 = ~n22615 & n24674;
  assign n24676 = ~n24666 & n24675;
  assign n3141 = n24673 | ~n24676;
  assign n24678 = ~n24215 & n24218;
  assign n24679 = n24215 & ~n24218;
  assign n24680 = ~n24678 & ~n24679;
  assign n24681 = n24267 & ~n24680;
  assign n24682 = ~n24267 & n24680;
  assign n24683 = ~n24681 & ~n24682;
  assign n24684 = n24307 & ~n24683;
  assign n24685 = ~n22755 & ~n24684;
  assign n24686 = ~n19824 & ~n24084;
  assign n24687 = n24685 & ~n24686;
  assign n24688 = ~n19756 & ~n24080;
  assign n24689 = ~n19851 & n24087;
  assign n24690 = ~n19720 & n24089;
  assign n24691 = ~n19756 & ~n24063;
  assign n24692 = ~n24689 & ~n24690;
  assign n24693 = ~n24691 & n24692;
  assign n24694 = n24086 & ~n24693;
  assign n24695 = n24687 & ~n24688;
  assign n3146 = n24694 | ~n24695;
  assign n24697 = ~n21150 & n24315;
  assign n24698 = n21222 & n24319;
  assign n24699 = P4_REG3_REG_24_ & ~P4_STATE_REG;
  assign n24700 = ~n21220 & n24087;
  assign n24701 = ~n21087 & n24089;
  assign n24702 = ~n21150 & ~n24063;
  assign n24703 = ~n24700 & ~n24701;
  assign n24704 = ~n24702 & n24703;
  assign n24705 = n24086 & ~n24704;
  assign n24706 = ~n24356 & n24359;
  assign n24707 = n24356 & ~n24359;
  assign n24708 = ~n24706 & ~n24707;
  assign n24709 = n24472 & ~n24708;
  assign n24710 = ~n24360 & ~n24475;
  assign n24711 = ~n24472 & ~n24710;
  assign n24712 = ~n24709 & ~n24711;
  assign n24713 = n24307 & ~n24712;
  assign n24714 = ~n24697 & ~n24698;
  assign n24715 = ~n24699 & n24714;
  assign n24716 = ~n24705 & n24715;
  assign n3151 = n24713 | ~n24716;
  assign n24718 = ~n20666 & ~n24080;
  assign n24719 = ~n20751 & ~n24084;
  assign n24720 = ~n20742 & n24087;
  assign n24721 = ~n20602 & n24089;
  assign n24722 = ~n20666 & ~n24063;
  assign n24723 = ~n24720 & ~n24721;
  assign n24724 = ~n24722 & n24723;
  assign n24725 = n24086 & ~n24724;
  assign n24726 = ~n24428 & ~n24445;
  assign n24727 = n24451 & ~n24726;
  assign n24728 = ~n24438 & n24455;
  assign n24729 = n24727 & ~n24728;
  assign n24730 = n24428 & ~n24445;
  assign n24731 = ~n24428 & n24445;
  assign n24732 = ~n24730 & ~n24731;
  assign n24733 = ~n24438 & n24732;
  assign n24734 = ~n24449 & ~n24455;
  assign n24735 = n24733 & ~n24734;
  assign n24736 = ~n24729 & ~n24735;
  assign n24737 = n24307 & n24736;
  assign n24738 = ~n24718 & ~n24719;
  assign n24739 = ~n22413 & n24738;
  assign n24740 = ~n24725 & n24739;
  assign n3156 = n24737 | ~n24740;
  assign n24742 = n24172 & ~n24178;
  assign n24743 = ~n24172 & n24178;
  assign n24744 = ~n24742 & ~n24743;
  assign n24745 = n24270 & ~n24744;
  assign n24746 = ~n24270 & n24744;
  assign n24747 = ~n24745 & ~n24746;
  assign n24748 = n24307 & ~n24747;
  assign n24749 = ~n22725 & ~n24748;
  assign n24750 = ~n19908 & ~n24084;
  assign n24751 = n24749 & ~n24750;
  assign n24752 = ~n19844 & ~n24080;
  assign n24753 = ~n19901 & n24087;
  assign n24754 = ~n19763 & n24089;
  assign n24755 = ~n19844 & ~n24063;
  assign n24756 = ~n24753 & ~n24754;
  assign n24757 = ~n24755 & n24756;
  assign n24758 = n24086 & ~n24757;
  assign n24759 = n24751 & ~n24752;
  assign n3161 = n24758 | ~n24759;
  assign n24761 = ~n20598 & ~n24080;
  assign n24762 = ~n20677 & ~n24084;
  assign n24763 = ~n20670 & n24087;
  assign n24764 = ~n20533 & n24089;
  assign n24765 = ~n20598 & ~n24063;
  assign n24766 = ~n24763 & ~n24764;
  assign n24767 = ~n24765 & n24766;
  assign n24768 = n24086 & ~n24767;
  assign n24769 = n24431 & ~n24437;
  assign n24770 = ~n24431 & n24437;
  assign n24771 = ~n24769 & ~n24770;
  assign n24772 = n24455 & ~n24771;
  assign n24773 = ~n24438 & ~n24449;
  assign n24774 = ~n24455 & ~n24773;
  assign n24775 = ~n24772 & ~n24774;
  assign n24776 = n24307 & ~n24775;
  assign n24777 = ~n24761 & ~n24762;
  assign n24778 = ~n22441 & n24777;
  assign n24779 = ~n24768 & n24778;
  assign n3166 = n24776 | ~n24779;
  assign n24781 = ~n21216 & n24315;
  assign n24782 = n21293 & n24319;
  assign n24783 = P4_REG3_REG_25_ & ~P4_STATE_REG;
  assign n24784 = ~n21289 & n24087;
  assign n24785 = ~n21154 & n24089;
  assign n24786 = ~n21216 & ~n24063;
  assign n24787 = ~n24784 & ~n24785;
  assign n24788 = ~n24786 & n24787;
  assign n24789 = n24086 & ~n24788;
  assign n24790 = ~n24473 & ~n24475;
  assign n24791 = ~n24333 & n24336;
  assign n24792 = n24333 & ~n24336;
  assign n24793 = ~n24791 & ~n24792;
  assign n24794 = n24790 & ~n24793;
  assign n24795 = ~n24337 & ~n24476;
  assign n24796 = ~n24790 & ~n24795;
  assign n24797 = ~n24794 & ~n24796;
  assign n24798 = n24307 & ~n24797;
  assign n24799 = ~n24781 & ~n24782;
  assign n24800 = ~n24783 & n24799;
  assign n24801 = ~n24789 & n24800;
  assign n3171 = n24798 | ~n24801;
  assign n24803 = ~n20304 & ~n24080;
  assign n24804 = ~n20397 & ~n24084;
  assign n24805 = ~n20390 & n24087;
  assign n24806 = ~n20247 & n24089;
  assign n24807 = ~n20304 & ~n24063;
  assign n24808 = ~n24805 & ~n24806;
  assign n24809 = ~n24807 & n24808;
  assign n24810 = n24086 & ~n24809;
  assign n24811 = ~n24121 & n24124;
  assign n24812 = n24121 & ~n24124;
  assign n24813 = ~n24811 & ~n24812;
  assign n24814 = n24609 & ~n24813;
  assign n24815 = ~n24125 & ~n24282;
  assign n24816 = ~n24609 & ~n24815;
  assign n24817 = ~n24814 & ~n24816;
  assign n24818 = n24307 & ~n24817;
  assign n24819 = ~n24803 & ~n24804;
  assign n24820 = ~n22533 & n24819;
  assign n24821 = ~n24810 & n24820;
  assign n3176 = n24818 | ~n24821;
  assign n24823 = ~n20953 & n24315;
  assign n24824 = n21025 & n24319;
  assign n24825 = P4_REG3_REG_21_ & ~P4_STATE_REG;
  assign n24826 = ~n21021 & n24087;
  assign n24827 = ~n20889 & n24089;
  assign n24828 = ~n20953 & ~n24063;
  assign n24829 = ~n24826 & ~n24827;
  assign n24830 = ~n24828 & n24829;
  assign n24831 = n24086 & ~n24830;
  assign n24832 = n24413 & ~n24461;
  assign n24833 = ~n24462 & n24637;
  assign n24834 = n24832 & ~n24833;
  assign n24835 = ~n24408 & n24411;
  assign n24836 = n24408 & ~n24411;
  assign n24837 = ~n24835 & ~n24836;
  assign n24838 = ~n24462 & n24837;
  assign n24839 = ~n24402 & ~n24637;
  assign n24840 = n24838 & ~n24839;
  assign n24841 = ~n24834 & ~n24840;
  assign n24842 = n24307 & n24841;
  assign n24843 = ~n24823 & ~n24824;
  assign n24844 = ~n24825 & n24843;
  assign n24845 = ~n24831 & n24844;
  assign n3181 = n24842 | ~n24845;
  assign n24847 = ~n22796 & ~n24261;
  assign n24848 = ~n24248 & ~n24847;
  assign n24849 = ~n24254 & n24257;
  assign n24850 = n24254 & ~n24257;
  assign n24851 = ~n24849 & ~n24850;
  assign n24852 = n24848 & ~n24851;
  assign n24853 = ~n24848 & n24851;
  assign n24854 = ~n24852 & ~n24853;
  assign n24855 = n24307 & ~n24854;
  assign n24856 = ~n22885 & ~n24855;
  assign n24857 = ~n19643 & ~n24084;
  assign n24858 = n24856 & ~n24857;
  assign n24859 = P4_REG3_REG_1_ & ~n24080;
  assign n24860 = ~n19659 & n24087;
  assign n24861 = ~n19599 & n24089;
  assign n24862 = P4_REG3_REG_1_ & ~n24063;
  assign n24863 = ~n24860 & ~n24861;
  assign n24864 = ~n24862 & n24863;
  assign n24865 = n24086 & ~n24864;
  assign n24866 = n24858 & ~n24859;
  assign n3186 = n24865 | ~n24866;
  assign n24868 = ~n20033 & ~n24080;
  assign n24869 = ~n20116 & ~n24084;
  assign n24870 = ~n20109 & n24087;
  assign n24871 = ~n19965 & n24089;
  assign n24872 = ~n20033 & ~n24063;
  assign n24873 = ~n24870 & ~n24871;
  assign n24874 = ~n24872 & n24873;
  assign n24875 = n24086 & ~n24874;
  assign n24876 = n24161 & ~n24167;
  assign n24877 = ~n24161 & n24167;
  assign n24878 = ~n24876 & ~n24877;
  assign n24879 = n24272 & ~n24878;
  assign n24880 = ~n24272 & n24878;
  assign n24881 = ~n24879 & ~n24880;
  assign n24882 = n24307 & ~n24881;
  assign n24883 = ~n22646 & ~n24882;
  assign n24884 = ~n24868 & ~n24869;
  assign n24885 = ~n24875 & n24884;
  assign n3191 = ~n24883 | ~n24885;
  assign n24887 = ~n21416 & n24315;
  assign n24888 = n21485 & n24319;
  assign n24889 = P4_REG3_REG_28_ & ~P4_STATE_REG;
  assign n24890 = ~n21483 & n24087;
  assign n24891 = ~n21416 & ~n24063;
  assign n24892 = ~n21353 & n24089;
  assign n24893 = ~n24890 & ~n24891;
  assign n24894 = ~n24892 & n24893;
  assign n24895 = n24086 & ~n24894;
  assign n24896 = n24337 & ~n24348;
  assign n24897 = ~n21353 & n22775;
  assign n24898 = n21422 & ~n22788;
  assign n24899 = ~n24897 & ~n24898;
  assign n24900 = ~n22793 & ~n24899;
  assign n24901 = n22793 & n24899;
  assign n24902 = ~n24900 & ~n24901;
  assign n24903 = ~n21353 & ~n22785;
  assign n24904 = n21422 & n22775;
  assign n24905 = ~n24903 & ~n24904;
  assign n24906 = n24902 & n24905;
  assign n24907 = ~n24348 & n24477;
  assign n24908 = ~n24896 & ~n24906;
  assign n24909 = ~n24347 & n24908;
  assign n24910 = ~n24907 & n24909;
  assign n24911 = ~n24902 & ~n24905;
  assign n24912 = ~n24910 & ~n24911;
  assign n24913 = ~n24337 & ~n24360;
  assign n24914 = ~n24347 & n24913;
  assign n24915 = ~n24906 & n24914;
  assign n24916 = ~n24472 & n24915;
  assign n24917 = ~n21420 & ~n22785;
  assign n24918 = n21485 & n22775;
  assign n24919 = ~n24917 & ~n24918;
  assign n24920 = ~n22793 & ~n24919;
  assign n24921 = n22793 & n24919;
  assign n24922 = ~n24920 & ~n24921;
  assign n24923 = ~n21420 & n22775;
  assign n24924 = n21485 & ~n22788;
  assign n24925 = ~n24923 & ~n24924;
  assign n24926 = ~n24922 & n24925;
  assign n24927 = n24922 & ~n24925;
  assign n24928 = ~n24926 & ~n24927;
  assign n24929 = n24912 & ~n24916;
  assign n24930 = ~n24928 & n24929;
  assign n24931 = ~n24472 & n24914;
  assign n24932 = ~n24337 & ~n24477;
  assign n24933 = ~n24347 & n24932;
  assign n24934 = ~n24911 & ~n24933;
  assign n24935 = ~n24348 & ~n24931;
  assign n24936 = n24934 & n24935;
  assign n24937 = ~n24906 & ~n24936;
  assign n24938 = n24928 & n24937;
  assign n24939 = ~n24930 & ~n24938;
  assign n24940 = n24307 & ~n24939;
  assign n24941 = ~n24887 & ~n24888;
  assign n24942 = ~n24889 & n24941;
  assign n24943 = ~n24895 & n24942;
  assign n3196 = n24940 | ~n24943;
  assign n24945 = ~n20814 & ~n24080;
  assign n24946 = ~n20895 & ~n24084;
  assign n24947 = ~n20889 & n24087;
  assign n24948 = ~n20742 & n24089;
  assign n24949 = ~n20814 & ~n24063;
  assign n24950 = ~n24947 & ~n24948;
  assign n24951 = ~n24949 & n24950;
  assign n24952 = n24086 & ~n24951;
  assign n24953 = ~n24388 & n24391;
  assign n24954 = n24388 & ~n24391;
  assign n24955 = ~n24953 & ~n24954;
  assign n24956 = n24459 & ~n24955;
  assign n24957 = ~n24392 & ~n24464;
  assign n24958 = ~n24459 & ~n24957;
  assign n24959 = ~n24956 & ~n24958;
  assign n24960 = n24307 & ~n24959;
  assign n24961 = ~n24945 & ~n24946;
  assign n24962 = ~n22266 & n24961;
  assign n24963 = ~n24952 & n24962;
  assign n3201 = n24960 | ~n24963;
  assign n24965 = ~n24222 & ~n24241;
  assign n24966 = n24247 & ~n24965;
  assign n24967 = ~n24233 & n24265;
  assign n24968 = n24966 & ~n24967;
  assign n24969 = n24222 & ~n24241;
  assign n24970 = ~n24222 & n24241;
  assign n24971 = ~n24969 & ~n24970;
  assign n24972 = ~n24233 & n24971;
  assign n24973 = ~n24245 & ~n24265;
  assign n24974 = n24972 & ~n24973;
  assign n24975 = ~n24968 & ~n24974;
  assign n24976 = n24307 & n24975;
  assign n24977 = ~n22825 & ~n24976;
  assign n24978 = ~n19770 & ~n24084;
  assign n24979 = n24977 & ~n24978;
  assign n24980 = ~P4_REG3_REG_3_ & ~n24080;
  assign n24981 = ~n19763 & n24087;
  assign n24982 = ~n19659 & n24089;
  assign n24983 = ~P4_REG3_REG_3_ & ~n24063;
  assign n24984 = ~n24981 & ~n24982;
  assign n24985 = ~n24983 & n24984;
  assign n24986 = n24086 & ~n24985;
  assign n24987 = n24979 & ~n24980;
  assign n3206 = n24986 | ~n24987;
  assign n24989 = ~n20171 & ~n24080;
  assign n24990 = ~n20254 & ~n24084;
  assign n24991 = ~n20247 & n24087;
  assign n24992 = ~n20109 & n24089;
  assign n24993 = ~n20171 & ~n24063;
  assign n24994 = ~n24991 & ~n24992;
  assign n24995 = ~n24993 & n24994;
  assign n24996 = n24086 & ~n24995;
  assign n24997 = n24140 & ~n24146;
  assign n24998 = ~n24140 & n24146;
  assign n24999 = ~n24997 & ~n24998;
  assign n25000 = n24277 & ~n24999;
  assign n25001 = ~n24277 & n24999;
  assign n25002 = ~n25000 & ~n25001;
  assign n25003 = n24307 & ~n25002;
  assign n25004 = ~n24989 & ~n24990;
  assign n25005 = ~n22592 & n25004;
  assign n25006 = ~n24996 & n25005;
  assign n3211 = n25003 | ~n25006;
  assign n25008 = ~n21083 & n24315;
  assign n25009 = n21158 & n24319;
  assign n25010 = P4_REG3_REG_23_ & ~P4_STATE_REG;
  assign n25011 = ~n21154 & n24087;
  assign n25012 = ~n21021 & n24089;
  assign n25013 = ~n21083 & ~n24063;
  assign n25014 = ~n25011 & ~n25012;
  assign n25015 = ~n25013 & n25014;
  assign n25016 = n24086 & ~n25015;
  assign n25017 = n24363 & ~n24369;
  assign n25018 = ~n24363 & n24369;
  assign n25019 = ~n25017 & ~n25018;
  assign n25020 = n24470 & ~n25019;
  assign n25021 = ~n24470 & n25019;
  assign n25022 = ~n25020 & ~n25021;
  assign n25023 = n24307 & ~n25022;
  assign n25024 = ~n25008 & ~n25009;
  assign n25025 = ~n25010 & n25024;
  assign n25026 = ~n25016 & n25025;
  assign n3216 = n25023 | ~n25026;
  assign n25028 = ~n20458 & ~n24080;
  assign n25029 = ~n20540 & ~n24084;
  assign n25030 = ~n20533 & n24087;
  assign n25031 = ~n20390 & n24089;
  assign n25032 = ~n20458 & ~n24063;
  assign n25033 = ~n25030 & ~n25031;
  assign n25034 = ~n25032 & n25033;
  assign n25035 = n24086 & ~n25034;
  assign n25036 = n24097 & ~n24103;
  assign n25037 = ~n24097 & n24103;
  assign n25038 = ~n25036 & ~n25037;
  assign n25039 = n24288 & ~n25038;
  assign n25040 = ~n24288 & n25038;
  assign n25041 = ~n25039 & ~n25040;
  assign n25042 = n24307 & ~n25041;
  assign n25043 = ~n25028 & ~n25029;
  assign n25044 = ~n22484 & n25043;
  assign n25045 = ~n25035 & n25044;
  assign n3221 = n25042 | ~n25045;
  assign n25047 = ~n21349 & n24315;
  assign n25048 = n21422 & n24319;
  assign n25049 = P4_REG3_REG_27_ & ~P4_STATE_REG;
  assign n25050 = ~n21349 & ~n24063;
  assign n25051 = ~n21289 & n24089;
  assign n25052 = ~n21420 & n24087;
  assign n25053 = ~n25050 & ~n25051;
  assign n25054 = ~n25052 & n25053;
  assign n25055 = n24086 & ~n25054;
  assign n25056 = ~n24347 & ~n24907;
  assign n25057 = ~n24896 & n25056;
  assign n25058 = ~n24931 & ~n25057;
  assign n25059 = ~n24902 & n24905;
  assign n25060 = n24902 & ~n24905;
  assign n25061 = ~n25059 & ~n25060;
  assign n25062 = n25058 & ~n25061;
  assign n25063 = ~n25058 & n25061;
  assign n25064 = ~n25062 & ~n25063;
  assign n25065 = n24307 & ~n25064;
  assign n25066 = ~n25047 & ~n25048;
  assign n25067 = ~n25049 & n25066;
  assign n25068 = ~n25055 & n25067;
  assign n3226 = n25065 | ~n25068;
  assign n25070 = ~n19958 & ~n24080;
  assign n25071 = ~n20047 & ~n24084;
  assign n25072 = ~n20040 & n24087;
  assign n25073 = ~n19901 & n24089;
  assign n25074 = ~n19958 & ~n24063;
  assign n25075 = ~n25072 & ~n25073;
  assign n25076 = ~n25074 & n25075;
  assign n25077 = n24086 & ~n25076;
  assign n25078 = ~n24195 & ~n24198;
  assign n25079 = n24200 & ~n25078;
  assign n25080 = ~n24202 & n24504;
  assign n25081 = n25079 & ~n25080;
  assign n25082 = ~n24195 & n24198;
  assign n25083 = n24195 & ~n24198;
  assign n25084 = ~n25082 & ~n25083;
  assign n25085 = ~n24202 & n25084;
  assign n25086 = ~n24189 & ~n24504;
  assign n25087 = n25085 & ~n25086;
  assign n25088 = ~n25081 & ~n25087;
  assign n25089 = n24307 & n25088;
  assign n25090 = ~n22669 & ~n25089;
  assign n25091 = ~n25070 & ~n25071;
  assign n25092 = ~n25077 & n25091;
  assign n3231 = ~n25090 | ~n25092;
  assign n25094 = P1_P3_STATE_REG_1_ & ~P1_P3_STATE_REG_0_;
  assign n25095 = P1_P3_BYTEENABLE_REG_3_ & n25094;
  assign n25096 = P1_P3_BE_N_REG_3_ & ~n25094;
  assign n3251 = n25095 | n25096;
  assign n25098 = P1_P3_BYTEENABLE_REG_2_ & n25094;
  assign n25099 = P1_P3_BE_N_REG_2_ & ~n25094;
  assign n3256 = n25098 | n25099;
  assign n25101 = P1_P3_BYTEENABLE_REG_1_ & n25094;
  assign n25102 = P1_P3_BE_N_REG_1_ & ~n25094;
  assign n3261 = n25101 | n25102;
  assign n25104 = P1_P3_BYTEENABLE_REG_0_ & n25094;
  assign n25105 = P1_P3_BE_N_REG_0_ & ~n25094;
  assign n3266 = n25104 | n25105;
  assign n25107 = P1_P3_STATE_REG_2_ & n25094;
  assign n25108 = P1_P3_REIP_REG_30_ & n25107;
  assign n25109 = ~P1_P3_STATE_REG_2_ & n25094;
  assign n25110 = P1_P3_REIP_REG_31_ & n25109;
  assign n25111 = P1_P3_ADDRESS_REG_29_ & ~n25094;
  assign n25112 = ~n25108 & ~n25110;
  assign n3271 = n25111 | ~n25112;
  assign n25114 = P1_P3_REIP_REG_29_ & n25107;
  assign n25115 = P1_P3_REIP_REG_30_ & n25109;
  assign n25116 = P1_P3_ADDRESS_REG_28_ & ~n25094;
  assign n25117 = ~n25114 & ~n25115;
  assign n3276 = n25116 | ~n25117;
  assign n25119 = P1_P3_REIP_REG_28_ & n25107;
  assign n25120 = P1_P3_REIP_REG_29_ & n25109;
  assign n25121 = P1_P3_ADDRESS_REG_27_ & ~n25094;
  assign n25122 = ~n25119 & ~n25120;
  assign n3281 = n25121 | ~n25122;
  assign n25124 = P1_P3_REIP_REG_27_ & n25107;
  assign n25125 = P1_P3_REIP_REG_28_ & n25109;
  assign n25126 = P1_P3_ADDRESS_REG_26_ & ~n25094;
  assign n25127 = ~n25124 & ~n25125;
  assign n3286 = n25126 | ~n25127;
  assign n25129 = P1_P3_REIP_REG_26_ & n25107;
  assign n25130 = P1_P3_REIP_REG_27_ & n25109;
  assign n25131 = P1_P3_ADDRESS_REG_25_ & ~n25094;
  assign n25132 = ~n25129 & ~n25130;
  assign n3291 = n25131 | ~n25132;
  assign n25134 = P1_P3_REIP_REG_25_ & n25107;
  assign n25135 = P1_P3_REIP_REG_26_ & n25109;
  assign n25136 = P1_P3_ADDRESS_REG_24_ & ~n25094;
  assign n25137 = ~n25134 & ~n25135;
  assign n3296 = n25136 | ~n25137;
  assign n25139 = P1_P3_REIP_REG_24_ & n25107;
  assign n25140 = P1_P3_REIP_REG_25_ & n25109;
  assign n25141 = P1_P3_ADDRESS_REG_23_ & ~n25094;
  assign n25142 = ~n25139 & ~n25140;
  assign n3301 = n25141 | ~n25142;
  assign n25144 = P1_P3_REIP_REG_23_ & n25107;
  assign n25145 = P1_P3_REIP_REG_24_ & n25109;
  assign n25146 = P1_P3_ADDRESS_REG_22_ & ~n25094;
  assign n25147 = ~n25144 & ~n25145;
  assign n3306 = n25146 | ~n25147;
  assign n25149 = P1_P3_REIP_REG_22_ & n25107;
  assign n25150 = P1_P3_REIP_REG_23_ & n25109;
  assign n25151 = P1_P3_ADDRESS_REG_21_ & ~n25094;
  assign n25152 = ~n25149 & ~n25150;
  assign n3311 = n25151 | ~n25152;
  assign n25154 = P1_P3_REIP_REG_21_ & n25107;
  assign n25155 = P1_P3_REIP_REG_22_ & n25109;
  assign n25156 = P1_P3_ADDRESS_REG_20_ & ~n25094;
  assign n25157 = ~n25154 & ~n25155;
  assign n3316 = n25156 | ~n25157;
  assign n25159 = P1_P3_REIP_REG_20_ & n25107;
  assign n25160 = P1_P3_REIP_REG_21_ & n25109;
  assign n25161 = P1_P3_ADDRESS_REG_19_ & ~n25094;
  assign n25162 = ~n25159 & ~n25160;
  assign n3321 = n25161 | ~n25162;
  assign n25164 = P1_P3_REIP_REG_19_ & n25107;
  assign n25165 = P1_P3_REIP_REG_20_ & n25109;
  assign n25166 = P1_P3_ADDRESS_REG_18_ & ~n25094;
  assign n25167 = ~n25164 & ~n25165;
  assign n3326 = n25166 | ~n25167;
  assign n25169 = P1_P3_REIP_REG_18_ & n25107;
  assign n25170 = P1_P3_REIP_REG_19_ & n25109;
  assign n25171 = P1_P3_ADDRESS_REG_17_ & ~n25094;
  assign n25172 = ~n25169 & ~n25170;
  assign n3331 = n25171 | ~n25172;
  assign n25174 = P1_P3_REIP_REG_17_ & n25107;
  assign n25175 = P1_P3_REIP_REG_18_ & n25109;
  assign n25176 = P1_P3_ADDRESS_REG_16_ & ~n25094;
  assign n25177 = ~n25174 & ~n25175;
  assign n3336 = n25176 | ~n25177;
  assign n25179 = P1_P3_REIP_REG_16_ & n25107;
  assign n25180 = P1_P3_REIP_REG_17_ & n25109;
  assign n25181 = P1_P3_ADDRESS_REG_15_ & ~n25094;
  assign n25182 = ~n25179 & ~n25180;
  assign n3341 = n25181 | ~n25182;
  assign n25184 = P1_P3_REIP_REG_15_ & n25107;
  assign n25185 = P1_P3_REIP_REG_16_ & n25109;
  assign n25186 = P1_P3_ADDRESS_REG_14_ & ~n25094;
  assign n25187 = ~n25184 & ~n25185;
  assign n3346 = n25186 | ~n25187;
  assign n25189 = P1_P3_REIP_REG_14_ & n25107;
  assign n25190 = P1_P3_REIP_REG_15_ & n25109;
  assign n25191 = P1_P3_ADDRESS_REG_13_ & ~n25094;
  assign n25192 = ~n25189 & ~n25190;
  assign n3351 = n25191 | ~n25192;
  assign n25194 = P1_P3_REIP_REG_13_ & n25107;
  assign n25195 = P1_P3_REIP_REG_14_ & n25109;
  assign n25196 = P1_P3_ADDRESS_REG_12_ & ~n25094;
  assign n25197 = ~n25194 & ~n25195;
  assign n3356 = n25196 | ~n25197;
  assign n25199 = P1_P3_REIP_REG_12_ & n25107;
  assign n25200 = P1_P3_REIP_REG_13_ & n25109;
  assign n25201 = P1_P3_ADDRESS_REG_11_ & ~n25094;
  assign n25202 = ~n25199 & ~n25200;
  assign n3361 = n25201 | ~n25202;
  assign n25204 = P1_P3_REIP_REG_11_ & n25107;
  assign n25205 = P1_P3_REIP_REG_12_ & n25109;
  assign n25206 = P1_P3_ADDRESS_REG_10_ & ~n25094;
  assign n25207 = ~n25204 & ~n25205;
  assign n3366 = n25206 | ~n25207;
  assign n25209 = P1_P3_REIP_REG_10_ & n25107;
  assign n25210 = P1_P3_REIP_REG_11_ & n25109;
  assign n25211 = P1_P3_ADDRESS_REG_9_ & ~n25094;
  assign n25212 = ~n25209 & ~n25210;
  assign n3371 = n25211 | ~n25212;
  assign n25214 = P1_P3_REIP_REG_9_ & n25107;
  assign n25215 = P1_P3_REIP_REG_10_ & n25109;
  assign n25216 = P1_P3_ADDRESS_REG_8_ & ~n25094;
  assign n25217 = ~n25214 & ~n25215;
  assign n3376 = n25216 | ~n25217;
  assign n25219 = P1_P3_REIP_REG_8_ & n25107;
  assign n25220 = P1_P3_REIP_REG_9_ & n25109;
  assign n25221 = P1_P3_ADDRESS_REG_7_ & ~n25094;
  assign n25222 = ~n25219 & ~n25220;
  assign n3381 = n25221 | ~n25222;
  assign n25224 = P1_P3_REIP_REG_7_ & n25107;
  assign n25225 = P1_P3_REIP_REG_8_ & n25109;
  assign n25226 = P1_P3_ADDRESS_REG_6_ & ~n25094;
  assign n25227 = ~n25224 & ~n25225;
  assign n3386 = n25226 | ~n25227;
  assign n25229 = P1_P3_REIP_REG_6_ & n25107;
  assign n25230 = P1_P3_REIP_REG_7_ & n25109;
  assign n25231 = P1_P3_ADDRESS_REG_5_ & ~n25094;
  assign n25232 = ~n25229 & ~n25230;
  assign n3391 = n25231 | ~n25232;
  assign n25234 = P1_P3_REIP_REG_5_ & n25107;
  assign n25235 = P1_P3_REIP_REG_6_ & n25109;
  assign n25236 = P1_P3_ADDRESS_REG_4_ & ~n25094;
  assign n25237 = ~n25234 & ~n25235;
  assign n3396 = n25236 | ~n25237;
  assign n25239 = P1_P3_REIP_REG_4_ & n25107;
  assign n25240 = P1_P3_REIP_REG_5_ & n25109;
  assign n25241 = P1_P3_ADDRESS_REG_3_ & ~n25094;
  assign n25242 = ~n25239 & ~n25240;
  assign n3401 = n25241 | ~n25242;
  assign n25244 = P1_P3_REIP_REG_3_ & n25107;
  assign n25245 = P1_P3_REIP_REG_4_ & n25109;
  assign n25246 = P1_P3_ADDRESS_REG_2_ & ~n25094;
  assign n25247 = ~n25244 & ~n25245;
  assign n3406 = n25246 | ~n25247;
  assign n25249 = P1_P3_REIP_REG_2_ & n25107;
  assign n25250 = P1_P3_REIP_REG_3_ & n25109;
  assign n25251 = P1_P3_ADDRESS_REG_1_ & ~n25094;
  assign n25252 = ~n25249 & ~n25250;
  assign n3411 = n25251 | ~n25252;
  assign n25254 = P1_P3_REIP_REG_1_ & n25107;
  assign n25255 = P1_P3_REIP_REG_2_ & n25109;
  assign n25256 = P1_P3_ADDRESS_REG_0_ & ~n25094;
  assign n25257 = ~n25254 & ~n25255;
  assign n3416 = n25256 | ~n25257;
  assign n25259 = ~P1_P3_STATE_REG_2_ & P1_P3_STATE_REG_1_;
  assign n25260 = NA & n25259;
  assign n25261 = P1_P3_STATE_REG_0_ & ~n25260;
  assign n25262 = ~HOLD & ~P1_P3_REQUESTPENDING_REG;
  assign n25263 = P1_P3_W_R_N_REG & ~P1_P3_ADS_N_REG;
  assign n25264 = P3_RD_REG & n25263;
  assign n25265 = P1_P3_D_C_N_REG & n25264;
  assign n25266 = P1_P3_M_IO_N_REG & n25265;
  assign n25267 = P1_READY22_REG & ~n25266;
  assign n25268 = n25259 & ~n25262;
  assign n25269 = n25267 & n25268;
  assign n25270 = ~P1_P3_STATE_REG_2_ & ~P1_P3_STATE_REG_1_;
  assign n25271 = HOLD & ~P1_P3_REQUESTPENDING_REG;
  assign n25272 = n25270 & n25271;
  assign n25273 = ~n25269 & ~n25272;
  assign n25274 = n25261 & ~n25273;
  assign n25275 = ~n25107 & ~n25274;
  assign n25276 = ~HOLD & P1_P3_REQUESTPENDING_REG;
  assign n25277 = P1_P3_STATE_REG_0_ & ~n25276;
  assign n25278 = ~n25262 & n25277;
  assign n25279 = ~NA & ~P1_P3_STATE_REG_0_;
  assign n25280 = n25262 & ~n25267;
  assign n25281 = ~n25267 & n25276;
  assign n25282 = ~n25280 & ~n25281;
  assign n25283 = P1_P3_STATE_REG_1_ & n25282;
  assign n25284 = ~n25278 & ~n25279;
  assign n25285 = ~n25283 & n25284;
  assign n25286 = P1_P3_STATE_REG_2_ & ~n25285;
  assign n3421 = ~n25275 | n25286;
  assign n25288 = P1_P3_STATE_REG_2_ & ~n25277;
  assign n25289 = P1_P3_STATE_REG_0_ & P1_P3_REQUESTPENDING_REG;
  assign n25290 = ~P1_P3_STATE_REG_2_ & n25289;
  assign n25291 = ~n25288 & ~n25290;
  assign n25292 = ~P1_P3_STATE_REG_1_ & ~n25291;
  assign n25293 = HOLD & ~n25267;
  assign n25294 = P1_P3_STATE_REG_0_ & ~n25293;
  assign n25295 = P1_P3_STATE_REG_2_ & ~n25294;
  assign n25296 = ~n25280 & ~n25295;
  assign n25297 = P1_P3_STATE_REG_1_ & n25296;
  assign n25298 = n25094 & n25267;
  assign n25299 = ~n25109 & ~n25298;
  assign n25300 = ~n25292 & ~n25297;
  assign n3426 = ~n25299 | ~n25300;
  assign n25302 = P1_P3_STATE_REG_1_ & ~n25281;
  assign n25303 = n25289 & ~n25302;
  assign n25304 = ~P1_P3_STATE_REG_2_ & ~n25303;
  assign n25305 = P1_P3_STATE_REG_2_ & n25277;
  assign n25306 = NA & ~P1_P3_STATE_REG_0_;
  assign n25307 = P1_P3_STATE_REG_2_ & ~n25276;
  assign n25308 = ~n25306 & ~n25307;
  assign n25309 = ~P1_P3_STATE_REG_1_ & ~n25308;
  assign n25310 = ~n25304 & ~n25305;
  assign n3431 = n25309 | ~n25310;
  assign n25312 = ~BS & ~n25270;
  assign n25313 = P1_P3_STATE_REG_0_ & n25259;
  assign n25314 = ~P1_P3_STATE_REG_1_ & ~P1_P3_STATE_REG_0_;
  assign n25315 = ~n25313 & ~n25314;
  assign n25316 = n25312 & ~n25315;
  assign n25317 = P1_P3_DATAWIDTH_REG_0_ & n25315;
  assign n3436 = n25316 | n25317;
  assign n25319 = P1_P3_DATAWIDTH_REG_1_ & n25315;
  assign n25320 = ~n25312 & ~n25315;
  assign n3441 = n25319 | n25320;
  assign n3446 = P1_P3_DATAWIDTH_REG_2_ & n25315;
  assign n3451 = P1_P3_DATAWIDTH_REG_3_ & n25315;
  assign n3456 = P1_P3_DATAWIDTH_REG_4_ & n25315;
  assign n3461 = P1_P3_DATAWIDTH_REG_5_ & n25315;
  assign n3466 = P1_P3_DATAWIDTH_REG_6_ & n25315;
  assign n3471 = P1_P3_DATAWIDTH_REG_7_ & n25315;
  assign n3476 = P1_P3_DATAWIDTH_REG_8_ & n25315;
  assign n3481 = P1_P3_DATAWIDTH_REG_9_ & n25315;
  assign n3486 = P1_P3_DATAWIDTH_REG_10_ & n25315;
  assign n3491 = P1_P3_DATAWIDTH_REG_11_ & n25315;
  assign n3496 = P1_P3_DATAWIDTH_REG_12_ & n25315;
  assign n3501 = P1_P3_DATAWIDTH_REG_13_ & n25315;
  assign n3506 = P1_P3_DATAWIDTH_REG_14_ & n25315;
  assign n3511 = P1_P3_DATAWIDTH_REG_15_ & n25315;
  assign n3516 = P1_P3_DATAWIDTH_REG_16_ & n25315;
  assign n3521 = P1_P3_DATAWIDTH_REG_17_ & n25315;
  assign n3526 = P1_P3_DATAWIDTH_REG_18_ & n25315;
  assign n3531 = P1_P3_DATAWIDTH_REG_19_ & n25315;
  assign n3536 = P1_P3_DATAWIDTH_REG_20_ & n25315;
  assign n3541 = P1_P3_DATAWIDTH_REG_21_ & n25315;
  assign n3546 = P1_P3_DATAWIDTH_REG_22_ & n25315;
  assign n3551 = P1_P3_DATAWIDTH_REG_23_ & n25315;
  assign n3556 = P1_P3_DATAWIDTH_REG_24_ & n25315;
  assign n3561 = P1_P3_DATAWIDTH_REG_25_ & n25315;
  assign n3566 = P1_P3_DATAWIDTH_REG_26_ & n25315;
  assign n3571 = P1_P3_DATAWIDTH_REG_27_ & n25315;
  assign n3576 = P1_P3_DATAWIDTH_REG_28_ & n25315;
  assign n3581 = P1_P3_DATAWIDTH_REG_29_ & n25315;
  assign n3586 = P1_P3_DATAWIDTH_REG_30_ & n25315;
  assign n3591 = P1_P3_DATAWIDTH_REG_31_ & n25315;
  assign n25352 = P1_P3_STATE2_REG_2_ & P1_P3_STATE2_REG_1_;
  assign n25353 = P1_P3_STATE2_REG_1_ & n25267;
  assign n25354 = ~P1_P3_STATE2_REG_0_ & ~n25353;
  assign n25355 = ~P1_P3_STATEBS16_REG & ~n25267;
  assign n25356 = P1_P3_STATE_REG_2_ & ~P1_P3_STATE_REG_1_;
  assign n25357 = ~n25259 & ~n25356;
  assign n25358 = ~P1_P3_STATE_REG_0_ & ~n25357;
  assign n25359 = n25355 & n25358;
  assign n25360 = P1_P3_INSTQUEUERD_ADDR_REG_1_ & P1_P3_INSTQUEUERD_ADDR_REG_0_;
  assign n25361 = ~P1_P3_INSTQUEUERD_ADDR_REG_2_ & n25360;
  assign n25362 = P1_P3_INSTQUEUERD_ADDR_REG_3_ & n25361;
  assign n25363 = P1_P3_INSTQUEUE_REG_11__5_ & n25362;
  assign n25364 = P1_P3_INSTQUEUERD_ADDR_REG_1_ & ~P1_P3_INSTQUEUERD_ADDR_REG_0_;
  assign n25365 = ~P1_P3_INSTQUEUERD_ADDR_REG_2_ & n25364;
  assign n25366 = P1_P3_INSTQUEUERD_ADDR_REG_3_ & n25365;
  assign n25367 = P1_P3_INSTQUEUE_REG_10__5_ & n25366;
  assign n25368 = ~n25363 & ~n25367;
  assign n25369 = ~P1_P3_INSTQUEUERD_ADDR_REG_1_ & P1_P3_INSTQUEUERD_ADDR_REG_0_;
  assign n25370 = ~P1_P3_INSTQUEUERD_ADDR_REG_2_ & n25369;
  assign n25371 = P1_P3_INSTQUEUERD_ADDR_REG_3_ & n25370;
  assign n25372 = P1_P3_INSTQUEUE_REG_9__5_ & n25371;
  assign n25373 = ~P1_P3_INSTQUEUERD_ADDR_REG_1_ & ~P1_P3_INSTQUEUERD_ADDR_REG_0_;
  assign n25374 = ~P1_P3_INSTQUEUERD_ADDR_REG_2_ & n25373;
  assign n25375 = P1_P3_INSTQUEUERD_ADDR_REG_3_ & n25374;
  assign n25376 = P1_P3_INSTQUEUE_REG_8__5_ & n25375;
  assign n25377 = ~n25372 & ~n25376;
  assign n25378 = P1_P3_INSTQUEUERD_ADDR_REG_3_ & P1_P3_INSTQUEUERD_ADDR_REG_2_;
  assign n25379 = n25360 & n25378;
  assign n25380 = P1_P3_INSTQUEUE_REG_15__5_ & n25379;
  assign n25381 = n25364 & n25378;
  assign n25382 = P1_P3_INSTQUEUE_REG_14__5_ & n25381;
  assign n25383 = n25369 & n25378;
  assign n25384 = P1_P3_INSTQUEUE_REG_13__5_ & n25383;
  assign n25385 = n25373 & n25378;
  assign n25386 = P1_P3_INSTQUEUE_REG_12__5_ & n25385;
  assign n25387 = ~n25380 & ~n25382;
  assign n25388 = ~n25384 & n25387;
  assign n25389 = ~n25386 & n25388;
  assign n25390 = ~P1_P3_INSTQUEUERD_ADDR_REG_3_ & P1_P3_INSTQUEUERD_ADDR_REG_2_;
  assign n25391 = n25360 & n25390;
  assign n25392 = P1_P3_INSTQUEUE_REG_7__5_ & n25391;
  assign n25393 = n25364 & n25390;
  assign n25394 = P1_P3_INSTQUEUE_REG_6__5_ & n25393;
  assign n25395 = n25369 & n25390;
  assign n25396 = P1_P3_INSTQUEUE_REG_5__5_ & n25395;
  assign n25397 = n25373 & n25390;
  assign n25398 = P1_P3_INSTQUEUE_REG_4__5_ & n25397;
  assign n25399 = ~n25392 & ~n25394;
  assign n25400 = ~n25396 & n25399;
  assign n25401 = ~n25398 & n25400;
  assign n25402 = ~P1_P3_INSTQUEUERD_ADDR_REG_3_ & n25361;
  assign n25403 = P1_P3_INSTQUEUE_REG_3__5_ & n25402;
  assign n25404 = ~P1_P3_INSTQUEUERD_ADDR_REG_3_ & ~P1_P3_INSTQUEUERD_ADDR_REG_2_;
  assign n25405 = n25364 & n25404;
  assign n25406 = P1_P3_INSTQUEUE_REG_2__5_ & n25405;
  assign n25407 = n25369 & n25404;
  assign n25408 = P1_P3_INSTQUEUE_REG_1__5_ & n25407;
  assign n25409 = ~P1_P3_INSTQUEUERD_ADDR_REG_3_ & n25374;
  assign n25410 = P1_P3_INSTQUEUE_REG_0__5_ & n25409;
  assign n25411 = ~n25403 & ~n25406;
  assign n25412 = ~n25408 & n25411;
  assign n25413 = ~n25410 & n25412;
  assign n25414 = n25368 & n25377;
  assign n25415 = n25389 & n25414;
  assign n25416 = n25401 & n25415;
  assign n25417 = n25413 & n25416;
  assign n25418 = P1_P3_INSTQUEUE_REG_11__6_ & n25362;
  assign n25419 = P1_P3_INSTQUEUE_REG_10__6_ & n25366;
  assign n25420 = ~n25418 & ~n25419;
  assign n25421 = P1_P3_INSTQUEUE_REG_9__6_ & n25371;
  assign n25422 = P1_P3_INSTQUEUE_REG_8__6_ & n25375;
  assign n25423 = ~n25421 & ~n25422;
  assign n25424 = P1_P3_INSTQUEUE_REG_15__6_ & n25379;
  assign n25425 = P1_P3_INSTQUEUE_REG_14__6_ & n25381;
  assign n25426 = P1_P3_INSTQUEUE_REG_13__6_ & n25383;
  assign n25427 = P1_P3_INSTQUEUE_REG_12__6_ & n25385;
  assign n25428 = ~n25424 & ~n25425;
  assign n25429 = ~n25426 & n25428;
  assign n25430 = ~n25427 & n25429;
  assign n25431 = P1_P3_INSTQUEUE_REG_7__6_ & n25391;
  assign n25432 = P1_P3_INSTQUEUE_REG_6__6_ & n25393;
  assign n25433 = P1_P3_INSTQUEUE_REG_5__6_ & n25395;
  assign n25434 = P1_P3_INSTQUEUE_REG_4__6_ & n25397;
  assign n25435 = ~n25431 & ~n25432;
  assign n25436 = ~n25433 & n25435;
  assign n25437 = ~n25434 & n25436;
  assign n25438 = P1_P3_INSTQUEUE_REG_3__6_ & n25402;
  assign n25439 = P1_P3_INSTQUEUE_REG_2__6_ & n25405;
  assign n25440 = P1_P3_INSTQUEUE_REG_1__6_ & n25407;
  assign n25441 = P1_P3_INSTQUEUE_REG_0__6_ & n25409;
  assign n25442 = ~n25438 & ~n25439;
  assign n25443 = ~n25440 & n25442;
  assign n25444 = ~n25441 & n25443;
  assign n25445 = n25420 & n25423;
  assign n25446 = n25430 & n25445;
  assign n25447 = n25437 & n25446;
  assign n25448 = n25444 & n25447;
  assign n25449 = n25417 & n25448;
  assign n25450 = P1_P3_INSTQUEUE_REG_11__4_ & n25362;
  assign n25451 = P1_P3_INSTQUEUE_REG_10__4_ & n25366;
  assign n25452 = ~n25450 & ~n25451;
  assign n25453 = P1_P3_INSTQUEUE_REG_9__4_ & n25371;
  assign n25454 = P1_P3_INSTQUEUE_REG_8__4_ & n25375;
  assign n25455 = ~n25453 & ~n25454;
  assign n25456 = P1_P3_INSTQUEUE_REG_15__4_ & n25379;
  assign n25457 = P1_P3_INSTQUEUE_REG_14__4_ & n25381;
  assign n25458 = P1_P3_INSTQUEUE_REG_13__4_ & n25383;
  assign n25459 = P1_P3_INSTQUEUE_REG_12__4_ & n25385;
  assign n25460 = ~n25456 & ~n25457;
  assign n25461 = ~n25458 & n25460;
  assign n25462 = ~n25459 & n25461;
  assign n25463 = P1_P3_INSTQUEUE_REG_7__4_ & n25391;
  assign n25464 = P1_P3_INSTQUEUE_REG_6__4_ & n25393;
  assign n25465 = P1_P3_INSTQUEUE_REG_5__4_ & n25395;
  assign n25466 = P1_P3_INSTQUEUE_REG_4__4_ & n25397;
  assign n25467 = ~n25463 & ~n25464;
  assign n25468 = ~n25465 & n25467;
  assign n25469 = ~n25466 & n25468;
  assign n25470 = P1_P3_INSTQUEUE_REG_3__4_ & n25402;
  assign n25471 = P1_P3_INSTQUEUE_REG_2__4_ & n25405;
  assign n25472 = P1_P3_INSTQUEUE_REG_1__4_ & n25407;
  assign n25473 = P1_P3_INSTQUEUE_REG_0__4_ & n25409;
  assign n25474 = ~n25470 & ~n25471;
  assign n25475 = ~n25472 & n25474;
  assign n25476 = ~n25473 & n25475;
  assign n25477 = n25452 & n25455;
  assign n25478 = n25462 & n25477;
  assign n25479 = n25469 & n25478;
  assign n25480 = n25476 & n25479;
  assign n25481 = P1_P3_INSTQUEUE_REG_11__7_ & n25362;
  assign n25482 = P1_P3_INSTQUEUE_REG_10__7_ & n25366;
  assign n25483 = ~n25481 & ~n25482;
  assign n25484 = P1_P3_INSTQUEUE_REG_9__7_ & n25371;
  assign n25485 = P1_P3_INSTQUEUE_REG_8__7_ & n25375;
  assign n25486 = ~n25484 & ~n25485;
  assign n25487 = P1_P3_INSTQUEUE_REG_15__7_ & n25379;
  assign n25488 = P1_P3_INSTQUEUE_REG_14__7_ & n25381;
  assign n25489 = P1_P3_INSTQUEUE_REG_13__7_ & n25383;
  assign n25490 = P1_P3_INSTQUEUE_REG_12__7_ & n25385;
  assign n25491 = ~n25487 & ~n25488;
  assign n25492 = ~n25489 & n25491;
  assign n25493 = ~n25490 & n25492;
  assign n25494 = P1_P3_INSTQUEUE_REG_7__7_ & n25391;
  assign n25495 = P1_P3_INSTQUEUE_REG_6__7_ & n25393;
  assign n25496 = P1_P3_INSTQUEUE_REG_5__7_ & n25395;
  assign n25497 = P1_P3_INSTQUEUE_REG_4__7_ & n25397;
  assign n25498 = ~n25494 & ~n25495;
  assign n25499 = ~n25496 & n25498;
  assign n25500 = ~n25497 & n25499;
  assign n25501 = P1_P3_INSTQUEUE_REG_3__7_ & n25402;
  assign n25502 = P1_P3_INSTQUEUE_REG_2__7_ & n25405;
  assign n25503 = P1_P3_INSTQUEUE_REG_1__7_ & n25407;
  assign n25504 = P1_P3_INSTQUEUE_REG_0__7_ & n25409;
  assign n25505 = ~n25501 & ~n25502;
  assign n25506 = ~n25503 & n25505;
  assign n25507 = ~n25504 & n25506;
  assign n25508 = n25483 & n25486;
  assign n25509 = n25493 & n25508;
  assign n25510 = n25500 & n25509;
  assign n25511 = n25507 & n25510;
  assign n25512 = P1_P3_INSTQUEUE_REG_11__3_ & n25362;
  assign n25513 = P1_P3_INSTQUEUE_REG_10__3_ & n25366;
  assign n25514 = ~n25512 & ~n25513;
  assign n25515 = P1_P3_INSTQUEUE_REG_9__3_ & n25371;
  assign n25516 = P1_P3_INSTQUEUE_REG_8__3_ & n25375;
  assign n25517 = ~n25515 & ~n25516;
  assign n25518 = P1_P3_INSTQUEUE_REG_15__3_ & n25379;
  assign n25519 = P1_P3_INSTQUEUE_REG_14__3_ & n25381;
  assign n25520 = P1_P3_INSTQUEUE_REG_13__3_ & n25383;
  assign n25521 = P1_P3_INSTQUEUE_REG_12__3_ & n25385;
  assign n25522 = ~n25518 & ~n25519;
  assign n25523 = ~n25520 & n25522;
  assign n25524 = ~n25521 & n25523;
  assign n25525 = P1_P3_INSTQUEUE_REG_7__3_ & n25391;
  assign n25526 = P1_P3_INSTQUEUE_REG_6__3_ & n25393;
  assign n25527 = P1_P3_INSTQUEUE_REG_5__3_ & n25395;
  assign n25528 = P1_P3_INSTQUEUE_REG_4__3_ & n25397;
  assign n25529 = ~n25525 & ~n25526;
  assign n25530 = ~n25527 & n25529;
  assign n25531 = ~n25528 & n25530;
  assign n25532 = P1_P3_INSTQUEUE_REG_3__3_ & n25402;
  assign n25533 = P1_P3_INSTQUEUE_REG_2__3_ & n25405;
  assign n25534 = P1_P3_INSTQUEUE_REG_1__3_ & n25407;
  assign n25535 = P1_P3_INSTQUEUE_REG_0__3_ & n25409;
  assign n25536 = ~n25532 & ~n25533;
  assign n25537 = ~n25534 & n25536;
  assign n25538 = ~n25535 & n25537;
  assign n25539 = n25514 & n25517;
  assign n25540 = n25524 & n25539;
  assign n25541 = n25531 & n25540;
  assign n25542 = n25538 & n25541;
  assign n25543 = P1_P3_INSTQUEUE_REG_11__2_ & n25362;
  assign n25544 = P1_P3_INSTQUEUE_REG_10__2_ & n25366;
  assign n25545 = ~n25543 & ~n25544;
  assign n25546 = P1_P3_INSTQUEUE_REG_9__2_ & n25371;
  assign n25547 = P1_P3_INSTQUEUE_REG_8__2_ & n25375;
  assign n25548 = ~n25546 & ~n25547;
  assign n25549 = P1_P3_INSTQUEUE_REG_15__2_ & n25379;
  assign n25550 = P1_P3_INSTQUEUE_REG_14__2_ & n25381;
  assign n25551 = P1_P3_INSTQUEUE_REG_13__2_ & n25383;
  assign n25552 = P1_P3_INSTQUEUE_REG_12__2_ & n25385;
  assign n25553 = ~n25549 & ~n25550;
  assign n25554 = ~n25551 & n25553;
  assign n25555 = ~n25552 & n25554;
  assign n25556 = P1_P3_INSTQUEUE_REG_7__2_ & n25391;
  assign n25557 = P1_P3_INSTQUEUE_REG_6__2_ & n25393;
  assign n25558 = P1_P3_INSTQUEUE_REG_5__2_ & n25395;
  assign n25559 = P1_P3_INSTQUEUE_REG_4__2_ & n25397;
  assign n25560 = ~n25556 & ~n25557;
  assign n25561 = ~n25558 & n25560;
  assign n25562 = ~n25559 & n25561;
  assign n25563 = P1_P3_INSTQUEUE_REG_3__2_ & n25402;
  assign n25564 = P1_P3_INSTQUEUE_REG_2__2_ & n25405;
  assign n25565 = P1_P3_INSTQUEUE_REG_1__2_ & n25407;
  assign n25566 = P1_P3_INSTQUEUE_REG_0__2_ & n25409;
  assign n25567 = ~n25563 & ~n25564;
  assign n25568 = ~n25565 & n25567;
  assign n25569 = ~n25566 & n25568;
  assign n25570 = n25545 & n25548;
  assign n25571 = n25555 & n25570;
  assign n25572 = n25562 & n25571;
  assign n25573 = n25569 & n25572;
  assign n25574 = ~n25511 & ~n25542;
  assign n25575 = n25573 & n25574;
  assign n25576 = n25449 & n25480;
  assign n25577 = n25575 & n25576;
  assign n25578 = P1_P3_INSTQUEUE_REG_11__1_ & n25362;
  assign n25579 = P1_P3_INSTQUEUE_REG_10__1_ & n25366;
  assign n25580 = ~n25578 & ~n25579;
  assign n25581 = P1_P3_INSTQUEUE_REG_9__1_ & n25371;
  assign n25582 = P1_P3_INSTQUEUE_REG_8__1_ & n25375;
  assign n25583 = ~n25581 & ~n25582;
  assign n25584 = P1_P3_INSTQUEUE_REG_15__1_ & n25379;
  assign n25585 = P1_P3_INSTQUEUE_REG_14__1_ & n25381;
  assign n25586 = P1_P3_INSTQUEUE_REG_13__1_ & n25383;
  assign n25587 = P1_P3_INSTQUEUE_REG_12__1_ & n25385;
  assign n25588 = ~n25584 & ~n25585;
  assign n25589 = ~n25586 & n25588;
  assign n25590 = ~n25587 & n25589;
  assign n25591 = P1_P3_INSTQUEUE_REG_7__1_ & n25391;
  assign n25592 = P1_P3_INSTQUEUE_REG_6__1_ & n25393;
  assign n25593 = P1_P3_INSTQUEUE_REG_5__1_ & n25395;
  assign n25594 = P1_P3_INSTQUEUE_REG_4__1_ & n25397;
  assign n25595 = ~n25591 & ~n25592;
  assign n25596 = ~n25593 & n25595;
  assign n25597 = ~n25594 & n25596;
  assign n25598 = P1_P3_INSTQUEUE_REG_3__1_ & n25402;
  assign n25599 = P1_P3_INSTQUEUE_REG_2__1_ & n25405;
  assign n25600 = P1_P3_INSTQUEUE_REG_1__1_ & n25407;
  assign n25601 = P1_P3_INSTQUEUE_REG_0__1_ & n25409;
  assign n25602 = ~n25598 & ~n25599;
  assign n25603 = ~n25600 & n25602;
  assign n25604 = ~n25601 & n25603;
  assign n25605 = n25580 & n25583;
  assign n25606 = n25590 & n25605;
  assign n25607 = n25597 & n25606;
  assign n25608 = n25604 & n25607;
  assign n25609 = P1_P3_INSTQUEUE_REG_11__0_ & n25362;
  assign n25610 = P1_P3_INSTQUEUE_REG_10__0_ & n25366;
  assign n25611 = ~n25609 & ~n25610;
  assign n25612 = P1_P3_INSTQUEUE_REG_9__0_ & n25371;
  assign n25613 = P1_P3_INSTQUEUE_REG_8__0_ & n25375;
  assign n25614 = ~n25612 & ~n25613;
  assign n25615 = P1_P3_INSTQUEUE_REG_15__0_ & n25379;
  assign n25616 = P1_P3_INSTQUEUE_REG_14__0_ & n25381;
  assign n25617 = P1_P3_INSTQUEUE_REG_13__0_ & n25383;
  assign n25618 = P1_P3_INSTQUEUE_REG_12__0_ & n25385;
  assign n25619 = ~n25615 & ~n25616;
  assign n25620 = ~n25617 & n25619;
  assign n25621 = ~n25618 & n25620;
  assign n25622 = P1_P3_INSTQUEUE_REG_7__0_ & n25391;
  assign n25623 = P1_P3_INSTQUEUE_REG_6__0_ & n25393;
  assign n25624 = P1_P3_INSTQUEUE_REG_5__0_ & n25395;
  assign n25625 = P1_P3_INSTQUEUE_REG_4__0_ & n25397;
  assign n25626 = ~n25622 & ~n25623;
  assign n25627 = ~n25624 & n25626;
  assign n25628 = ~n25625 & n25627;
  assign n25629 = P1_P3_INSTQUEUE_REG_3__0_ & n25402;
  assign n25630 = P1_P3_INSTQUEUE_REG_2__0_ & n25405;
  assign n25631 = P1_P3_INSTQUEUE_REG_1__0_ & n25407;
  assign n25632 = P1_P3_INSTQUEUE_REG_0__0_ & n25409;
  assign n25633 = ~n25629 & ~n25630;
  assign n25634 = ~n25631 & n25633;
  assign n25635 = ~n25632 & n25634;
  assign n25636 = n25611 & n25614;
  assign n25637 = n25621 & n25636;
  assign n25638 = n25628 & n25637;
  assign n25639 = n25635 & n25638;
  assign n25640 = n25608 & ~n25639;
  assign n25641 = n25577 & n25640;
  assign n25642 = n25359 & n25641;
  assign n25643 = ~P1_P3_STATE2_REG_1_ & ~n25642;
  assign n25644 = ~n25267 & n25358;
  assign n25645 = ~n25573 & ~n25608;
  assign n25646 = n25644 & n25645;
  assign n25647 = ~n25267 & ~n25573;
  assign n25648 = n25608 & n25647;
  assign n25649 = ~n25267 & n25573;
  assign n25650 = n25608 & ~n25644;
  assign n25651 = n25649 & ~n25650;
  assign n25652 = ~n25646 & ~n25648;
  assign n25653 = ~n25651 & n25652;
  assign n25654 = P1_P3_INSTQUEUERD_ADDR_REG_4_ & ~P1_P3_INSTQUEUEWR_ADDR_REG_4_;
  assign n25655 = ~P1_P3_INSTQUEUERD_ADDR_REG_3_ & P1_P3_INSTQUEUEWR_ADDR_REG_3_;
  assign n25656 = P1_P3_INSTQUEUERD_ADDR_REG_3_ & ~P1_P3_INSTQUEUEWR_ADDR_REG_3_;
  assign n25657 = ~P1_P3_INSTQUEUERD_ADDR_REG_2_ & P1_P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n25658 = P1_P3_INSTQUEUERD_ADDR_REG_2_ & ~P1_P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n25659 = P1_P3_INSTQUEUERD_ADDR_REG_0_ & ~P1_P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n25660 = P1_P3_INSTQUEUEWR_ADDR_REG_1_ & ~n25659;
  assign n25661 = ~P1_P3_INSTQUEUEWR_ADDR_REG_1_ & n25659;
  assign n25662 = ~P1_P3_INSTQUEUERD_ADDR_REG_1_ & ~n25661;
  assign n25663 = ~n25660 & ~n25662;
  assign n25664 = ~n25658 & ~n25663;
  assign n25665 = ~n25657 & ~n25664;
  assign n25666 = ~n25656 & ~n25665;
  assign n25667 = ~n25655 & ~n25666;
  assign n25668 = ~P1_P3_INSTQUEUERD_ADDR_REG_4_ & P1_P3_INSTQUEUEWR_ADDR_REG_4_;
  assign n25669 = n25667 & ~n25668;
  assign n25670 = ~n25654 & ~n25669;
  assign n25671 = ~n25654 & ~n25668;
  assign n25672 = ~n25667 & ~n25671;
  assign n25673 = n25667 & n25671;
  assign n25674 = ~n25672 & ~n25673;
  assign n25675 = ~n25655 & ~n25656;
  assign n25676 = ~n25665 & ~n25675;
  assign n25677 = n25665 & n25675;
  assign n25678 = ~n25676 & ~n25677;
  assign n25679 = ~P1_P3_INSTQUEUERD_ADDR_REG_1_ & P1_P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n25680 = P1_P3_INSTQUEUERD_ADDR_REG_1_ & ~P1_P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n25681 = ~n25679 & ~n25680;
  assign n25682 = ~n25659 & ~n25681;
  assign n25683 = n25659 & n25681;
  assign n25684 = ~n25682 & ~n25683;
  assign n25685 = ~n25657 & ~n25658;
  assign n25686 = ~n25663 & ~n25685;
  assign n25687 = n25663 & n25685;
  assign n25688 = ~n25686 & ~n25687;
  assign n25689 = n25674 & n25678;
  assign n25690 = n25684 & n25689;
  assign n25691 = n25688 & n25690;
  assign n25692 = n25670 & ~n25691;
  assign n25693 = ~n25608 & ~n25692;
  assign n25694 = n25608 & ~n25692;
  assign n25695 = ~n25693 & ~n25694;
  assign n25696 = ~n25511 & n25542;
  assign n25697 = ~n25417 & ~n25448;
  assign n25698 = n25480 & n25697;
  assign n25699 = n25696 & n25698;
  assign n25700 = n25639 & n25699;
  assign n25701 = n25695 & n25700;
  assign n25702 = ~n25573 & ~n25701;
  assign n25703 = ~n25542 & ~n25639;
  assign n25704 = ~n25511 & n25703;
  assign n25705 = n25576 & n25704;
  assign n25706 = ~n25693 & n25705;
  assign n25707 = ~n25694 & n25706;
  assign n25708 = n25573 & ~n25707;
  assign n25709 = ~n25702 & ~n25708;
  assign n25710 = n25653 & n25709;
  assign n25711 = ~P1_P3_FLUSH_REG & ~P1_P3_MORE_REG;
  assign n25712 = n25710 & ~n25711;
  assign n25713 = ~n25608 & n25639;
  assign n25714 = ~n25573 & n25713;
  assign n25715 = n25699 & n25714;
  assign n25716 = ~n25692 & n25715;
  assign n25717 = n25608 & n25639;
  assign n25718 = ~n25573 & n25717;
  assign n25719 = n25699 & n25718;
  assign n25720 = ~n25692 & n25719;
  assign n25721 = n25641 & ~n25692;
  assign n25722 = ~n25608 & ~n25639;
  assign n25723 = n25577 & n25722;
  assign n25724 = ~n25692 & n25723;
  assign n25725 = ~n25716 & ~n25720;
  assign n25726 = ~n25721 & n25725;
  assign n25727 = ~n25724 & n25726;
  assign n25728 = ~n25417 & n25448;
  assign n25729 = ~n25480 & n25728;
  assign n25730 = n25575 & n25729;
  assign n25731 = n25722 & n25730;
  assign n25732 = ~P1_P3_INSTQUEUERD_ADDR_REG_0_ & P1_P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n25733 = ~n25659 & ~n25732;
  assign n25734 = n25684 & n25733;
  assign n25735 = ~n25688 & ~n25734;
  assign n25736 = n25689 & ~n25735;
  assign n25737 = n25670 & ~n25736;
  assign n25738 = n25731 & ~n25737;
  assign n25739 = n25717 & n25730;
  assign n25740 = ~n25737 & n25739;
  assign n25741 = n25575 & n25698;
  assign n25742 = n25640 & n25741;
  assign n25743 = n25674 & ~n25735;
  assign n25744 = n25678 & n25743;
  assign n25745 = n25670 & ~n25744;
  assign n25746 = n25742 & ~n25745;
  assign n25747 = n25722 & n25741;
  assign n25748 = ~n25684 & ~n25733;
  assign n25749 = n25689 & ~n25748;
  assign n25750 = n25688 & n25749;
  assign n25751 = n25670 & ~n25750;
  assign n25752 = n25747 & ~n25751;
  assign n25753 = ~n25738 & ~n25740;
  assign n25754 = ~n25746 & n25753;
  assign n25755 = ~n25752 & n25754;
  assign n25756 = n25727 & n25755;
  assign n25757 = ~n25710 & ~n25756;
  assign n25758 = ~n25608 & ~n25751;
  assign n25759 = n25608 & ~n25745;
  assign n25760 = ~n25758 & ~n25759;
  assign n25761 = ~n25639 & n25741;
  assign n25762 = n25760 & n25761;
  assign n25763 = n25542 & n25573;
  assign n25764 = n25417 & ~n25448;
  assign n25765 = n25763 & n25764;
  assign n25766 = n25717 & n25765;
  assign n25767 = ~n25511 & n25766;
  assign n25768 = n25577 & ~n25639;
  assign n25769 = ~n25715 & ~n25767;
  assign n25770 = ~n25768 & n25769;
  assign n25771 = n25448 & n25542;
  assign n25772 = ~n25480 & n25573;
  assign n25773 = ~n25511 & n25717;
  assign n25774 = n25772 & n25773;
  assign n25775 = n25417 & ~n25573;
  assign n25776 = n25480 & n25511;
  assign n25777 = n25775 & n25776;
  assign n25778 = ~n25774 & ~n25777;
  assign n25779 = n25771 & ~n25778;
  assign n25780 = n25722 & n25776;
  assign n25781 = n25765 & n25780;
  assign n25782 = n25542 & ~n25573;
  assign n25783 = n25511 & n25713;
  assign n25784 = n25698 & n25782;
  assign n25785 = n25783 & n25784;
  assign n25786 = ~n25608 & n25741;
  assign n25787 = ~n25785 & ~n25786;
  assign n25788 = ~n25779 & ~n25781;
  assign n25789 = n25787 & n25788;
  assign n25790 = n25448 & ~n25511;
  assign n25791 = ~n25764 & ~n25790;
  assign n25792 = n25542 & n25791;
  assign n25793 = ~n25573 & ~n25792;
  assign n25794 = ~n25511 & ~n25764;
  assign n25795 = ~n25728 & n25794;
  assign n25796 = ~n25542 & n25795;
  assign n25797 = n25640 & ~n25796;
  assign n25798 = n25697 & n25717;
  assign n25799 = n25417 & n25511;
  assign n25800 = ~n25574 & ~n25799;
  assign n25801 = ~n25608 & n25800;
  assign n25802 = n25448 & n25480;
  assign n25803 = n25639 & n25802;
  assign n25804 = ~n25798 & ~n25801;
  assign n25805 = ~n25803 & n25804;
  assign n25806 = ~n25797 & n25805;
  assign n25807 = n25573 & ~n25806;
  assign n25808 = ~n25542 & ~n25802;
  assign n25809 = n25417 & n25808;
  assign n25810 = n25511 & n25608;
  assign n25811 = n25639 & ~n25810;
  assign n25812 = n25542 & ~n25811;
  assign n25813 = ~n25417 & n25812;
  assign n25814 = ~n25511 & ~n25697;
  assign n25815 = ~n25640 & n25814;
  assign n25816 = ~n25480 & ~n25815;
  assign n25817 = n25448 & ~n25608;
  assign n25818 = n25511 & n25817;
  assign n25819 = n25480 & ~n25608;
  assign n25820 = n25728 & n25819;
  assign n25821 = ~n25697 & n25713;
  assign n25822 = ~n25818 & ~n25820;
  assign n25823 = ~n25821 & n25822;
  assign n25824 = ~n25809 & ~n25813;
  assign n25825 = ~n25816 & n25824;
  assign n25826 = n25823 & n25825;
  assign n25827 = ~n25793 & ~n25807;
  assign n25828 = n25826 & n25827;
  assign n25829 = n25789 & n25828;
  assign n25830 = ~n25766 & n25829;
  assign n25831 = P1_P3_INSTQUEUERD_ADDR_REG_0_ & ~n25830;
  assign n25832 = n25770 & ~n25831;
  assign n25833 = ~P1_P3_INSTQUEUERD_ADDR_REG_2_ & ~n25832;
  assign n25834 = P1_P3_INSTQUEUERD_ADDR_REG_1_ & n25833;
  assign n25835 = P1_P3_INSTQUEUERD_ADDR_REG_2_ & ~n25770;
  assign n25836 = ~P1_P3_INSTQUEUERD_ADDR_REG_1_ & n25835;
  assign n25837 = ~P1_P3_INSTQUEUERD_ADDR_REG_2_ & P1_P3_INSTQUEUERD_ADDR_REG_1_;
  assign n25838 = P1_P3_INSTQUEUERD_ADDR_REG_2_ & ~P1_P3_INSTQUEUERD_ADDR_REG_1_;
  assign n25839 = ~n25837 & ~n25838;
  assign n25840 = n25719 & ~n25839;
  assign n25841 = P1_P3_INSTQUEUERD_ADDR_REG_2_ & ~n25360;
  assign n25842 = ~n25361 & ~n25841;
  assign n25843 = ~n25717 & ~n25722;
  assign n25844 = n25842 & ~n25843;
  assign n25845 = n25730 & n25844;
  assign n25846 = ~n25840 & ~n25845;
  assign n25847 = n25608 & n25771;
  assign n25848 = ~n25772 & ~n25777;
  assign n25849 = n25847 & ~n25848;
  assign n25850 = n25776 & ~n25843;
  assign n25851 = n25765 & n25850;
  assign n25852 = ~n25849 & ~n25851;
  assign n25853 = n25787 & n25852;
  assign n25854 = n25828 & n25853;
  assign n25855 = n25841 & ~n25854;
  assign n25856 = n25846 & ~n25855;
  assign n25857 = ~n25834 & ~n25836;
  assign n25858 = n25856 & n25857;
  assign n25859 = n25480 & n25639;
  assign n25860 = ~n25542 & ~n25713;
  assign n25861 = n25794 & ~n25859;
  assign n25862 = n25860 & n25861;
  assign n25863 = ~n25820 & n25862;
  assign n25864 = n25573 & ~n25863;
  assign n25865 = ~n25573 & ~n25700;
  assign n25866 = n25640 & ~n25795;
  assign n25867 = ~n25864 & ~n25865;
  assign n25868 = ~n25866 & n25867;
  assign n25869 = n25737 & n25739;
  assign n25870 = n25692 & n25719;
  assign n25871 = n25692 & n25723;
  assign n25872 = ~n25870 & ~n25871;
  assign n25873 = ~n25267 & ~n25872;
  assign n25874 = ~n25869 & ~n25873;
  assign n25875 = n25731 & n25737;
  assign n25876 = ~n25728 & n25772;
  assign n25877 = ~n25875 & ~n25876;
  assign n25878 = n25692 & n25715;
  assign n25879 = n25641 & n25692;
  assign n25880 = ~n25878 & ~n25879;
  assign n25881 = n25644 & ~n25880;
  assign n25882 = n25877 & ~n25881;
  assign n25883 = n25868 & n25874;
  assign n25884 = n25882 & n25883;
  assign n25885 = ~n25858 & ~n25884;
  assign n25886 = P1_P3_INSTQUEUERD_ADDR_REG_2_ & n25884;
  assign n25887 = ~n25885 & ~n25886;
  assign n25888 = P1_P3_INSTQUEUERD_ADDR_REG_1_ & n25390;
  assign n25889 = ~n25832 & n25888;
  assign n25890 = P1_P3_INSTQUEUERD_ADDR_REG_2_ & n25360;
  assign n25891 = P1_P3_INSTQUEUERD_ADDR_REG_3_ & ~n25890;
  assign n25892 = ~n25853 & n25891;
  assign n25893 = P1_P3_INSTQUEUERD_ADDR_REG_2_ & P1_P3_INSTQUEUERD_ADDR_REG_1_;
  assign n25894 = ~P1_P3_INSTQUEUERD_ADDR_REG_3_ & n25893;
  assign n25895 = P1_P3_INSTQUEUERD_ADDR_REG_3_ & ~n25893;
  assign n25896 = ~n25894 & ~n25895;
  assign n25897 = n25719 & ~n25896;
  assign n25898 = ~n25892 & ~n25897;
  assign n25899 = ~n25480 & n25767;
  assign n25900 = n25480 & n25767;
  assign n25901 = ~n25641 & ~n25723;
  assign n25902 = ~n25715 & n25901;
  assign n25903 = ~n25899 & ~n25900;
  assign n25904 = n25902 & n25903;
  assign n25905 = n25828 & n25904;
  assign n25906 = n25895 & ~n25905;
  assign n25907 = P1_P3_INSTQUEUERD_ADDR_REG_3_ & ~P1_P3_INSTQUEUERD_ADDR_REG_0_;
  assign n25908 = ~n25828 & n25907;
  assign n25909 = ~n25360 & n25404;
  assign n25910 = ~P1_P3_INSTQUEUERD_ADDR_REG_2_ & ~n25360;
  assign n25911 = P1_P3_INSTQUEUERD_ADDR_REG_3_ & ~n25910;
  assign n25912 = ~n25909 & ~n25911;
  assign n25913 = ~n25843 & n25912;
  assign n25914 = n25730 & n25913;
  assign n25915 = ~n25908 & ~n25914;
  assign n25916 = n25898 & ~n25906;
  assign n25917 = n25915 & n25916;
  assign n25918 = ~n25889 & n25917;
  assign n25919 = ~n25884 & ~n25918;
  assign n25920 = P1_P3_INSTQUEUERD_ADDR_REG_3_ & n25884;
  assign n25921 = ~n25919 & ~n25920;
  assign n25922 = ~n25887 & ~n25921;
  assign n25923 = P1_P3_INSTQUEUERD_ADDR_REG_4_ & n25884;
  assign n25924 = P1_P3_INSTQUEUERD_ADDR_REG_3_ & n25893;
  assign n25925 = ~P1_P3_INSTQUEUERD_ADDR_REG_4_ & n25924;
  assign n25926 = P1_P3_INSTQUEUERD_ADDR_REG_4_ & ~n25924;
  assign n25927 = ~n25925 & ~n25926;
  assign n25928 = n25719 & ~n25927;
  assign n25929 = ~n25884 & n25928;
  assign n25930 = ~n25923 & ~n25929;
  assign n25931 = ~n25922 & n25930;
  assign n25932 = ~P1_P3_INSTQUEUEWR_ADDR_REG_3_ & ~n25921;
  assign n25933 = ~P1_P3_INSTQUEUEWR_ADDR_REG_4_ & ~n25930;
  assign n25934 = P1_P3_INSTQUEUEWR_ADDR_REG_2_ & n25887;
  assign n25935 = P1_P3_INSTQUEUEWR_ADDR_REG_3_ & n25921;
  assign n25936 = n25728 & n25774;
  assign n25937 = ~n25731 & ~n25936;
  assign n25938 = n25766 & n25776;
  assign n25939 = n25829 & ~n25938;
  assign n25940 = n25937 & n25939;
  assign n25941 = ~P1_P3_INSTQUEUERD_ADDR_REG_0_ & ~n25940;
  assign n25942 = P1_P3_INSTQUEUERD_ADDR_REG_0_ & ~n25770;
  assign n25943 = P1_P3_INSTQUEUERD_ADDR_REG_0_ & n25719;
  assign n25944 = ~n25941 & ~n25942;
  assign n25945 = ~n25943 & n25944;
  assign n25946 = ~n25884 & ~n25945;
  assign n25947 = P1_P3_INSTQUEUERD_ADDR_REG_0_ & n25884;
  assign n25948 = ~n25946 & ~n25947;
  assign n25949 = P1_P3_INSTQUEUEWR_ADDR_REG_0_ & n25948;
  assign n25950 = ~P1_P3_INSTQUEUEWR_ADDR_REG_1_ & ~n25949;
  assign n25951 = ~P1_P3_INSTQUEUEWR_ADDR_REG_2_ & ~n25887;
  assign n25952 = ~P1_P3_INSTQUEUERD_ADDR_REG_1_ & ~n25832;
  assign n25953 = ~P1_P3_INSTQUEUERD_ADDR_REG_1_ & n25719;
  assign n25954 = ~n25360 & ~n25373;
  assign n25955 = ~n25937 & n25954;
  assign n25956 = ~n25953 & ~n25955;
  assign n25957 = n25364 & ~n25939;
  assign n25958 = n25956 & ~n25957;
  assign n25959 = ~n25952 & n25958;
  assign n25960 = ~n25884 & ~n25959;
  assign n25961 = P1_P3_INSTQUEUERD_ADDR_REG_1_ & n25884;
  assign n25962 = ~n25960 & ~n25961;
  assign n25963 = P1_P3_INSTQUEUEWR_ADDR_REG_1_ & n25949;
  assign n25964 = ~n25962 & ~n25963;
  assign n25965 = ~n25950 & ~n25951;
  assign n25966 = ~n25964 & n25965;
  assign n25967 = ~n25934 & ~n25935;
  assign n25968 = ~n25966 & n25967;
  assign n25969 = ~n25932 & ~n25933;
  assign n25970 = ~n25968 & n25969;
  assign n25971 = P1_P3_INSTQUEUEWR_ADDR_REG_4_ & n25930;
  assign n25972 = ~n25970 & ~n25971;
  assign n25973 = ~n25712 & ~n25757;
  assign n25974 = ~n25762 & n25973;
  assign n25975 = n25931 & n25974;
  assign n25976 = ~n25972 & n25975;
  assign n25977 = n25643 & n25976;
  assign n25978 = P1_P3_STATE2_REG_0_ & ~n25977;
  assign n25979 = ~n25354 & ~n25978;
  assign n25980 = P1_P3_STATE2_REG_2_ & n25979;
  assign n25981 = P1_P3_STATE2_REG_0_ & ~n25980;
  assign n25982 = n25352 & n25981;
  assign n25983 = P1_P3_STATE2_REG_3_ & ~n25981;
  assign n3596 = n25982 | n25983;
  assign n25985 = ~P1_P3_STATE2_REG_2_ & ~n25267;
  assign n25986 = P1_P3_STATE2_REG_0_ & ~n25985;
  assign n25987 = ~P1_P3_STATE2_REG_0_ & ~P1_P3_STATEBS16_REG;
  assign n25988 = ~n25986 & ~n25987;
  assign n25989 = P1_P3_STATE2_REG_1_ & n25988;
  assign n25990 = P1_P3_STATE2_REG_2_ & ~P1_P3_STATE2_REG_1_;
  assign n25991 = ~n25989 & ~n25990;
  assign n25992 = P1_P3_STATE2_REG_2_ & ~n25981;
  assign n3601 = ~n25991 | n25992;
  assign n25994 = P1_P3_STATE2_REG_0_ & n25990;
  assign n25995 = ~n25980 & n25994;
  assign n25996 = ~P1_P3_STATE2_REG_2_ & P1_P3_STATE2_REG_0_;
  assign n25997 = n25267 & n25996;
  assign n25998 = ~n25980 & ~n25997;
  assign n25999 = P1_P3_STATE2_REG_1_ & ~n25998;
  assign n26000 = ~P1_P3_STATE2_REG_3_ & ~P1_P3_STATE2_REG_1_;
  assign n26001 = ~n25267 & n26000;
  assign n26002 = n25981 & n26001;
  assign n26003 = P1_P3_STATE2_REG_1_ & ~P1_P3_STATE2_REG_0_;
  assign n26004 = ~P1_P3_STATE2_REG_2_ & n26003;
  assign n26005 = ~P1_P3_STATEBS16_REG & n26004;
  assign n26006 = ~n25995 & ~n25999;
  assign n26007 = ~n26002 & n26006;
  assign n3606 = n26005 | ~n26007;
  assign n26009 = P1_P3_STATE2_REG_3_ & ~P1_P3_INSTQUEUERD_ADDR_REG_4_;
  assign n26010 = ~P1_P3_STATE2_REG_2_ & ~P1_P3_STATE2_REG_1_;
  assign n26011 = n26009 & n26010;
  assign n26012 = ~n25980 & ~n26011;
  assign n26013 = ~P1_P3_STATE2_REG_0_ & n26012;
  assign n26014 = P1_P3_INSTADDRPOINTER_REG_0_ & P1_P3_INSTADDRPOINTER_REG_31_;
  assign n26015 = P1_P3_INSTADDRPOINTER_REG_0_ & ~P1_P3_INSTADDRPOINTER_REG_31_;
  assign n26016 = ~n26014 & ~n26015;
  assign n26017 = P1_P3_FLUSH_REG & n26016;
  assign n26018 = P1_P3_INSTQUEUERD_ADDR_REG_0_ & ~P1_P3_FLUSH_REG;
  assign n26019 = ~n26017 & ~n26018;
  assign n26020 = P1_P3_INSTADDRPOINTER_REG_0_ & ~P1_P3_INSTADDRPOINTER_REG_1_;
  assign n26021 = ~P1_P3_INSTADDRPOINTER_REG_0_ & P1_P3_INSTADDRPOINTER_REG_1_;
  assign n26022 = ~n26020 & ~n26021;
  assign n26023 = P1_P3_INSTADDRPOINTER_REG_31_ & ~n26022;
  assign n26024 = P1_P3_INSTADDRPOINTER_REG_1_ & ~P1_P3_INSTADDRPOINTER_REG_31_;
  assign n26025 = ~n26023 & ~n26024;
  assign n26026 = ~n26016 & n26025;
  assign n26027 = P1_P3_FLUSH_REG & n26026;
  assign n26028 = P1_P3_INSTQUEUERD_ADDR_REG_1_ & ~P1_P3_FLUSH_REG;
  assign n26029 = ~n26027 & ~n26028;
  assign n26030 = n26019 & n26029;
  assign n26031 = P1_P3_INSTQUEUERD_ADDR_REG_3_ & ~P1_P3_FLUSH_REG;
  assign n26032 = ~n26016 & ~n26025;
  assign n26033 = P1_P3_FLUSH_REG & n26032;
  assign n26034 = P1_P3_INSTQUEUERD_ADDR_REG_2_ & ~P1_P3_FLUSH_REG;
  assign n26035 = ~n26033 & ~n26034;
  assign n26036 = ~n26030 & n26031;
  assign n26037 = ~n26035 & n26036;
  assign n26038 = P1_P3_INSTQUEUERD_ADDR_REG_4_ & ~P1_P3_FLUSH_REG;
  assign n26039 = ~n26037 & ~n26038;
  assign n26040 = n25352 & n26039;
  assign n26041 = ~n25980 & ~n26040;
  assign n26042 = P1_P3_STATE2_REG_0_ & ~n26041;
  assign n26043 = P1_P3_STATE2_REG_3_ & P1_P3_STATE2_REG_0_;
  assign n26044 = n26010 & n26043;
  assign n26045 = ~n25997 & ~n26044;
  assign n26046 = ~n25976 & n25994;
  assign n26047 = n26045 & ~n26046;
  assign n26048 = ~n26013 & ~n26042;
  assign n3611 = ~n26047 | ~n26048;
  assign n26050 = P1_P3_INSTQUEUEWR_ADDR_REG_1_ & P1_P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n26051 = P1_P3_INSTQUEUEWR_ADDR_REG_2_ & n26050;
  assign n26052 = P1_P3_INSTQUEUEWR_ADDR_REG_3_ & n26051;
  assign n26053 = P1_P3_STATE2_REG_3_ & ~n26052;
  assign n26054 = ~P1_P3_STATE2_REG_2_ & P1_P3_STATE2_REG_1_;
  assign n26055 = ~n25990 & ~n26054;
  assign n26056 = ~n26009 & n26055;
  assign n26057 = ~P1_P3_STATE2_REG_0_ & ~n26056;
  assign n26058 = ~n26053 & n26057;
  assign n26059 = ~P1_P3_INSTQUEUEWR_ADDR_REG_2_ & n26050;
  assign n26060 = P1_P3_INSTQUEUEWR_ADDR_REG_2_ & ~n26050;
  assign n26061 = ~n26059 & ~n26060;
  assign n26062 = ~P1_P3_INSTQUEUEWR_ADDR_REG_3_ & n26051;
  assign n26063 = P1_P3_INSTQUEUEWR_ADDR_REG_3_ & ~n26051;
  assign n26064 = ~n26062 & ~n26063;
  assign n26065 = ~n26061 & ~n26064;
  assign n26066 = ~P1_P3_INSTQUEUEWR_ADDR_REG_1_ & P1_P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n26067 = P1_P3_INSTQUEUEWR_ADDR_REG_1_ & ~P1_P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n26068 = ~n26066 & ~n26067;
  assign n26069 = ~P1_P3_INSTQUEUEWR_ADDR_REG_0_ & ~n26068;
  assign n26070 = n26065 & n26069;
  assign n26071 = ~n26052 & ~n26070;
  assign n26072 = ~P1_P3_STATE2_REG_3_ & ~P1_P3_STATE2_REG_2_;
  assign n26073 = ~P1_P3_STATEBS16_REG & n26072;
  assign n26074 = ~P1_P3_STATE2_REG_2_ & ~n26073;
  assign n26075 = P1_P3_INSTQUEUEWR_ADDR_REG_0_ & ~n26068;
  assign n26076 = ~P1_P3_INSTQUEUEWR_ADDR_REG_0_ & n26068;
  assign n26077 = ~n26075 & ~n26076;
  assign n26078 = ~P1_P3_INSTQUEUEWR_ADDR_REG_0_ & ~n26077;
  assign n26079 = P1_P3_INSTQUEUEWR_ADDR_REG_0_ & n26077;
  assign n26080 = ~n26078 & ~n26079;
  assign n26081 = ~P1_P3_INSTQUEUEWR_ADDR_REG_0_ & ~n26080;
  assign n26082 = ~n26061 & ~n26069;
  assign n26083 = n26061 & n26069;
  assign n26084 = ~n26082 & ~n26083;
  assign n26085 = P1_P3_INSTQUEUEWR_ADDR_REG_0_ & ~n26077;
  assign n26086 = ~n26084 & ~n26085;
  assign n26087 = n26084 & n26085;
  assign n26088 = ~n26086 & ~n26087;
  assign n26089 = ~n26061 & n26064;
  assign n26090 = n26069 & n26089;
  assign n26091 = ~n26061 & n26069;
  assign n26092 = ~n26064 & ~n26091;
  assign n26093 = ~n26090 & ~n26092;
  assign n26094 = n26084 & ~n26093;
  assign n26095 = ~n26085 & ~n26093;
  assign n26096 = ~n26094 & ~n26095;
  assign n26097 = ~n26084 & n26093;
  assign n26098 = n26085 & n26097;
  assign n26099 = n26096 & ~n26098;
  assign n26100 = ~n26088 & ~n26099;
  assign n26101 = n26081 & n26100;
  assign n26102 = ~n26084 & ~n26093;
  assign n26103 = n26085 & n26102;
  assign n26104 = ~n26101 & ~n26103;
  assign n26105 = n26074 & ~n26104;
  assign n26106 = n26071 & ~n26105;
  assign n26107 = n26058 & ~n26106;
  assign n26108 = P1_P3_INSTQUEUE_REG_15__7_ & ~n26107;
  assign n26109 = P1_P3_STATEBS16_REG & n26072;
  assign n26110 = n26057 & n26109;
  assign n26111 = P1_BUF2_REG_23_ & n26110;
  assign n26112 = n26103 & n26111;
  assign n26113 = P1_P3_STATE2_REG_3_ & n26057;
  assign n26114 = ~n25511 & n26113;
  assign n26115 = n26052 & n26114;
  assign n26116 = ~n26112 & ~n26115;
  assign n26117 = P1_BUF2_REG_31_ & n26110;
  assign n26118 = n26101 & n26117;
  assign n26119 = n26116 & ~n26118;
  assign n26120 = n26104 & n26109;
  assign n26121 = n26074 & ~n26120;
  assign n26122 = ~n26071 & ~n26121;
  assign n26123 = P1_BUF2_REG_7_ & n26057;
  assign n26124 = n26122 & n26123;
  assign n26125 = ~n26108 & n26119;
  assign n3616 = n26124 | ~n26125;
  assign n26127 = P1_P3_INSTQUEUE_REG_15__6_ & ~n26107;
  assign n26128 = P1_BUF2_REG_22_ & n26110;
  assign n26129 = n26103 & n26128;
  assign n26130 = ~n25448 & n26113;
  assign n26131 = n26052 & n26130;
  assign n26132 = ~n26129 & ~n26131;
  assign n26133 = P1_BUF2_REG_30_ & n26110;
  assign n26134 = n26101 & n26133;
  assign n26135 = n26132 & ~n26134;
  assign n26136 = P1_BUF2_REG_6_ & n26057;
  assign n26137 = n26122 & n26136;
  assign n26138 = ~n26127 & n26135;
  assign n3621 = n26137 | ~n26138;
  assign n26140 = P1_P3_INSTQUEUE_REG_15__5_ & ~n26107;
  assign n26141 = P1_BUF2_REG_21_ & n26110;
  assign n26142 = n26103 & n26141;
  assign n26143 = ~n25417 & n26113;
  assign n26144 = n26052 & n26143;
  assign n26145 = ~n26142 & ~n26144;
  assign n26146 = P1_BUF2_REG_29_ & n26110;
  assign n26147 = n26101 & n26146;
  assign n26148 = n26145 & ~n26147;
  assign n26149 = P1_BUF2_REG_5_ & n26057;
  assign n26150 = n26122 & n26149;
  assign n26151 = ~n26140 & n26148;
  assign n3626 = n26150 | ~n26151;
  assign n26153 = P1_P3_INSTQUEUE_REG_15__4_ & ~n26107;
  assign n26154 = P1_BUF2_REG_20_ & n26110;
  assign n26155 = n26103 & n26154;
  assign n26156 = ~n25480 & n26113;
  assign n26157 = n26052 & n26156;
  assign n26158 = ~n26155 & ~n26157;
  assign n26159 = P1_BUF2_REG_28_ & n26110;
  assign n26160 = n26101 & n26159;
  assign n26161 = n26158 & ~n26160;
  assign n26162 = P1_BUF2_REG_4_ & n26057;
  assign n26163 = n26122 & n26162;
  assign n26164 = ~n26153 & n26161;
  assign n3631 = n26163 | ~n26164;
  assign n26166 = P1_P3_INSTQUEUE_REG_15__3_ & ~n26107;
  assign n26167 = P1_BUF2_REG_19_ & n26110;
  assign n26168 = n26103 & n26167;
  assign n26169 = ~n25542 & n26113;
  assign n26170 = n26052 & n26169;
  assign n26171 = ~n26168 & ~n26170;
  assign n26172 = P1_BUF2_REG_27_ & n26110;
  assign n26173 = n26101 & n26172;
  assign n26174 = n26171 & ~n26173;
  assign n26175 = P1_BUF2_REG_3_ & n26057;
  assign n26176 = n26122 & n26175;
  assign n26177 = ~n26166 & n26174;
  assign n3636 = n26176 | ~n26177;
  assign n26179 = P1_P3_INSTQUEUE_REG_15__2_ & ~n26107;
  assign n26180 = P1_BUF2_REG_18_ & n26110;
  assign n26181 = n26103 & n26180;
  assign n26182 = ~n25573 & n26113;
  assign n26183 = n26052 & n26182;
  assign n26184 = ~n26181 & ~n26183;
  assign n26185 = P1_BUF2_REG_26_ & n26110;
  assign n26186 = n26101 & n26185;
  assign n26187 = n26184 & ~n26186;
  assign n26188 = P1_BUF2_REG_2_ & n26057;
  assign n26189 = n26122 & n26188;
  assign n26190 = ~n26179 & n26187;
  assign n3641 = n26189 | ~n26190;
  assign n26192 = P1_P3_INSTQUEUE_REG_15__1_ & ~n26107;
  assign n26193 = P1_BUF2_REG_17_ & n26110;
  assign n26194 = n26103 & n26193;
  assign n26195 = ~n25608 & n26113;
  assign n26196 = n26052 & n26195;
  assign n26197 = ~n26194 & ~n26196;
  assign n26198 = P1_BUF2_REG_25_ & n26110;
  assign n26199 = n26101 & n26198;
  assign n26200 = n26197 & ~n26199;
  assign n26201 = P1_BUF2_REG_1_ & n26057;
  assign n26202 = n26122 & n26201;
  assign n26203 = ~n26192 & n26200;
  assign n3646 = n26202 | ~n26203;
  assign n26205 = P1_P3_INSTQUEUE_REG_15__0_ & ~n26107;
  assign n26206 = P1_BUF2_REG_16_ & n26110;
  assign n26207 = n26103 & n26206;
  assign n26208 = ~n25639 & n26113;
  assign n26209 = n26052 & n26208;
  assign n26210 = ~n26207 & ~n26209;
  assign n26211 = P1_BUF2_REG_24_ & n26110;
  assign n26212 = n26101 & n26211;
  assign n26213 = n26210 & ~n26212;
  assign n26214 = P1_BUF2_REG_0_ & n26057;
  assign n26215 = n26122 & n26214;
  assign n26216 = ~n26205 & n26213;
  assign n3651 = n26215 | ~n26216;
  assign n26218 = P1_P3_INSTQUEUEWR_ADDR_REG_3_ & P1_P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n26219 = P1_P3_INSTQUEUEWR_ADDR_REG_2_ & ~P1_P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n26220 = n26218 & n26219;
  assign n26221 = P1_P3_STATE2_REG_3_ & ~n26220;
  assign n26222 = n26057 & ~n26221;
  assign n26223 = n26065 & n26075;
  assign n26224 = ~n26220 & ~n26223;
  assign n26225 = P1_P3_INSTQUEUEWR_ADDR_REG_0_ & ~n26080;
  assign n26226 = n26100 & n26225;
  assign n26227 = n26078 & n26102;
  assign n26228 = ~n26226 & ~n26227;
  assign n26229 = n26074 & ~n26228;
  assign n26230 = n26224 & ~n26229;
  assign n26231 = n26222 & ~n26230;
  assign n26232 = P1_P3_INSTQUEUE_REG_14__7_ & ~n26231;
  assign n26233 = n26111 & n26227;
  assign n26234 = n26114 & n26220;
  assign n26235 = ~n26233 & ~n26234;
  assign n26236 = n26117 & n26226;
  assign n26237 = n26235 & ~n26236;
  assign n26238 = n26109 & n26228;
  assign n26239 = n26074 & ~n26238;
  assign n26240 = ~n26224 & ~n26239;
  assign n26241 = n26123 & n26240;
  assign n26242 = ~n26232 & n26237;
  assign n3656 = n26241 | ~n26242;
  assign n26244 = P1_P3_INSTQUEUE_REG_14__6_ & ~n26231;
  assign n26245 = n26128 & n26227;
  assign n26246 = n26130 & n26220;
  assign n26247 = ~n26245 & ~n26246;
  assign n26248 = n26133 & n26226;
  assign n26249 = n26247 & ~n26248;
  assign n26250 = n26136 & n26240;
  assign n26251 = ~n26244 & n26249;
  assign n3661 = n26250 | ~n26251;
  assign n26253 = P1_P3_INSTQUEUE_REG_14__5_ & ~n26231;
  assign n26254 = n26141 & n26227;
  assign n26255 = n26143 & n26220;
  assign n26256 = ~n26254 & ~n26255;
  assign n26257 = n26146 & n26226;
  assign n26258 = n26256 & ~n26257;
  assign n26259 = n26149 & n26240;
  assign n26260 = ~n26253 & n26258;
  assign n3666 = n26259 | ~n26260;
  assign n26262 = P1_P3_INSTQUEUE_REG_14__4_ & ~n26231;
  assign n26263 = n26154 & n26227;
  assign n26264 = n26156 & n26220;
  assign n26265 = ~n26263 & ~n26264;
  assign n26266 = n26159 & n26226;
  assign n26267 = n26265 & ~n26266;
  assign n26268 = n26162 & n26240;
  assign n26269 = ~n26262 & n26267;
  assign n3671 = n26268 | ~n26269;
  assign n26271 = P1_P3_INSTQUEUE_REG_14__3_ & ~n26231;
  assign n26272 = n26167 & n26227;
  assign n26273 = n26169 & n26220;
  assign n26274 = ~n26272 & ~n26273;
  assign n26275 = n26172 & n26226;
  assign n26276 = n26274 & ~n26275;
  assign n26277 = n26175 & n26240;
  assign n26278 = ~n26271 & n26276;
  assign n3676 = n26277 | ~n26278;
  assign n26280 = P1_P3_INSTQUEUE_REG_14__2_ & ~n26231;
  assign n26281 = n26180 & n26227;
  assign n26282 = n26182 & n26220;
  assign n26283 = ~n26281 & ~n26282;
  assign n26284 = n26185 & n26226;
  assign n26285 = n26283 & ~n26284;
  assign n26286 = n26188 & n26240;
  assign n26287 = ~n26280 & n26285;
  assign n3681 = n26286 | ~n26287;
  assign n26289 = P1_P3_INSTQUEUE_REG_14__1_ & ~n26231;
  assign n26290 = n26193 & n26227;
  assign n26291 = n26195 & n26220;
  assign n26292 = ~n26290 & ~n26291;
  assign n26293 = n26198 & n26226;
  assign n26294 = n26292 & ~n26293;
  assign n26295 = n26201 & n26240;
  assign n26296 = ~n26289 & n26294;
  assign n3686 = n26295 | ~n26296;
  assign n26298 = P1_P3_INSTQUEUE_REG_14__0_ & ~n26231;
  assign n26299 = n26206 & n26227;
  assign n26300 = n26208 & n26220;
  assign n26301 = ~n26299 & ~n26300;
  assign n26302 = n26211 & n26226;
  assign n26303 = n26301 & ~n26302;
  assign n26304 = n26214 & n26240;
  assign n26305 = ~n26298 & n26303;
  assign n3691 = n26304 | ~n26305;
  assign n26307 = P1_P3_INSTQUEUEWR_ADDR_REG_3_ & P1_P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n26308 = n26066 & n26307;
  assign n26309 = P1_P3_STATE2_REG_3_ & ~n26308;
  assign n26310 = n26057 & ~n26309;
  assign n26311 = n26065 & n26076;
  assign n26312 = ~n26308 & ~n26311;
  assign n26313 = ~P1_P3_INSTQUEUEWR_ADDR_REG_0_ & n26080;
  assign n26314 = n26100 & n26313;
  assign n26315 = n26079 & n26102;
  assign n26316 = ~n26314 & ~n26315;
  assign n26317 = n26074 & ~n26316;
  assign n26318 = n26312 & ~n26317;
  assign n26319 = n26310 & ~n26318;
  assign n26320 = P1_P3_INSTQUEUE_REG_13__7_ & ~n26319;
  assign n26321 = n26111 & n26315;
  assign n26322 = n26114 & n26308;
  assign n26323 = ~n26321 & ~n26322;
  assign n26324 = n26117 & n26314;
  assign n26325 = n26323 & ~n26324;
  assign n26326 = n26109 & n26316;
  assign n26327 = n26074 & ~n26326;
  assign n26328 = ~n26312 & ~n26327;
  assign n26329 = n26123 & n26328;
  assign n26330 = ~n26320 & n26325;
  assign n3696 = n26329 | ~n26330;
  assign n26332 = P1_P3_INSTQUEUE_REG_13__6_ & ~n26319;
  assign n26333 = n26128 & n26315;
  assign n26334 = n26130 & n26308;
  assign n26335 = ~n26333 & ~n26334;
  assign n26336 = n26133 & n26314;
  assign n26337 = n26335 & ~n26336;
  assign n26338 = n26136 & n26328;
  assign n26339 = ~n26332 & n26337;
  assign n3701 = n26338 | ~n26339;
  assign n26341 = P1_P3_INSTQUEUE_REG_13__5_ & ~n26319;
  assign n26342 = n26141 & n26315;
  assign n26343 = n26143 & n26308;
  assign n26344 = ~n26342 & ~n26343;
  assign n26345 = n26146 & n26314;
  assign n26346 = n26344 & ~n26345;
  assign n26347 = n26149 & n26328;
  assign n26348 = ~n26341 & n26346;
  assign n3706 = n26347 | ~n26348;
  assign n26350 = P1_P3_INSTQUEUE_REG_13__4_ & ~n26319;
  assign n26351 = n26154 & n26315;
  assign n26352 = n26156 & n26308;
  assign n26353 = ~n26351 & ~n26352;
  assign n26354 = n26159 & n26314;
  assign n26355 = n26353 & ~n26354;
  assign n26356 = n26162 & n26328;
  assign n26357 = ~n26350 & n26355;
  assign n3711 = n26356 | ~n26357;
  assign n26359 = P1_P3_INSTQUEUE_REG_13__3_ & ~n26319;
  assign n26360 = n26167 & n26315;
  assign n26361 = n26169 & n26308;
  assign n26362 = ~n26360 & ~n26361;
  assign n26363 = n26172 & n26314;
  assign n26364 = n26362 & ~n26363;
  assign n26365 = n26175 & n26328;
  assign n26366 = ~n26359 & n26364;
  assign n3716 = n26365 | ~n26366;
  assign n26368 = P1_P3_INSTQUEUE_REG_13__2_ & ~n26319;
  assign n26369 = n26180 & n26315;
  assign n26370 = n26182 & n26308;
  assign n26371 = ~n26369 & ~n26370;
  assign n26372 = n26185 & n26314;
  assign n26373 = n26371 & ~n26372;
  assign n26374 = n26188 & n26328;
  assign n26375 = ~n26368 & n26373;
  assign n3721 = n26374 | ~n26375;
  assign n26377 = P1_P3_INSTQUEUE_REG_13__1_ & ~n26319;
  assign n26378 = n26193 & n26315;
  assign n26379 = n26195 & n26308;
  assign n26380 = ~n26378 & ~n26379;
  assign n26381 = n26198 & n26314;
  assign n26382 = n26380 & ~n26381;
  assign n26383 = n26201 & n26328;
  assign n26384 = ~n26377 & n26382;
  assign n3726 = n26383 | ~n26384;
  assign n26386 = P1_P3_INSTQUEUE_REG_13__0_ & ~n26319;
  assign n26387 = n26206 & n26315;
  assign n26388 = n26208 & n26308;
  assign n26389 = ~n26387 & ~n26388;
  assign n26390 = n26211 & n26314;
  assign n26391 = n26389 & ~n26390;
  assign n26392 = n26214 & n26328;
  assign n26393 = ~n26386 & n26391;
  assign n3731 = n26392 | ~n26393;
  assign n26395 = P1_P3_INSTQUEUEWR_ADDR_REG_3_ & ~P1_P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n26396 = n26219 & n26395;
  assign n26397 = P1_P3_STATE2_REG_3_ & ~n26396;
  assign n26398 = n26057 & ~n26397;
  assign n26399 = P1_P3_INSTQUEUEWR_ADDR_REG_0_ & n26080;
  assign n26400 = n26100 & n26399;
  assign n26401 = ~P1_P3_INSTQUEUEWR_ADDR_REG_0_ & n26077;
  assign n26402 = n26102 & n26401;
  assign n26403 = ~n26400 & ~n26402;
  assign n26404 = n26074 & ~n26403;
  assign n26405 = n26065 & n26068;
  assign n26406 = ~n26404 & ~n26405;
  assign n26407 = n26398 & ~n26406;
  assign n26408 = P1_P3_INSTQUEUE_REG_12__7_ & ~n26407;
  assign n26409 = n26111 & n26402;
  assign n26410 = n26114 & n26396;
  assign n26411 = ~n26409 & ~n26410;
  assign n26412 = n26117 & n26400;
  assign n26413 = n26411 & ~n26412;
  assign n26414 = n26109 & n26403;
  assign n26415 = n26074 & ~n26414;
  assign n26416 = n26405 & ~n26415;
  assign n26417 = n26123 & n26416;
  assign n26418 = ~n26408 & n26413;
  assign n3736 = n26417 | ~n26418;
  assign n26420 = P1_P3_INSTQUEUE_REG_12__6_ & ~n26407;
  assign n26421 = n26128 & n26402;
  assign n26422 = n26130 & n26396;
  assign n26423 = ~n26421 & ~n26422;
  assign n26424 = n26133 & n26400;
  assign n26425 = n26423 & ~n26424;
  assign n26426 = n26136 & n26416;
  assign n26427 = ~n26420 & n26425;
  assign n3741 = n26426 | ~n26427;
  assign n26429 = P1_P3_INSTQUEUE_REG_12__5_ & ~n26407;
  assign n26430 = n26141 & n26402;
  assign n26431 = n26143 & n26396;
  assign n26432 = ~n26430 & ~n26431;
  assign n26433 = n26146 & n26400;
  assign n26434 = n26432 & ~n26433;
  assign n26435 = n26149 & n26416;
  assign n26436 = ~n26429 & n26434;
  assign n3746 = n26435 | ~n26436;
  assign n26438 = P1_P3_INSTQUEUE_REG_12__4_ & ~n26407;
  assign n26439 = n26154 & n26402;
  assign n26440 = n26156 & n26396;
  assign n26441 = ~n26439 & ~n26440;
  assign n26442 = n26159 & n26400;
  assign n26443 = n26441 & ~n26442;
  assign n26444 = n26162 & n26416;
  assign n26445 = ~n26438 & n26443;
  assign n3751 = n26444 | ~n26445;
  assign n26447 = P1_P3_INSTQUEUE_REG_12__3_ & ~n26407;
  assign n26448 = n26167 & n26402;
  assign n26449 = n26169 & n26396;
  assign n26450 = ~n26448 & ~n26449;
  assign n26451 = n26172 & n26400;
  assign n26452 = n26450 & ~n26451;
  assign n26453 = n26175 & n26416;
  assign n26454 = ~n26447 & n26452;
  assign n3756 = n26453 | ~n26454;
  assign n26456 = P1_P3_INSTQUEUE_REG_12__2_ & ~n26407;
  assign n26457 = n26180 & n26402;
  assign n26458 = n26182 & n26396;
  assign n26459 = ~n26457 & ~n26458;
  assign n26460 = n26185 & n26400;
  assign n26461 = n26459 & ~n26460;
  assign n26462 = n26188 & n26416;
  assign n26463 = ~n26456 & n26461;
  assign n3761 = n26462 | ~n26463;
  assign n26465 = P1_P3_INSTQUEUE_REG_12__1_ & ~n26407;
  assign n26466 = n26193 & n26402;
  assign n26467 = n26195 & n26396;
  assign n26468 = ~n26466 & ~n26467;
  assign n26469 = n26198 & n26400;
  assign n26470 = n26468 & ~n26469;
  assign n26471 = n26201 & n26416;
  assign n26472 = ~n26465 & n26470;
  assign n3766 = n26471 | ~n26472;
  assign n26474 = P1_P3_INSTQUEUE_REG_12__0_ & ~n26407;
  assign n26475 = n26206 & n26402;
  assign n26476 = n26208 & n26396;
  assign n26477 = ~n26475 & ~n26476;
  assign n26478 = n26211 & n26400;
  assign n26479 = n26477 & ~n26478;
  assign n26480 = n26214 & n26416;
  assign n26481 = ~n26474 & n26479;
  assign n3771 = n26480 | ~n26481;
  assign n26483 = P1_P3_INSTQUEUEWR_ADDR_REG_3_ & ~P1_P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n26484 = n26050 & n26483;
  assign n26485 = P1_P3_STATE2_REG_3_ & ~n26484;
  assign n26486 = n26057 & ~n26485;
  assign n26487 = n26061 & ~n26064;
  assign n26488 = n26069 & n26487;
  assign n26489 = ~n26484 & ~n26488;
  assign n26490 = n26088 & ~n26099;
  assign n26491 = n26081 & n26490;
  assign n26492 = n26085 & n26094;
  assign n26493 = ~n26491 & ~n26492;
  assign n26494 = n26074 & ~n26493;
  assign n26495 = n26489 & ~n26494;
  assign n26496 = n26486 & ~n26495;
  assign n26497 = P1_P3_INSTQUEUE_REG_11__7_ & ~n26496;
  assign n26498 = n26111 & n26492;
  assign n26499 = n26114 & n26484;
  assign n26500 = ~n26498 & ~n26499;
  assign n26501 = n26117 & n26491;
  assign n26502 = n26500 & ~n26501;
  assign n26503 = n26109 & n26493;
  assign n26504 = n26074 & ~n26503;
  assign n26505 = ~n26489 & ~n26504;
  assign n26506 = n26123 & n26505;
  assign n26507 = ~n26497 & n26502;
  assign n3776 = n26506 | ~n26507;
  assign n26509 = P1_P3_INSTQUEUE_REG_11__6_ & ~n26496;
  assign n26510 = n26128 & n26492;
  assign n26511 = n26130 & n26484;
  assign n26512 = ~n26510 & ~n26511;
  assign n26513 = n26133 & n26491;
  assign n26514 = n26512 & ~n26513;
  assign n26515 = n26136 & n26505;
  assign n26516 = ~n26509 & n26514;
  assign n3781 = n26515 | ~n26516;
  assign n26518 = P1_P3_INSTQUEUE_REG_11__5_ & ~n26496;
  assign n26519 = n26141 & n26492;
  assign n26520 = n26143 & n26484;
  assign n26521 = ~n26519 & ~n26520;
  assign n26522 = n26146 & n26491;
  assign n26523 = n26521 & ~n26522;
  assign n26524 = n26149 & n26505;
  assign n26525 = ~n26518 & n26523;
  assign n3786 = n26524 | ~n26525;
  assign n26527 = P1_P3_INSTQUEUE_REG_11__4_ & ~n26496;
  assign n26528 = n26154 & n26492;
  assign n26529 = n26156 & n26484;
  assign n26530 = ~n26528 & ~n26529;
  assign n26531 = n26159 & n26491;
  assign n26532 = n26530 & ~n26531;
  assign n26533 = n26162 & n26505;
  assign n26534 = ~n26527 & n26532;
  assign n3791 = n26533 | ~n26534;
  assign n26536 = P1_P3_INSTQUEUE_REG_11__3_ & ~n26496;
  assign n26537 = n26167 & n26492;
  assign n26538 = n26169 & n26484;
  assign n26539 = ~n26537 & ~n26538;
  assign n26540 = n26172 & n26491;
  assign n26541 = n26539 & ~n26540;
  assign n26542 = n26175 & n26505;
  assign n26543 = ~n26536 & n26541;
  assign n3796 = n26542 | ~n26543;
  assign n26545 = P1_P3_INSTQUEUE_REG_11__2_ & ~n26496;
  assign n26546 = n26180 & n26492;
  assign n26547 = n26182 & n26484;
  assign n26548 = ~n26546 & ~n26547;
  assign n26549 = n26185 & n26491;
  assign n26550 = n26548 & ~n26549;
  assign n26551 = n26188 & n26505;
  assign n26552 = ~n26545 & n26550;
  assign n3801 = n26551 | ~n26552;
  assign n26554 = P1_P3_INSTQUEUE_REG_11__1_ & ~n26496;
  assign n26555 = n26193 & n26492;
  assign n26556 = n26195 & n26484;
  assign n26557 = ~n26555 & ~n26556;
  assign n26558 = n26198 & n26491;
  assign n26559 = n26557 & ~n26558;
  assign n26560 = n26201 & n26505;
  assign n26561 = ~n26554 & n26559;
  assign n3806 = n26560 | ~n26561;
  assign n26563 = P1_P3_INSTQUEUE_REG_11__0_ & ~n26496;
  assign n26564 = n26206 & n26492;
  assign n26565 = n26208 & n26484;
  assign n26566 = ~n26564 & ~n26565;
  assign n26567 = n26211 & n26491;
  assign n26568 = n26566 & ~n26567;
  assign n26569 = n26214 & n26505;
  assign n26570 = ~n26563 & n26568;
  assign n3811 = n26569 | ~n26570;
  assign n26572 = ~P1_P3_INSTQUEUEWR_ADDR_REG_2_ & ~P1_P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n26573 = n26218 & n26572;
  assign n26574 = P1_P3_STATE2_REG_3_ & ~n26573;
  assign n26575 = n26057 & ~n26574;
  assign n26576 = n26075 & n26487;
  assign n26577 = ~n26573 & ~n26576;
  assign n26578 = n26225 & n26490;
  assign n26579 = n26078 & n26094;
  assign n26580 = ~n26578 & ~n26579;
  assign n26581 = n26074 & ~n26580;
  assign n26582 = n26577 & ~n26581;
  assign n26583 = n26575 & ~n26582;
  assign n26584 = P1_P3_INSTQUEUE_REG_10__7_ & ~n26583;
  assign n26585 = n26111 & n26579;
  assign n26586 = n26114 & n26573;
  assign n26587 = ~n26585 & ~n26586;
  assign n26588 = n26117 & n26578;
  assign n26589 = n26587 & ~n26588;
  assign n26590 = n26109 & n26580;
  assign n26591 = n26074 & ~n26590;
  assign n26592 = ~n26577 & ~n26591;
  assign n26593 = n26123 & n26592;
  assign n26594 = ~n26584 & n26589;
  assign n3816 = n26593 | ~n26594;
  assign n26596 = P1_P3_INSTQUEUE_REG_10__6_ & ~n26583;
  assign n26597 = n26128 & n26579;
  assign n26598 = n26130 & n26573;
  assign n26599 = ~n26597 & ~n26598;
  assign n26600 = n26133 & n26578;
  assign n26601 = n26599 & ~n26600;
  assign n26602 = n26136 & n26592;
  assign n26603 = ~n26596 & n26601;
  assign n3821 = n26602 | ~n26603;
  assign n26605 = P1_P3_INSTQUEUE_REG_10__5_ & ~n26583;
  assign n26606 = n26141 & n26579;
  assign n26607 = n26143 & n26573;
  assign n26608 = ~n26606 & ~n26607;
  assign n26609 = n26146 & n26578;
  assign n26610 = n26608 & ~n26609;
  assign n26611 = n26149 & n26592;
  assign n26612 = ~n26605 & n26610;
  assign n3826 = n26611 | ~n26612;
  assign n26614 = P1_P3_INSTQUEUE_REG_10__4_ & ~n26583;
  assign n26615 = n26154 & n26579;
  assign n26616 = n26156 & n26573;
  assign n26617 = ~n26615 & ~n26616;
  assign n26618 = n26159 & n26578;
  assign n26619 = n26617 & ~n26618;
  assign n26620 = n26162 & n26592;
  assign n26621 = ~n26614 & n26619;
  assign n3831 = n26620 | ~n26621;
  assign n26623 = P1_P3_INSTQUEUE_REG_10__3_ & ~n26583;
  assign n26624 = n26167 & n26579;
  assign n26625 = n26169 & n26573;
  assign n26626 = ~n26624 & ~n26625;
  assign n26627 = n26172 & n26578;
  assign n26628 = n26626 & ~n26627;
  assign n26629 = n26175 & n26592;
  assign n26630 = ~n26623 & n26628;
  assign n3836 = n26629 | ~n26630;
  assign n26632 = P1_P3_INSTQUEUE_REG_10__2_ & ~n26583;
  assign n26633 = n26180 & n26579;
  assign n26634 = n26182 & n26573;
  assign n26635 = ~n26633 & ~n26634;
  assign n26636 = n26185 & n26578;
  assign n26637 = n26635 & ~n26636;
  assign n26638 = n26188 & n26592;
  assign n26639 = ~n26632 & n26637;
  assign n3841 = n26638 | ~n26639;
  assign n26641 = P1_P3_INSTQUEUE_REG_10__1_ & ~n26583;
  assign n26642 = n26193 & n26579;
  assign n26643 = n26195 & n26573;
  assign n26644 = ~n26642 & ~n26643;
  assign n26645 = n26198 & n26578;
  assign n26646 = n26644 & ~n26645;
  assign n26647 = n26201 & n26592;
  assign n26648 = ~n26641 & n26646;
  assign n3846 = n26647 | ~n26648;
  assign n26650 = P1_P3_INSTQUEUE_REG_10__0_ & ~n26583;
  assign n26651 = n26206 & n26579;
  assign n26652 = n26208 & n26573;
  assign n26653 = ~n26651 & ~n26652;
  assign n26654 = n26211 & n26578;
  assign n26655 = n26653 & ~n26654;
  assign n26656 = n26214 & n26592;
  assign n26657 = ~n26650 & n26655;
  assign n3851 = n26656 | ~n26657;
  assign n26659 = n26066 & n26483;
  assign n26660 = P1_P3_STATE2_REG_3_ & ~n26659;
  assign n26661 = n26057 & ~n26660;
  assign n26662 = n26076 & n26487;
  assign n26663 = ~n26659 & ~n26662;
  assign n26664 = n26313 & n26490;
  assign n26665 = n26079 & n26094;
  assign n26666 = ~n26664 & ~n26665;
  assign n26667 = n26074 & ~n26666;
  assign n26668 = n26663 & ~n26667;
  assign n26669 = n26661 & ~n26668;
  assign n26670 = P1_P3_INSTQUEUE_REG_9__7_ & ~n26669;
  assign n26671 = n26111 & n26665;
  assign n26672 = n26114 & n26659;
  assign n26673 = ~n26671 & ~n26672;
  assign n26674 = n26117 & n26664;
  assign n26675 = n26673 & ~n26674;
  assign n26676 = n26109 & n26666;
  assign n26677 = n26074 & ~n26676;
  assign n26678 = ~n26663 & ~n26677;
  assign n26679 = n26123 & n26678;
  assign n26680 = ~n26670 & n26675;
  assign n3856 = n26679 | ~n26680;
  assign n26682 = P1_P3_INSTQUEUE_REG_9__6_ & ~n26669;
  assign n26683 = n26128 & n26665;
  assign n26684 = n26130 & n26659;
  assign n26685 = ~n26683 & ~n26684;
  assign n26686 = n26133 & n26664;
  assign n26687 = n26685 & ~n26686;
  assign n26688 = n26136 & n26678;
  assign n26689 = ~n26682 & n26687;
  assign n3861 = n26688 | ~n26689;
  assign n26691 = P1_P3_INSTQUEUE_REG_9__5_ & ~n26669;
  assign n26692 = n26141 & n26665;
  assign n26693 = n26143 & n26659;
  assign n26694 = ~n26692 & ~n26693;
  assign n26695 = n26146 & n26664;
  assign n26696 = n26694 & ~n26695;
  assign n26697 = n26149 & n26678;
  assign n26698 = ~n26691 & n26696;
  assign n3866 = n26697 | ~n26698;
  assign n26700 = P1_P3_INSTQUEUE_REG_9__4_ & ~n26669;
  assign n26701 = n26154 & n26665;
  assign n26702 = n26156 & n26659;
  assign n26703 = ~n26701 & ~n26702;
  assign n26704 = n26159 & n26664;
  assign n26705 = n26703 & ~n26704;
  assign n26706 = n26162 & n26678;
  assign n26707 = ~n26700 & n26705;
  assign n3871 = n26706 | ~n26707;
  assign n26709 = P1_P3_INSTQUEUE_REG_9__3_ & ~n26669;
  assign n26710 = n26167 & n26665;
  assign n26711 = n26169 & n26659;
  assign n26712 = ~n26710 & ~n26711;
  assign n26713 = n26172 & n26664;
  assign n26714 = n26712 & ~n26713;
  assign n26715 = n26175 & n26678;
  assign n26716 = ~n26709 & n26714;
  assign n3876 = n26715 | ~n26716;
  assign n26718 = P1_P3_INSTQUEUE_REG_9__2_ & ~n26669;
  assign n26719 = n26180 & n26665;
  assign n26720 = n26182 & n26659;
  assign n26721 = ~n26719 & ~n26720;
  assign n26722 = n26185 & n26664;
  assign n26723 = n26721 & ~n26722;
  assign n26724 = n26188 & n26678;
  assign n26725 = ~n26718 & n26723;
  assign n3881 = n26724 | ~n26725;
  assign n26727 = P1_P3_INSTQUEUE_REG_9__1_ & ~n26669;
  assign n26728 = n26193 & n26665;
  assign n26729 = n26195 & n26659;
  assign n26730 = ~n26728 & ~n26729;
  assign n26731 = n26198 & n26664;
  assign n26732 = n26730 & ~n26731;
  assign n26733 = n26201 & n26678;
  assign n26734 = ~n26727 & n26732;
  assign n3886 = n26733 | ~n26734;
  assign n26736 = P1_P3_INSTQUEUE_REG_9__0_ & ~n26669;
  assign n26737 = n26206 & n26665;
  assign n26738 = n26208 & n26659;
  assign n26739 = ~n26737 & ~n26738;
  assign n26740 = n26211 & n26664;
  assign n26741 = n26739 & ~n26740;
  assign n26742 = n26214 & n26678;
  assign n26743 = ~n26736 & n26741;
  assign n3891 = n26742 | ~n26743;
  assign n26745 = n26395 & n26572;
  assign n26746 = P1_P3_STATE2_REG_3_ & ~n26745;
  assign n26747 = n26057 & ~n26746;
  assign n26748 = n26399 & n26490;
  assign n26749 = n26094 & n26401;
  assign n26750 = ~n26748 & ~n26749;
  assign n26751 = n26074 & ~n26750;
  assign n26752 = n26068 & n26487;
  assign n26753 = ~n26751 & ~n26752;
  assign n26754 = n26747 & ~n26753;
  assign n26755 = P1_P3_INSTQUEUE_REG_8__7_ & ~n26754;
  assign n26756 = n26111 & n26749;
  assign n26757 = n26114 & n26745;
  assign n26758 = ~n26756 & ~n26757;
  assign n26759 = n26117 & n26748;
  assign n26760 = n26758 & ~n26759;
  assign n26761 = n26109 & n26750;
  assign n26762 = n26074 & ~n26761;
  assign n26763 = n26752 & ~n26762;
  assign n26764 = n26123 & n26763;
  assign n26765 = ~n26755 & n26760;
  assign n3896 = n26764 | ~n26765;
  assign n26767 = P1_P3_INSTQUEUE_REG_8__6_ & ~n26754;
  assign n26768 = n26128 & n26749;
  assign n26769 = n26130 & n26745;
  assign n26770 = ~n26768 & ~n26769;
  assign n26771 = n26133 & n26748;
  assign n26772 = n26770 & ~n26771;
  assign n26773 = n26136 & n26763;
  assign n26774 = ~n26767 & n26772;
  assign n3901 = n26773 | ~n26774;
  assign n26776 = P1_P3_INSTQUEUE_REG_8__5_ & ~n26754;
  assign n26777 = n26141 & n26749;
  assign n26778 = n26143 & n26745;
  assign n26779 = ~n26777 & ~n26778;
  assign n26780 = n26146 & n26748;
  assign n26781 = n26779 & ~n26780;
  assign n26782 = n26149 & n26763;
  assign n26783 = ~n26776 & n26781;
  assign n3906 = n26782 | ~n26783;
  assign n26785 = P1_P3_INSTQUEUE_REG_8__4_ & ~n26754;
  assign n26786 = n26154 & n26749;
  assign n26787 = n26156 & n26745;
  assign n26788 = ~n26786 & ~n26787;
  assign n26789 = n26159 & n26748;
  assign n26790 = n26788 & ~n26789;
  assign n26791 = n26162 & n26763;
  assign n26792 = ~n26785 & n26790;
  assign n3911 = n26791 | ~n26792;
  assign n26794 = P1_P3_INSTQUEUE_REG_8__3_ & ~n26754;
  assign n26795 = n26167 & n26749;
  assign n26796 = n26169 & n26745;
  assign n26797 = ~n26795 & ~n26796;
  assign n26798 = n26172 & n26748;
  assign n26799 = n26797 & ~n26798;
  assign n26800 = n26175 & n26763;
  assign n26801 = ~n26794 & n26799;
  assign n3916 = n26800 | ~n26801;
  assign n26803 = P1_P3_INSTQUEUE_REG_8__2_ & ~n26754;
  assign n26804 = n26180 & n26749;
  assign n26805 = n26182 & n26745;
  assign n26806 = ~n26804 & ~n26805;
  assign n26807 = n26185 & n26748;
  assign n26808 = n26806 & ~n26807;
  assign n26809 = n26188 & n26763;
  assign n26810 = ~n26803 & n26808;
  assign n3921 = n26809 | ~n26810;
  assign n26812 = P1_P3_INSTQUEUE_REG_8__1_ & ~n26754;
  assign n26813 = n26193 & n26749;
  assign n26814 = n26195 & n26745;
  assign n26815 = ~n26813 & ~n26814;
  assign n26816 = n26198 & n26748;
  assign n26817 = n26815 & ~n26816;
  assign n26818 = n26201 & n26763;
  assign n26819 = ~n26812 & n26817;
  assign n3926 = n26818 | ~n26819;
  assign n26821 = P1_P3_INSTQUEUE_REG_8__0_ & ~n26754;
  assign n26822 = n26206 & n26749;
  assign n26823 = n26208 & n26745;
  assign n26824 = ~n26822 & ~n26823;
  assign n26825 = n26211 & n26748;
  assign n26826 = n26824 & ~n26825;
  assign n26827 = n26214 & n26763;
  assign n26828 = ~n26821 & n26826;
  assign n3931 = n26827 | ~n26828;
  assign n26830 = P1_P3_STATE2_REG_3_ & ~n26062;
  assign n26831 = n26057 & ~n26830;
  assign n26832 = ~n26062 & ~n26090;
  assign n26833 = ~n26088 & n26099;
  assign n26834 = n26081 & n26833;
  assign n26835 = ~n26098 & ~n26834;
  assign n26836 = n26074 & ~n26835;
  assign n26837 = n26832 & ~n26836;
  assign n26838 = n26831 & ~n26837;
  assign n26839 = P1_P3_INSTQUEUE_REG_7__7_ & ~n26838;
  assign n26840 = n26098 & n26111;
  assign n26841 = n26062 & n26114;
  assign n26842 = ~n26840 & ~n26841;
  assign n26843 = n26117 & n26834;
  assign n26844 = n26842 & ~n26843;
  assign n26845 = n26109 & n26835;
  assign n26846 = n26074 & ~n26845;
  assign n26847 = ~n26832 & ~n26846;
  assign n26848 = n26123 & n26847;
  assign n26849 = ~n26839 & n26844;
  assign n3936 = n26848 | ~n26849;
  assign n26851 = P1_P3_INSTQUEUE_REG_7__6_ & ~n26838;
  assign n26852 = n26098 & n26128;
  assign n26853 = n26062 & n26130;
  assign n26854 = ~n26852 & ~n26853;
  assign n26855 = n26133 & n26834;
  assign n26856 = n26854 & ~n26855;
  assign n26857 = n26136 & n26847;
  assign n26858 = ~n26851 & n26856;
  assign n3941 = n26857 | ~n26858;
  assign n26860 = P1_P3_INSTQUEUE_REG_7__5_ & ~n26838;
  assign n26861 = n26098 & n26141;
  assign n26862 = n26062 & n26143;
  assign n26863 = ~n26861 & ~n26862;
  assign n26864 = n26146 & n26834;
  assign n26865 = n26863 & ~n26864;
  assign n26866 = n26149 & n26847;
  assign n26867 = ~n26860 & n26865;
  assign n3946 = n26866 | ~n26867;
  assign n26869 = P1_P3_INSTQUEUE_REG_7__4_ & ~n26838;
  assign n26870 = n26098 & n26154;
  assign n26871 = n26062 & n26156;
  assign n26872 = ~n26870 & ~n26871;
  assign n26873 = n26159 & n26834;
  assign n26874 = n26872 & ~n26873;
  assign n26875 = n26162 & n26847;
  assign n26876 = ~n26869 & n26874;
  assign n3951 = n26875 | ~n26876;
  assign n26878 = P1_P3_INSTQUEUE_REG_7__3_ & ~n26838;
  assign n26879 = n26098 & n26167;
  assign n26880 = n26062 & n26169;
  assign n26881 = ~n26879 & ~n26880;
  assign n26882 = n26172 & n26834;
  assign n26883 = n26881 & ~n26882;
  assign n26884 = n26175 & n26847;
  assign n26885 = ~n26878 & n26883;
  assign n3956 = n26884 | ~n26885;
  assign n26887 = P1_P3_INSTQUEUE_REG_7__2_ & ~n26838;
  assign n26888 = n26098 & n26180;
  assign n26889 = n26062 & n26182;
  assign n26890 = ~n26888 & ~n26889;
  assign n26891 = n26185 & n26834;
  assign n26892 = n26890 & ~n26891;
  assign n26893 = n26188 & n26847;
  assign n26894 = ~n26887 & n26892;
  assign n3961 = n26893 | ~n26894;
  assign n26896 = P1_P3_INSTQUEUE_REG_7__1_ & ~n26838;
  assign n26897 = n26098 & n26193;
  assign n26898 = n26062 & n26195;
  assign n26899 = ~n26897 & ~n26898;
  assign n26900 = n26198 & n26834;
  assign n26901 = n26899 & ~n26900;
  assign n26902 = n26201 & n26847;
  assign n26903 = ~n26896 & n26901;
  assign n3966 = n26902 | ~n26903;
  assign n26905 = P1_P3_INSTQUEUE_REG_7__0_ & ~n26838;
  assign n26906 = n26098 & n26206;
  assign n26907 = n26062 & n26208;
  assign n26908 = ~n26906 & ~n26907;
  assign n26909 = n26211 & n26834;
  assign n26910 = n26908 & ~n26909;
  assign n26911 = n26214 & n26847;
  assign n26912 = ~n26905 & n26910;
  assign n3971 = n26911 | ~n26912;
  assign n26914 = ~P1_P3_INSTQUEUEWR_ADDR_REG_3_ & P1_P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n26915 = n26219 & n26914;
  assign n26916 = P1_P3_STATE2_REG_3_ & ~n26915;
  assign n26917 = n26057 & ~n26916;
  assign n26918 = n26075 & n26089;
  assign n26919 = ~n26915 & ~n26918;
  assign n26920 = n26225 & n26833;
  assign n26921 = n26078 & n26097;
  assign n26922 = ~n26920 & ~n26921;
  assign n26923 = n26074 & ~n26922;
  assign n26924 = n26919 & ~n26923;
  assign n26925 = n26917 & ~n26924;
  assign n26926 = P1_P3_INSTQUEUE_REG_6__7_ & ~n26925;
  assign n26927 = n26111 & n26921;
  assign n26928 = n26114 & n26915;
  assign n26929 = ~n26927 & ~n26928;
  assign n26930 = n26117 & n26920;
  assign n26931 = n26929 & ~n26930;
  assign n26932 = n26109 & n26922;
  assign n26933 = n26074 & ~n26932;
  assign n26934 = ~n26919 & ~n26933;
  assign n26935 = n26123 & n26934;
  assign n26936 = ~n26926 & n26931;
  assign n3976 = n26935 | ~n26936;
  assign n26938 = P1_P3_INSTQUEUE_REG_6__6_ & ~n26925;
  assign n26939 = n26128 & n26921;
  assign n26940 = n26130 & n26915;
  assign n26941 = ~n26939 & ~n26940;
  assign n26942 = n26133 & n26920;
  assign n26943 = n26941 & ~n26942;
  assign n26944 = n26136 & n26934;
  assign n26945 = ~n26938 & n26943;
  assign n3981 = n26944 | ~n26945;
  assign n26947 = P1_P3_INSTQUEUE_REG_6__5_ & ~n26925;
  assign n26948 = n26141 & n26921;
  assign n26949 = n26143 & n26915;
  assign n26950 = ~n26948 & ~n26949;
  assign n26951 = n26146 & n26920;
  assign n26952 = n26950 & ~n26951;
  assign n26953 = n26149 & n26934;
  assign n26954 = ~n26947 & n26952;
  assign n3986 = n26953 | ~n26954;
  assign n26956 = P1_P3_INSTQUEUE_REG_6__4_ & ~n26925;
  assign n26957 = n26154 & n26921;
  assign n26958 = n26156 & n26915;
  assign n26959 = ~n26957 & ~n26958;
  assign n26960 = n26159 & n26920;
  assign n26961 = n26959 & ~n26960;
  assign n26962 = n26162 & n26934;
  assign n26963 = ~n26956 & n26961;
  assign n3991 = n26962 | ~n26963;
  assign n26965 = P1_P3_INSTQUEUE_REG_6__3_ & ~n26925;
  assign n26966 = n26167 & n26921;
  assign n26967 = n26169 & n26915;
  assign n26968 = ~n26966 & ~n26967;
  assign n26969 = n26172 & n26920;
  assign n26970 = n26968 & ~n26969;
  assign n26971 = n26175 & n26934;
  assign n26972 = ~n26965 & n26970;
  assign n3996 = n26971 | ~n26972;
  assign n26974 = P1_P3_INSTQUEUE_REG_6__2_ & ~n26925;
  assign n26975 = n26180 & n26921;
  assign n26976 = n26182 & n26915;
  assign n26977 = ~n26975 & ~n26976;
  assign n26978 = n26185 & n26920;
  assign n26979 = n26977 & ~n26978;
  assign n26980 = n26188 & n26934;
  assign n26981 = ~n26974 & n26979;
  assign n4001 = n26980 | ~n26981;
  assign n26983 = P1_P3_INSTQUEUE_REG_6__1_ & ~n26925;
  assign n26984 = n26193 & n26921;
  assign n26985 = n26195 & n26915;
  assign n26986 = ~n26984 & ~n26985;
  assign n26987 = n26198 & n26920;
  assign n26988 = n26986 & ~n26987;
  assign n26989 = n26201 & n26934;
  assign n26990 = ~n26983 & n26988;
  assign n4006 = n26989 | ~n26990;
  assign n26992 = P1_P3_INSTQUEUE_REG_6__0_ & ~n26925;
  assign n26993 = n26206 & n26921;
  assign n26994 = n26208 & n26915;
  assign n26995 = ~n26993 & ~n26994;
  assign n26996 = n26211 & n26920;
  assign n26997 = n26995 & ~n26996;
  assign n26998 = n26214 & n26934;
  assign n26999 = ~n26992 & n26997;
  assign n4011 = n26998 | ~n26999;
  assign n27001 = ~P1_P3_INSTQUEUEWR_ADDR_REG_3_ & P1_P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n27002 = n26066 & n27001;
  assign n27003 = P1_P3_STATE2_REG_3_ & ~n27002;
  assign n27004 = n26057 & ~n27003;
  assign n27005 = n26076 & n26089;
  assign n27006 = ~n27002 & ~n27005;
  assign n27007 = n26313 & n26833;
  assign n27008 = n26079 & n26097;
  assign n27009 = ~n27007 & ~n27008;
  assign n27010 = n26074 & ~n27009;
  assign n27011 = n27006 & ~n27010;
  assign n27012 = n27004 & ~n27011;
  assign n27013 = P1_P3_INSTQUEUE_REG_5__7_ & ~n27012;
  assign n27014 = n26111 & n27008;
  assign n27015 = n26114 & n27002;
  assign n27016 = ~n27014 & ~n27015;
  assign n27017 = n26117 & n27007;
  assign n27018 = n27016 & ~n27017;
  assign n27019 = n26109 & n27009;
  assign n27020 = n26074 & ~n27019;
  assign n27021 = ~n27006 & ~n27020;
  assign n27022 = n26123 & n27021;
  assign n27023 = ~n27013 & n27018;
  assign n4016 = n27022 | ~n27023;
  assign n27025 = P1_P3_INSTQUEUE_REG_5__6_ & ~n27012;
  assign n27026 = n26128 & n27008;
  assign n27027 = n26130 & n27002;
  assign n27028 = ~n27026 & ~n27027;
  assign n27029 = n26133 & n27007;
  assign n27030 = n27028 & ~n27029;
  assign n27031 = n26136 & n27021;
  assign n27032 = ~n27025 & n27030;
  assign n4021 = n27031 | ~n27032;
  assign n27034 = P1_P3_INSTQUEUE_REG_5__5_ & ~n27012;
  assign n27035 = n26141 & n27008;
  assign n27036 = n26143 & n27002;
  assign n27037 = ~n27035 & ~n27036;
  assign n27038 = n26146 & n27007;
  assign n27039 = n27037 & ~n27038;
  assign n27040 = n26149 & n27021;
  assign n27041 = ~n27034 & n27039;
  assign n4026 = n27040 | ~n27041;
  assign n27043 = P1_P3_INSTQUEUE_REG_5__4_ & ~n27012;
  assign n27044 = n26154 & n27008;
  assign n27045 = n26156 & n27002;
  assign n27046 = ~n27044 & ~n27045;
  assign n27047 = n26159 & n27007;
  assign n27048 = n27046 & ~n27047;
  assign n27049 = n26162 & n27021;
  assign n27050 = ~n27043 & n27048;
  assign n4031 = n27049 | ~n27050;
  assign n27052 = P1_P3_INSTQUEUE_REG_5__3_ & ~n27012;
  assign n27053 = n26167 & n27008;
  assign n27054 = n26169 & n27002;
  assign n27055 = ~n27053 & ~n27054;
  assign n27056 = n26172 & n27007;
  assign n27057 = n27055 & ~n27056;
  assign n27058 = n26175 & n27021;
  assign n27059 = ~n27052 & n27057;
  assign n4036 = n27058 | ~n27059;
  assign n27061 = P1_P3_INSTQUEUE_REG_5__2_ & ~n27012;
  assign n27062 = n26180 & n27008;
  assign n27063 = n26182 & n27002;
  assign n27064 = ~n27062 & ~n27063;
  assign n27065 = n26185 & n27007;
  assign n27066 = n27064 & ~n27065;
  assign n27067 = n26188 & n27021;
  assign n27068 = ~n27061 & n27066;
  assign n4041 = n27067 | ~n27068;
  assign n27070 = P1_P3_INSTQUEUE_REG_5__1_ & ~n27012;
  assign n27071 = n26193 & n27008;
  assign n27072 = n26195 & n27002;
  assign n27073 = ~n27071 & ~n27072;
  assign n27074 = n26198 & n27007;
  assign n27075 = n27073 & ~n27074;
  assign n27076 = n26201 & n27021;
  assign n27077 = ~n27070 & n27075;
  assign n4046 = n27076 | ~n27077;
  assign n27079 = P1_P3_INSTQUEUE_REG_5__0_ & ~n27012;
  assign n27080 = n26206 & n27008;
  assign n27081 = n26208 & n27002;
  assign n27082 = ~n27080 & ~n27081;
  assign n27083 = n26211 & n27007;
  assign n27084 = n27082 & ~n27083;
  assign n27085 = n26214 & n27021;
  assign n27086 = ~n27079 & n27084;
  assign n4051 = n27085 | ~n27086;
  assign n27088 = n26097 & n26401;
  assign n27089 = n26111 & n27088;
  assign n27090 = ~P1_P3_INSTQUEUEWR_ADDR_REG_3_ & ~P1_P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n27091 = n26219 & n27090;
  assign n27092 = n26114 & n27091;
  assign n27093 = n26074 & ~n26109;
  assign n27094 = n26068 & n26089;
  assign n27095 = ~n27093 & n27094;
  assign n27096 = n26123 & n27095;
  assign n27097 = ~n27089 & ~n27092;
  assign n27098 = ~n27096 & n27097;
  assign n27099 = n26399 & n26833;
  assign n27100 = n26117 & n27099;
  assign n27101 = n27098 & ~n27100;
  assign n27102 = P1_P3_STATE2_REG_3_ & ~n27091;
  assign n27103 = n26057 & ~n27102;
  assign n27104 = ~n27088 & ~n27099;
  assign n27105 = n26074 & ~n27104;
  assign n27106 = ~n27094 & ~n27105;
  assign n27107 = n27103 & ~n27106;
  assign n27108 = P1_P3_INSTQUEUE_REG_4__7_ & ~n27107;
  assign n4056 = ~n27101 | n27108;
  assign n27110 = n26128 & n27088;
  assign n27111 = n26130 & n27091;
  assign n27112 = n26136 & n27095;
  assign n27113 = ~n27110 & ~n27111;
  assign n27114 = ~n27112 & n27113;
  assign n27115 = n26133 & n27099;
  assign n27116 = n27114 & ~n27115;
  assign n27117 = P1_P3_INSTQUEUE_REG_4__6_ & ~n27107;
  assign n4061 = ~n27116 | n27117;
  assign n27119 = n26141 & n27088;
  assign n27120 = n26143 & n27091;
  assign n27121 = n26149 & n27095;
  assign n27122 = ~n27119 & ~n27120;
  assign n27123 = ~n27121 & n27122;
  assign n27124 = n26146 & n27099;
  assign n27125 = n27123 & ~n27124;
  assign n27126 = P1_P3_INSTQUEUE_REG_4__5_ & ~n27107;
  assign n4066 = ~n27125 | n27126;
  assign n27128 = n26154 & n27088;
  assign n27129 = n26156 & n27091;
  assign n27130 = n26162 & n27095;
  assign n27131 = ~n27128 & ~n27129;
  assign n27132 = ~n27130 & n27131;
  assign n27133 = n26159 & n27099;
  assign n27134 = n27132 & ~n27133;
  assign n27135 = P1_P3_INSTQUEUE_REG_4__4_ & ~n27107;
  assign n4071 = ~n27134 | n27135;
  assign n27137 = n26167 & n27088;
  assign n27138 = n26169 & n27091;
  assign n27139 = n26175 & n27095;
  assign n27140 = ~n27137 & ~n27138;
  assign n27141 = ~n27139 & n27140;
  assign n27142 = n26172 & n27099;
  assign n27143 = n27141 & ~n27142;
  assign n27144 = P1_P3_INSTQUEUE_REG_4__3_ & ~n27107;
  assign n4076 = ~n27143 | n27144;
  assign n27146 = n26180 & n27088;
  assign n27147 = n26182 & n27091;
  assign n27148 = n26188 & n27095;
  assign n27149 = ~n27146 & ~n27147;
  assign n27150 = ~n27148 & n27149;
  assign n27151 = n26185 & n27099;
  assign n27152 = n27150 & ~n27151;
  assign n27153 = P1_P3_INSTQUEUE_REG_4__2_ & ~n27107;
  assign n4081 = ~n27152 | n27153;
  assign n27155 = n26193 & n27088;
  assign n27156 = n26195 & n27091;
  assign n27157 = n26201 & n27095;
  assign n27158 = ~n27155 & ~n27156;
  assign n27159 = ~n27157 & n27158;
  assign n27160 = n26198 & n27099;
  assign n27161 = n27159 & ~n27160;
  assign n27162 = P1_P3_INSTQUEUE_REG_4__1_ & ~n27107;
  assign n4086 = ~n27161 | n27162;
  assign n27164 = n26206 & n27088;
  assign n27165 = n26208 & n27091;
  assign n27166 = n26214 & n27095;
  assign n27167 = ~n27164 & ~n27165;
  assign n27168 = ~n27166 & n27167;
  assign n27169 = n26211 & n27099;
  assign n27170 = n27168 & ~n27169;
  assign n27171 = P1_P3_INSTQUEUE_REG_4__0_ & ~n27107;
  assign n4091 = ~n27170 | n27171;
  assign n27173 = n26084 & n26093;
  assign n27174 = n26085 & n27173;
  assign n27175 = n26111 & n27174;
  assign n27176 = ~P1_P3_INSTQUEUEWR_ADDR_REG_3_ & ~P1_P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n27177 = n26050 & n27176;
  assign n27178 = n26114 & n27177;
  assign n27179 = n26061 & n26064;
  assign n27180 = n26069 & n27179;
  assign n27181 = ~n27177 & ~n27180;
  assign n27182 = ~n27093 & ~n27181;
  assign n27183 = n26123 & n27182;
  assign n27184 = ~n27175 & ~n27178;
  assign n27185 = ~n27183 & n27184;
  assign n27186 = n26088 & n26099;
  assign n27187 = n26081 & n27186;
  assign n27188 = n26117 & n27187;
  assign n27189 = n27185 & ~n27188;
  assign n27190 = P1_P3_STATE2_REG_3_ & ~n27177;
  assign n27191 = n26057 & ~n27190;
  assign n27192 = ~n27174 & ~n27187;
  assign n27193 = n26074 & ~n27192;
  assign n27194 = n27181 & ~n27193;
  assign n27195 = n27191 & ~n27194;
  assign n27196 = P1_P3_INSTQUEUE_REG_3__7_ & ~n27195;
  assign n4096 = ~n27189 | n27196;
  assign n27198 = n26128 & n27174;
  assign n27199 = n26130 & n27177;
  assign n27200 = n26136 & n27182;
  assign n27201 = ~n27198 & ~n27199;
  assign n27202 = ~n27200 & n27201;
  assign n27203 = n26133 & n27187;
  assign n27204 = n27202 & ~n27203;
  assign n27205 = P1_P3_INSTQUEUE_REG_3__6_ & ~n27195;
  assign n4101 = ~n27204 | n27205;
  assign n27207 = n26141 & n27174;
  assign n27208 = n26143 & n27177;
  assign n27209 = n26149 & n27182;
  assign n27210 = ~n27207 & ~n27208;
  assign n27211 = ~n27209 & n27210;
  assign n27212 = n26146 & n27187;
  assign n27213 = n27211 & ~n27212;
  assign n27214 = P1_P3_INSTQUEUE_REG_3__5_ & ~n27195;
  assign n4106 = ~n27213 | n27214;
  assign n27216 = n26154 & n27174;
  assign n27217 = n26156 & n27177;
  assign n27218 = n26162 & n27182;
  assign n27219 = ~n27216 & ~n27217;
  assign n27220 = ~n27218 & n27219;
  assign n27221 = n26159 & n27187;
  assign n27222 = n27220 & ~n27221;
  assign n27223 = P1_P3_INSTQUEUE_REG_3__4_ & ~n27195;
  assign n4111 = ~n27222 | n27223;
  assign n27225 = n26167 & n27174;
  assign n27226 = n26169 & n27177;
  assign n27227 = n26175 & n27182;
  assign n27228 = ~n27225 & ~n27226;
  assign n27229 = ~n27227 & n27228;
  assign n27230 = n26172 & n27187;
  assign n27231 = n27229 & ~n27230;
  assign n27232 = P1_P3_INSTQUEUE_REG_3__3_ & ~n27195;
  assign n4116 = ~n27231 | n27232;
  assign n27234 = n26180 & n27174;
  assign n27235 = n26182 & n27177;
  assign n27236 = n26188 & n27182;
  assign n27237 = ~n27234 & ~n27235;
  assign n27238 = ~n27236 & n27237;
  assign n27239 = n26185 & n27187;
  assign n27240 = n27238 & ~n27239;
  assign n27241 = P1_P3_INSTQUEUE_REG_3__2_ & ~n27195;
  assign n4121 = ~n27240 | n27241;
  assign n27243 = n26193 & n27174;
  assign n27244 = n26195 & n27177;
  assign n27245 = n26201 & n27182;
  assign n27246 = ~n27243 & ~n27244;
  assign n27247 = ~n27245 & n27246;
  assign n27248 = n26198 & n27187;
  assign n27249 = n27247 & ~n27248;
  assign n27250 = P1_P3_INSTQUEUE_REG_3__1_ & ~n27195;
  assign n4126 = ~n27249 | n27250;
  assign n27252 = n26206 & n27174;
  assign n27253 = n26208 & n27177;
  assign n27254 = n26214 & n27182;
  assign n27255 = ~n27252 & ~n27253;
  assign n27256 = ~n27254 & n27255;
  assign n27257 = n26211 & n27187;
  assign n27258 = n27256 & ~n27257;
  assign n27259 = P1_P3_INSTQUEUE_REG_3__0_ & ~n27195;
  assign n4131 = ~n27258 | n27259;
  assign n27261 = n26078 & n27173;
  assign n27262 = n26111 & n27261;
  assign n27263 = n26572 & n26914;
  assign n27264 = n26114 & n27263;
  assign n27265 = n26075 & n27179;
  assign n27266 = ~n27263 & ~n27265;
  assign n27267 = ~n27093 & ~n27266;
  assign n27268 = n26123 & n27267;
  assign n27269 = ~n27262 & ~n27264;
  assign n27270 = ~n27268 & n27269;
  assign n27271 = n26225 & n27186;
  assign n27272 = n26117 & n27271;
  assign n27273 = n27270 & ~n27272;
  assign n27274 = P1_P3_STATE2_REG_3_ & ~n27263;
  assign n27275 = n26057 & ~n27274;
  assign n27276 = ~n27261 & ~n27271;
  assign n27277 = n26074 & ~n27276;
  assign n27278 = n27266 & ~n27277;
  assign n27279 = n27275 & ~n27278;
  assign n27280 = P1_P3_INSTQUEUE_REG_2__7_ & ~n27279;
  assign n4136 = ~n27273 | n27280;
  assign n27282 = n26128 & n27261;
  assign n27283 = n26130 & n27263;
  assign n27284 = n26136 & n27267;
  assign n27285 = ~n27282 & ~n27283;
  assign n27286 = ~n27284 & n27285;
  assign n27287 = n26133 & n27271;
  assign n27288 = n27286 & ~n27287;
  assign n27289 = P1_P3_INSTQUEUE_REG_2__6_ & ~n27279;
  assign n4141 = ~n27288 | n27289;
  assign n27291 = n26141 & n27261;
  assign n27292 = n26143 & n27263;
  assign n27293 = n26149 & n27267;
  assign n27294 = ~n27291 & ~n27292;
  assign n27295 = ~n27293 & n27294;
  assign n27296 = n26146 & n27271;
  assign n27297 = n27295 & ~n27296;
  assign n27298 = P1_P3_INSTQUEUE_REG_2__5_ & ~n27279;
  assign n4146 = ~n27297 | n27298;
  assign n27300 = n26154 & n27261;
  assign n27301 = n26156 & n27263;
  assign n27302 = n26162 & n27267;
  assign n27303 = ~n27300 & ~n27301;
  assign n27304 = ~n27302 & n27303;
  assign n27305 = n26159 & n27271;
  assign n27306 = n27304 & ~n27305;
  assign n27307 = P1_P3_INSTQUEUE_REG_2__4_ & ~n27279;
  assign n4151 = ~n27306 | n27307;
  assign n27309 = n26167 & n27261;
  assign n27310 = n26169 & n27263;
  assign n27311 = n26175 & n27267;
  assign n27312 = ~n27309 & ~n27310;
  assign n27313 = ~n27311 & n27312;
  assign n27314 = n26172 & n27271;
  assign n27315 = n27313 & ~n27314;
  assign n27316 = P1_P3_INSTQUEUE_REG_2__3_ & ~n27279;
  assign n4156 = ~n27315 | n27316;
  assign n27318 = n26180 & n27261;
  assign n27319 = n26182 & n27263;
  assign n27320 = n26188 & n27267;
  assign n27321 = ~n27318 & ~n27319;
  assign n27322 = ~n27320 & n27321;
  assign n27323 = n26185 & n27271;
  assign n27324 = n27322 & ~n27323;
  assign n27325 = P1_P3_INSTQUEUE_REG_2__2_ & ~n27279;
  assign n4161 = ~n27324 | n27325;
  assign n27327 = n26193 & n27261;
  assign n27328 = n26195 & n27263;
  assign n27329 = n26201 & n27267;
  assign n27330 = ~n27327 & ~n27328;
  assign n27331 = ~n27329 & n27330;
  assign n27332 = n26198 & n27271;
  assign n27333 = n27331 & ~n27332;
  assign n27334 = P1_P3_INSTQUEUE_REG_2__1_ & ~n27279;
  assign n4166 = ~n27333 | n27334;
  assign n27336 = n26206 & n27261;
  assign n27337 = n26208 & n27263;
  assign n27338 = n26214 & n27267;
  assign n27339 = ~n27336 & ~n27337;
  assign n27340 = ~n27338 & n27339;
  assign n27341 = n26211 & n27271;
  assign n27342 = n27340 & ~n27341;
  assign n27343 = P1_P3_INSTQUEUE_REG_2__0_ & ~n27279;
  assign n4171 = ~n27342 | n27343;
  assign n27345 = n26079 & n27173;
  assign n27346 = n26111 & n27345;
  assign n27347 = n26066 & n27176;
  assign n27348 = n26114 & n27347;
  assign n27349 = n26076 & n27179;
  assign n27350 = ~n27347 & ~n27349;
  assign n27351 = ~n27093 & ~n27350;
  assign n27352 = n26123 & n27351;
  assign n27353 = ~n27346 & ~n27348;
  assign n27354 = ~n27352 & n27353;
  assign n27355 = n26313 & n27186;
  assign n27356 = n26117 & n27355;
  assign n27357 = n27354 & ~n27356;
  assign n27358 = P1_P3_STATE2_REG_3_ & ~n27347;
  assign n27359 = n26057 & ~n27358;
  assign n27360 = ~n27345 & ~n27355;
  assign n27361 = n26074 & ~n27360;
  assign n27362 = n27350 & ~n27361;
  assign n27363 = n27359 & ~n27362;
  assign n27364 = P1_P3_INSTQUEUE_REG_1__7_ & ~n27363;
  assign n4176 = ~n27357 | n27364;
  assign n27366 = n26128 & n27345;
  assign n27367 = n26130 & n27347;
  assign n27368 = n26136 & n27351;
  assign n27369 = ~n27366 & ~n27367;
  assign n27370 = ~n27368 & n27369;
  assign n27371 = n26133 & n27355;
  assign n27372 = n27370 & ~n27371;
  assign n27373 = P1_P3_INSTQUEUE_REG_1__6_ & ~n27363;
  assign n4181 = ~n27372 | n27373;
  assign n27375 = n26141 & n27345;
  assign n27376 = n26143 & n27347;
  assign n27377 = n26149 & n27351;
  assign n27378 = ~n27375 & ~n27376;
  assign n27379 = ~n27377 & n27378;
  assign n27380 = n26146 & n27355;
  assign n27381 = n27379 & ~n27380;
  assign n27382 = P1_P3_INSTQUEUE_REG_1__5_ & ~n27363;
  assign n4186 = ~n27381 | n27382;
  assign n27384 = n26154 & n27345;
  assign n27385 = n26156 & n27347;
  assign n27386 = n26162 & n27351;
  assign n27387 = ~n27384 & ~n27385;
  assign n27388 = ~n27386 & n27387;
  assign n27389 = n26159 & n27355;
  assign n27390 = n27388 & ~n27389;
  assign n27391 = P1_P3_INSTQUEUE_REG_1__4_ & ~n27363;
  assign n4191 = ~n27390 | n27391;
  assign n27393 = n26167 & n27345;
  assign n27394 = n26169 & n27347;
  assign n27395 = n26175 & n27351;
  assign n27396 = ~n27393 & ~n27394;
  assign n27397 = ~n27395 & n27396;
  assign n27398 = n26172 & n27355;
  assign n27399 = n27397 & ~n27398;
  assign n27400 = P1_P3_INSTQUEUE_REG_1__3_ & ~n27363;
  assign n4196 = ~n27399 | n27400;
  assign n27402 = n26180 & n27345;
  assign n27403 = n26182 & n27347;
  assign n27404 = n26188 & n27351;
  assign n27405 = ~n27402 & ~n27403;
  assign n27406 = ~n27404 & n27405;
  assign n27407 = n26185 & n27355;
  assign n27408 = n27406 & ~n27407;
  assign n27409 = P1_P3_INSTQUEUE_REG_1__2_ & ~n27363;
  assign n4201 = ~n27408 | n27409;
  assign n27411 = n26193 & n27345;
  assign n27412 = n26195 & n27347;
  assign n27413 = n26201 & n27351;
  assign n27414 = ~n27411 & ~n27412;
  assign n27415 = ~n27413 & n27414;
  assign n27416 = n26198 & n27355;
  assign n27417 = n27415 & ~n27416;
  assign n27418 = P1_P3_INSTQUEUE_REG_1__1_ & ~n27363;
  assign n4206 = ~n27417 | n27418;
  assign n27420 = n26206 & n27345;
  assign n27421 = n26208 & n27347;
  assign n27422 = n26214 & n27351;
  assign n27423 = ~n27420 & ~n27421;
  assign n27424 = ~n27422 & n27423;
  assign n27425 = n26211 & n27355;
  assign n27426 = n27424 & ~n27425;
  assign n27427 = P1_P3_INSTQUEUE_REG_1__0_ & ~n27363;
  assign n4211 = ~n27426 | n27427;
  assign n27429 = n26401 & n27173;
  assign n27430 = n26111 & n27429;
  assign n27431 = n26572 & n27090;
  assign n27432 = n26114 & n27431;
  assign n27433 = n26068 & n27179;
  assign n27434 = ~n27093 & n27433;
  assign n27435 = n26123 & n27434;
  assign n27436 = ~n27430 & ~n27432;
  assign n27437 = ~n27435 & n27436;
  assign n27438 = n26399 & n27186;
  assign n27439 = n26117 & n27438;
  assign n27440 = n27437 & ~n27439;
  assign n27441 = P1_P3_STATE2_REG_3_ & ~n27431;
  assign n27442 = n26057 & ~n27441;
  assign n27443 = ~n27429 & ~n27438;
  assign n27444 = n26074 & ~n27443;
  assign n27445 = ~n27433 & ~n27444;
  assign n27446 = n27442 & ~n27445;
  assign n27447 = P1_P3_INSTQUEUE_REG_0__7_ & ~n27446;
  assign n4216 = ~n27440 | n27447;
  assign n27449 = n26128 & n27429;
  assign n27450 = n26130 & n27431;
  assign n27451 = n26136 & n27434;
  assign n27452 = ~n27449 & ~n27450;
  assign n27453 = ~n27451 & n27452;
  assign n27454 = n26133 & n27438;
  assign n27455 = n27453 & ~n27454;
  assign n27456 = P1_P3_INSTQUEUE_REG_0__6_ & ~n27446;
  assign n4221 = ~n27455 | n27456;
  assign n27458 = n26141 & n27429;
  assign n27459 = n26143 & n27431;
  assign n27460 = n26149 & n27434;
  assign n27461 = ~n27458 & ~n27459;
  assign n27462 = ~n27460 & n27461;
  assign n27463 = n26146 & n27438;
  assign n27464 = n27462 & ~n27463;
  assign n27465 = P1_P3_INSTQUEUE_REG_0__5_ & ~n27446;
  assign n4226 = ~n27464 | n27465;
  assign n27467 = n26154 & n27429;
  assign n27468 = n26156 & n27431;
  assign n27469 = n26162 & n27434;
  assign n27470 = ~n27467 & ~n27468;
  assign n27471 = ~n27469 & n27470;
  assign n27472 = n26159 & n27438;
  assign n27473 = n27471 & ~n27472;
  assign n27474 = P1_P3_INSTQUEUE_REG_0__4_ & ~n27446;
  assign n4231 = ~n27473 | n27474;
  assign n27476 = n26167 & n27429;
  assign n27477 = n26169 & n27431;
  assign n27478 = n26175 & n27434;
  assign n27479 = ~n27476 & ~n27477;
  assign n27480 = ~n27478 & n27479;
  assign n27481 = n26172 & n27438;
  assign n27482 = n27480 & ~n27481;
  assign n27483 = P1_P3_INSTQUEUE_REG_0__3_ & ~n27446;
  assign n4236 = ~n27482 | n27483;
  assign n27485 = n26180 & n27429;
  assign n27486 = n26182 & n27431;
  assign n27487 = n26188 & n27434;
  assign n27488 = ~n27485 & ~n27486;
  assign n27489 = ~n27487 & n27488;
  assign n27490 = n26185 & n27438;
  assign n27491 = n27489 & ~n27490;
  assign n27492 = P1_P3_INSTQUEUE_REG_0__2_ & ~n27446;
  assign n4241 = ~n27491 | n27492;
  assign n27494 = n26193 & n27429;
  assign n27495 = n26195 & n27431;
  assign n27496 = n26201 & n27434;
  assign n27497 = ~n27494 & ~n27495;
  assign n27498 = ~n27496 & n27497;
  assign n27499 = n26198 & n27438;
  assign n27500 = n27498 & ~n27499;
  assign n27501 = P1_P3_INSTQUEUE_REG_0__1_ & ~n27446;
  assign n4246 = ~n27500 | n27501;
  assign n27503 = n26206 & n27429;
  assign n27504 = n26208 & n27431;
  assign n27505 = n26214 & n27434;
  assign n27506 = ~n27503 & ~n27504;
  assign n27507 = ~n27505 & n27506;
  assign n27508 = n26211 & n27438;
  assign n27509 = n27507 & ~n27508;
  assign n27510 = P1_P3_INSTQUEUE_REG_0__0_ & ~n27446;
  assign n4251 = ~n27509 | n27510;
  assign n27512 = P1_P3_STATE2_REG_3_ & ~P1_P3_STATE2_REG_0_;
  assign n27513 = P1_P3_STATE2_REG_0_ & P1_P3_FLUSH_REG;
  assign n27514 = n25352 & n27513;
  assign n27515 = ~n27512 & ~n27514;
  assign n27516 = ~n25884 & n25994;
  assign n27517 = n27515 & ~n27516;
  assign n27518 = P1_P3_INSTQUEUERD_ADDR_REG_4_ & n27517;
  assign n27519 = ~n25927 & n26000;
  assign n27520 = n25719 & n27519;
  assign n27521 = ~n27517 & n27520;
  assign n4256 = n27518 | n27521;
  assign n27523 = ~n25918 & n26000;
  assign n27524 = ~n25391 & ~n25891;
  assign n27525 = n26009 & ~n27524;
  assign n27526 = ~n27523 & ~n27525;
  assign n27527 = ~n27517 & ~n27526;
  assign n27528 = P1_P3_INSTQUEUERD_ADDR_REG_3_ & n27517;
  assign n4261 = n27527 | n27528;
  assign n27530 = ~n25842 & n26009;
  assign n27531 = P1_P3_STATE2_REG_1_ & ~n26016;
  assign n27532 = ~n26025 & n27531;
  assign n27533 = ~n27530 & ~n27532;
  assign n27534 = ~n25858 & n26000;
  assign n27535 = n27533 & ~n27534;
  assign n27536 = ~n27517 & ~n27535;
  assign n27537 = P1_P3_INSTQUEUERD_ADDR_REG_2_ & n27517;
  assign n4266 = n27536 | n27537;
  assign n27539 = n25954 & n26009;
  assign n27540 = n26025 & n27531;
  assign n27541 = ~n27539 & ~n27540;
  assign n27542 = ~n25959 & n26000;
  assign n27543 = n27541 & ~n27542;
  assign n27544 = ~n27517 & ~n27543;
  assign n27545 = P1_P3_INSTQUEUERD_ADDR_REG_1_ & n27517;
  assign n4271 = n27544 | n27545;
  assign n27547 = P1_P3_STATE2_REG_1_ & n26016;
  assign n27548 = ~P1_P3_INSTQUEUERD_ADDR_REG_0_ & n26009;
  assign n27549 = ~n27547 & ~n27548;
  assign n27550 = ~n25945 & n26000;
  assign n27551 = n27549 & ~n27550;
  assign n27552 = ~n27517 & ~n27551;
  assign n27553 = P1_P3_INSTQUEUERD_ADDR_REG_0_ & n27517;
  assign n4276 = n27552 | n27553;
  assign n27555 = P1_P3_STATE2_REG_0_ & n25352;
  assign n27556 = ~n26039 & n27555;
  assign n27557 = ~n26057 & ~n27514;
  assign n27558 = ~n27556 & n27557;
  assign n4281 = P1_P3_INSTQUEUEWR_ADDR_REG_4_ & n27558;
  assign n27560 = P1_P3_STATE2_REG_3_ & ~n26051;
  assign n27561 = ~n27558 & ~n27560;
  assign n27562 = P1_P3_INSTQUEUEWR_ADDR_REG_3_ & ~n27561;
  assign n27563 = ~n26000 & ~n26073;
  assign n27564 = ~n26093 & ~n27563;
  assign n27565 = P1_P3_STATE2_REG_3_ & n26062;
  assign n27566 = ~n27564 & ~n27565;
  assign n27567 = n26081 & ~n26088;
  assign n27568 = ~n26099 & ~n27567;
  assign n27569 = ~n26834 & ~n27568;
  assign n27570 = n26109 & ~n27569;
  assign n27571 = n27566 & ~n27570;
  assign n27572 = ~n27558 & ~n27571;
  assign n4286 = n27562 | n27572;
  assign n27574 = ~n26084 & ~n27563;
  assign n27575 = P1_P3_STATE2_REG_3_ & ~P1_P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n27576 = n26050 & n27575;
  assign n27577 = ~n27574 & ~n27576;
  assign n27578 = ~n26081 & ~n26088;
  assign n27579 = n26081 & n26088;
  assign n27580 = ~n27578 & ~n27579;
  assign n27581 = n26109 & ~n27580;
  assign n27582 = n27577 & ~n27581;
  assign n27583 = ~n27558 & ~n27582;
  assign n27584 = P1_P3_STATE2_REG_3_ & ~n26050;
  assign n27585 = ~n27558 & ~n27584;
  assign n27586 = P1_P3_INSTQUEUEWR_ADDR_REG_2_ & ~n27585;
  assign n4291 = n27583 | n27586;
  assign n27588 = ~n26077 & ~n27563;
  assign n27589 = P1_P3_STATE2_REG_3_ & ~P1_P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n27590 = ~n26080 & n26109;
  assign n27591 = ~n27589 & ~n27590;
  assign n27592 = P1_P3_INSTQUEUEWR_ADDR_REG_0_ & ~n27591;
  assign n27593 = n26109 & n26313;
  assign n27594 = ~n27588 & ~n27592;
  assign n27595 = ~n27593 & n27594;
  assign n27596 = ~n27558 & ~n27595;
  assign n27597 = P1_P3_STATE2_REG_3_ & ~P1_P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n27598 = ~n27558 & ~n27597;
  assign n27599 = P1_P3_INSTQUEUEWR_ADDR_REG_1_ & ~n27598;
  assign n4296 = n27596 | n27599;
  assign n27601 = ~n26000 & ~n26072;
  assign n27602 = ~n27558 & n27601;
  assign n27603 = P1_P3_INSTQUEUEWR_ADDR_REG_0_ & ~n27602;
  assign n27604 = ~n26040 & ~n27597;
  assign n27605 = ~n27558 & ~n27604;
  assign n4301 = n27603 | n27605;
  assign n27607 = ~P1_P3_STATE2_REG_1_ & n26072;
  assign n27608 = ~P1_P3_STATE2_REG_0_ & n27607;
  assign n27609 = n25648 & n25692;
  assign n27610 = ~n25480 & ~n25639;
  assign n27611 = n25737 & n27610;
  assign n27612 = n25646 & n25692;
  assign n27613 = ~n25876 & ~n27611;
  assign n27614 = ~n27612 & n27613;
  assign n27615 = n25697 & n25745;
  assign n27616 = n25449 & n25644;
  assign n27617 = n25692 & n27616;
  assign n27618 = ~n27615 & ~n27617;
  assign n27619 = n25608 & ~n27618;
  assign n27620 = ~n25448 & n25751;
  assign n27621 = ~n25267 & n25417;
  assign n27622 = n25692 & n27621;
  assign n27623 = ~n27620 & ~n27622;
  assign n27624 = ~n25608 & ~n27623;
  assign n27625 = n25639 & n25737;
  assign n27626 = ~n27619 & ~n27624;
  assign n27627 = ~n27625 & n27626;
  assign n27628 = n25573 & ~n27627;
  assign n27629 = n25868 & ~n27609;
  assign n27630 = n27614 & n27629;
  assign n27631 = ~n27628 & n27630;
  assign n27632 = n25994 & ~n27631;
  assign n27633 = ~n27608 & ~n27632;
  assign n27634 = P1_P3_STATE2_REG_2_ & ~n27633;
  assign n27635 = ~P1_P3_INSTADDRPOINTER_REG_0_ & n25938;
  assign n27636 = ~P1_P3_INSTADDRPOINTER_REG_0_ & n25781;
  assign n27637 = ~n27635 & ~n27636;
  assign n27638 = ~P1_P3_INSTADDRPOINTER_REG_0_ & ~n25828;
  assign n27639 = P1_P3_INSTADDRPOINTER_REG_0_ & n25899;
  assign n27640 = P1_P3_INSTADDRPOINTER_REG_0_ & n25900;
  assign n27641 = n25640 & n25771;
  assign n27642 = n25777 & n27641;
  assign n27643 = ~P1_P3_INSTADDRPOINTER_REG_0_ & n27642;
  assign n27644 = n25717 & n25771;
  assign n27645 = n25777 & n27644;
  assign n27646 = ~P1_P3_INSTADDRPOINTER_REG_0_ & n27645;
  assign n27647 = ~n27643 & ~n27646;
  assign n27648 = P1_P3_INSTADDRPOINTER_REG_0_ & n25715;
  assign n27649 = n27647 & ~n27648;
  assign n27650 = n25842 & n27524;
  assign n27651 = P1_P3_INSTQUEUERD_ADDR_REG_0_ & ~n25954;
  assign n27652 = n27650 & n27651;
  assign n27653 = P1_P3_INSTQUEUE_REG_0__0_ & n27652;
  assign n27654 = ~P1_P3_INSTQUEUERD_ADDR_REG_0_ & ~n25954;
  assign n27655 = n27650 & n27654;
  assign n27656 = P1_P3_INSTQUEUE_REG_1__0_ & n27655;
  assign n27657 = P1_P3_INSTQUEUERD_ADDR_REG_0_ & n25954;
  assign n27658 = n27650 & n27657;
  assign n27659 = P1_P3_INSTQUEUE_REG_2__0_ & n27658;
  assign n27660 = ~P1_P3_INSTQUEUERD_ADDR_REG_0_ & n25954;
  assign n27661 = n27650 & n27660;
  assign n27662 = P1_P3_INSTQUEUE_REG_3__0_ & n27661;
  assign n27663 = ~n27653 & ~n27656;
  assign n27664 = ~n27659 & n27663;
  assign n27665 = ~n27662 & n27664;
  assign n27666 = ~n25842 & n27524;
  assign n27667 = n27651 & n27666;
  assign n27668 = P1_P3_INSTQUEUE_REG_4__0_ & n27667;
  assign n27669 = n27654 & n27666;
  assign n27670 = P1_P3_INSTQUEUE_REG_5__0_ & n27669;
  assign n27671 = n27657 & n27666;
  assign n27672 = P1_P3_INSTQUEUE_REG_6__0_ & n27671;
  assign n27673 = n27660 & n27666;
  assign n27674 = P1_P3_INSTQUEUE_REG_7__0_ & n27673;
  assign n27675 = ~n27668 & ~n27670;
  assign n27676 = ~n27672 & n27675;
  assign n27677 = ~n27674 & n27676;
  assign n27678 = n25842 & ~n27524;
  assign n27679 = n27651 & n27678;
  assign n27680 = P1_P3_INSTQUEUE_REG_8__0_ & n27679;
  assign n27681 = n27654 & n27678;
  assign n27682 = P1_P3_INSTQUEUE_REG_9__0_ & n27681;
  assign n27683 = n27657 & n27678;
  assign n27684 = P1_P3_INSTQUEUE_REG_10__0_ & n27683;
  assign n27685 = n27660 & n27678;
  assign n27686 = P1_P3_INSTQUEUE_REG_11__0_ & n27685;
  assign n27687 = ~n27680 & ~n27682;
  assign n27688 = ~n27684 & n27687;
  assign n27689 = ~n27686 & n27688;
  assign n27690 = ~n25842 & ~n27524;
  assign n27691 = n27651 & n27690;
  assign n27692 = P1_P3_INSTQUEUE_REG_12__0_ & n27691;
  assign n27693 = n27654 & n27690;
  assign n27694 = P1_P3_INSTQUEUE_REG_13__0_ & n27693;
  assign n27695 = n27657 & n27690;
  assign n27696 = P1_P3_INSTQUEUE_REG_14__0_ & n27695;
  assign n27697 = n27660 & n27690;
  assign n27698 = P1_P3_INSTQUEUE_REG_15__0_ & n27697;
  assign n27699 = ~n27692 & ~n27694;
  assign n27700 = ~n27696 & n27699;
  assign n27701 = ~n27698 & n27700;
  assign n27702 = n27665 & n27677;
  assign n27703 = n27689 & n27702;
  assign n27704 = n27701 & n27703;
  assign n27705 = ~P1_P3_INSTADDRPOINTER_REG_0_ & ~n27704;
  assign n27706 = P1_P3_INSTADDRPOINTER_REG_0_ & n27704;
  assign n27707 = ~n27705 & ~n27706;
  assign n27708 = P1_P3_INSTQUEUE_REG_0__7_ & n27652;
  assign n27709 = P1_P3_INSTQUEUE_REG_1__7_ & n27655;
  assign n27710 = P1_P3_INSTQUEUE_REG_2__7_ & n27658;
  assign n27711 = P1_P3_INSTQUEUE_REG_3__7_ & n27661;
  assign n27712 = ~n27708 & ~n27709;
  assign n27713 = ~n27710 & n27712;
  assign n27714 = ~n27711 & n27713;
  assign n27715 = P1_P3_INSTQUEUE_REG_4__7_ & n27667;
  assign n27716 = P1_P3_INSTQUEUE_REG_5__7_ & n27669;
  assign n27717 = P1_P3_INSTQUEUE_REG_6__7_ & n27671;
  assign n27718 = P1_P3_INSTQUEUE_REG_7__7_ & n27673;
  assign n27719 = ~n27715 & ~n27716;
  assign n27720 = ~n27717 & n27719;
  assign n27721 = ~n27718 & n27720;
  assign n27722 = P1_P3_INSTQUEUE_REG_8__7_ & n27679;
  assign n27723 = P1_P3_INSTQUEUE_REG_9__7_ & n27681;
  assign n27724 = P1_P3_INSTQUEUE_REG_10__7_ & n27683;
  assign n27725 = P1_P3_INSTQUEUE_REG_11__7_ & n27685;
  assign n27726 = ~n27722 & ~n27723;
  assign n27727 = ~n27724 & n27726;
  assign n27728 = ~n27725 & n27727;
  assign n27729 = P1_P3_INSTQUEUE_REG_12__7_ & n27691;
  assign n27730 = P1_P3_INSTQUEUE_REG_13__7_ & n27693;
  assign n27731 = P1_P3_INSTQUEUE_REG_14__7_ & n27695;
  assign n27732 = P1_P3_INSTQUEUE_REG_15__7_ & n27697;
  assign n27733 = ~n27729 & ~n27730;
  assign n27734 = ~n27731 & n27733;
  assign n27735 = ~n27732 & n27734;
  assign n27736 = n27714 & n27721;
  assign n27737 = n27728 & n27736;
  assign n27738 = n27735 & n27737;
  assign n27739 = n25747 & ~n27738;
  assign n27740 = ~n27707 & n27739;
  assign n27741 = n25747 & n27738;
  assign n27742 = ~n27707 & n27741;
  assign n27743 = ~n27639 & ~n27640;
  assign n27744 = n27649 & n27743;
  assign n27745 = ~n27740 & n27744;
  assign n27746 = ~n27742 & n27745;
  assign n27747 = n25713 & n25741;
  assign n27748 = ~P1_P3_INSTADDRPOINTER_REG_0_ & n27747;
  assign n27749 = ~P1_P3_INSTADDRPOINTER_REG_0_ & n25785;
  assign n27750 = n25542 & n25728;
  assign n27751 = n25774 & n27750;
  assign n27752 = ~P1_P3_INSTADDRPOINTER_REG_0_ & n27751;
  assign n27753 = ~P1_P3_INSTADDRPOINTER_REG_0_ & n27704;
  assign n27754 = P1_P3_INSTADDRPOINTER_REG_0_ & ~n27704;
  assign n27755 = ~n27753 & ~n27754;
  assign n27756 = n25742 & ~n27755;
  assign n27757 = n25417 & n25771;
  assign n27758 = n25774 & n27757;
  assign n27759 = ~P1_P3_INSTADDRPOINTER_REG_0_ & n27758;
  assign n27760 = ~n27748 & ~n27749;
  assign n27761 = ~n27752 & n27760;
  assign n27762 = ~n27756 & n27761;
  assign n27763 = ~n27759 & n27762;
  assign n27764 = P1_P3_INSTADDRPOINTER_REG_0_ & n25641;
  assign n27765 = P1_P3_INSTADDRPOINTER_REG_0_ & n25719;
  assign n27766 = P1_P3_INSTADDRPOINTER_REG_0_ & n25723;
  assign n27767 = ~P1_P3_INSTADDRPOINTER_REG_0_ & n25739;
  assign n27768 = ~P1_P3_INSTADDRPOINTER_REG_0_ & n25731;
  assign n27769 = ~n27764 & ~n27765;
  assign n27770 = ~n27766 & n27769;
  assign n27771 = ~n27767 & n27770;
  assign n27772 = ~n27768 & n27771;
  assign n27773 = n27763 & n27772;
  assign n27774 = n27637 & ~n27638;
  assign n27775 = n27746 & n27774;
  assign n27776 = n27773 & n27775;
  assign n27777 = n27634 & ~n27776;
  assign n27778 = ~P1_P3_STATE2_REG_2_ & ~n27633;
  assign n27779 = P1_P3_REIP_REG_0_ & n27778;
  assign n27780 = P1_P3_INSTADDRPOINTER_REG_0_ & n27633;
  assign n27781 = ~n27777 & ~n27779;
  assign n4306 = n27780 | ~n27781;
  assign n27783 = P1_P3_INSTADDRPOINTER_REG_1_ & n27633;
  assign n27784 = P1_P3_REIP_REG_1_ & n27778;
  assign n27785 = ~n25828 & ~n26022;
  assign n27786 = n25938 & ~n26022;
  assign n27787 = n25781 & ~n26022;
  assign n27788 = ~n27786 & ~n27787;
  assign n27789 = ~P1_P3_INSTADDRPOINTER_REG_1_ & n27754;
  assign n27790 = P1_P3_INSTADDRPOINTER_REG_1_ & ~n27754;
  assign n27791 = ~n27789 & ~n27790;
  assign n27792 = P1_P3_INSTQUEUE_REG_0__1_ & n27652;
  assign n27793 = P1_P3_INSTQUEUE_REG_1__1_ & n27655;
  assign n27794 = P1_P3_INSTQUEUE_REG_2__1_ & n27658;
  assign n27795 = P1_P3_INSTQUEUE_REG_3__1_ & n27661;
  assign n27796 = ~n27792 & ~n27793;
  assign n27797 = ~n27794 & n27796;
  assign n27798 = ~n27795 & n27797;
  assign n27799 = P1_P3_INSTQUEUE_REG_4__1_ & n27667;
  assign n27800 = P1_P3_INSTQUEUE_REG_5__1_ & n27669;
  assign n27801 = P1_P3_INSTQUEUE_REG_6__1_ & n27671;
  assign n27802 = P1_P3_INSTQUEUE_REG_7__1_ & n27673;
  assign n27803 = ~n27799 & ~n27800;
  assign n27804 = ~n27801 & n27803;
  assign n27805 = ~n27802 & n27804;
  assign n27806 = P1_P3_INSTQUEUE_REG_8__1_ & n27679;
  assign n27807 = P1_P3_INSTQUEUE_REG_9__1_ & n27681;
  assign n27808 = P1_P3_INSTQUEUE_REG_10__1_ & n27683;
  assign n27809 = P1_P3_INSTQUEUE_REG_11__1_ & n27685;
  assign n27810 = ~n27806 & ~n27807;
  assign n27811 = ~n27808 & n27810;
  assign n27812 = ~n27809 & n27811;
  assign n27813 = P1_P3_INSTQUEUE_REG_12__1_ & n27691;
  assign n27814 = P1_P3_INSTQUEUE_REG_13__1_ & n27693;
  assign n27815 = P1_P3_INSTQUEUE_REG_14__1_ & n27695;
  assign n27816 = P1_P3_INSTQUEUE_REG_15__1_ & n27697;
  assign n27817 = ~n27813 & ~n27814;
  assign n27818 = ~n27815 & n27817;
  assign n27819 = ~n27816 & n27818;
  assign n27820 = n27798 & n27805;
  assign n27821 = n27812 & n27820;
  assign n27822 = n27819 & n27821;
  assign n27823 = ~n27791 & ~n27822;
  assign n27824 = ~P1_P3_INSTADDRPOINTER_REG_1_ & ~n27754;
  assign n27825 = n27822 & n27824;
  assign n27826 = n27754 & n27822;
  assign n27827 = P1_P3_INSTADDRPOINTER_REG_1_ & n27826;
  assign n27828 = ~n27823 & ~n27825;
  assign n27829 = ~n27827 & n27828;
  assign n27830 = n27741 & ~n27829;
  assign n27831 = ~n26022 & n27758;
  assign n27832 = ~n26022 & n27751;
  assign n27833 = ~n26022 & n27747;
  assign n27834 = n25785 & ~n26022;
  assign n27835 = ~n27831 & ~n27832;
  assign n27836 = ~n27833 & n27835;
  assign n27837 = ~n27834 & n27836;
  assign n27838 = ~P1_P3_INSTADDRPOINTER_REG_1_ & n25641;
  assign n27839 = ~P1_P3_INSTADDRPOINTER_REG_1_ & n25719;
  assign n27840 = ~P1_P3_INSTADDRPOINTER_REG_1_ & n25723;
  assign n27841 = n25739 & ~n26022;
  assign n27842 = n25731 & ~n26022;
  assign n27843 = ~n27838 & ~n27839;
  assign n27844 = ~n27840 & n27843;
  assign n27845 = ~n27841 & n27844;
  assign n27846 = ~n27842 & n27845;
  assign n27847 = ~P1_P3_INSTADDRPOINTER_REG_1_ & n27706;
  assign n27848 = P1_P3_INSTADDRPOINTER_REG_1_ & ~n27706;
  assign n27849 = ~n27847 & ~n27848;
  assign n27850 = ~n27704 & n27822;
  assign n27851 = n27704 & ~n27822;
  assign n27852 = ~n27850 & ~n27851;
  assign n27853 = ~n27849 & n27852;
  assign n27854 = ~P1_P3_INSTADDRPOINTER_REG_1_ & ~n27706;
  assign n27855 = ~n27852 & n27854;
  assign n27856 = n27706 & ~n27852;
  assign n27857 = P1_P3_INSTADDRPOINTER_REG_1_ & n27856;
  assign n27858 = ~n27853 & ~n27855;
  assign n27859 = ~n27857 & n27858;
  assign n27860 = n25742 & ~n27859;
  assign n27861 = n27837 & n27846;
  assign n27862 = ~n27860 & n27861;
  assign n27863 = ~P1_P3_INSTADDRPOINTER_REG_1_ & n25899;
  assign n27864 = ~P1_P3_INSTADDRPOINTER_REG_1_ & n25900;
  assign n27865 = ~n26022 & n27642;
  assign n27866 = ~n26022 & n27645;
  assign n27867 = ~n27865 & ~n27866;
  assign n27868 = ~P1_P3_INSTADDRPOINTER_REG_1_ & n25715;
  assign n27869 = n27867 & ~n27868;
  assign n27870 = n27739 & ~n27829;
  assign n27871 = ~n27863 & ~n27864;
  assign n27872 = n27869 & n27871;
  assign n27873 = ~n27870 & n27872;
  assign n27874 = ~n27785 & n27788;
  assign n27875 = ~n27830 & n27874;
  assign n27876 = n27862 & n27875;
  assign n27877 = n27873 & n27876;
  assign n27878 = n27634 & ~n27877;
  assign n27879 = ~n27783 & ~n27784;
  assign n4311 = n27878 | ~n27879;
  assign n27881 = P1_P3_INSTADDRPOINTER_REG_2_ & n27633;
  assign n27882 = P1_P3_REIP_REG_2_ & n27778;
  assign n27883 = P1_P3_INSTADDRPOINTER_REG_0_ & P1_P3_INSTADDRPOINTER_REG_1_;
  assign n27884 = ~P1_P3_INSTADDRPOINTER_REG_2_ & n27883;
  assign n27885 = P1_P3_INSTADDRPOINTER_REG_2_ & ~n27883;
  assign n27886 = ~n27884 & ~n27885;
  assign n27887 = ~n25828 & ~n27886;
  assign n27888 = P1_P3_INSTADDRPOINTER_REG_1_ & ~P1_P3_INSTADDRPOINTER_REG_2_;
  assign n27889 = ~P1_P3_INSTADDRPOINTER_REG_1_ & P1_P3_INSTADDRPOINTER_REG_2_;
  assign n27890 = ~n27888 & ~n27889;
  assign n27891 = n25899 & ~n27890;
  assign n27892 = n25900 & ~n27890;
  assign n27893 = n27642 & ~n27886;
  assign n27894 = n27645 & ~n27886;
  assign n27895 = ~n27893 & ~n27894;
  assign n27896 = n25715 & ~n27890;
  assign n27897 = n27895 & ~n27896;
  assign n27898 = ~n27891 & ~n27892;
  assign n27899 = n27897 & n27898;
  assign n27900 = ~n27754 & ~n27822;
  assign n27901 = P1_P3_INSTADDRPOINTER_REG_1_ & ~n27900;
  assign n27902 = ~n27826 & ~n27901;
  assign n27903 = P1_P3_INSTQUEUE_REG_0__2_ & n27652;
  assign n27904 = P1_P3_INSTQUEUE_REG_1__2_ & n27655;
  assign n27905 = P1_P3_INSTQUEUE_REG_2__2_ & n27658;
  assign n27906 = P1_P3_INSTQUEUE_REG_3__2_ & n27661;
  assign n27907 = ~n27903 & ~n27904;
  assign n27908 = ~n27905 & n27907;
  assign n27909 = ~n27906 & n27908;
  assign n27910 = P1_P3_INSTQUEUE_REG_4__2_ & n27667;
  assign n27911 = P1_P3_INSTQUEUE_REG_5__2_ & n27669;
  assign n27912 = P1_P3_INSTQUEUE_REG_6__2_ & n27671;
  assign n27913 = P1_P3_INSTQUEUE_REG_7__2_ & n27673;
  assign n27914 = ~n27910 & ~n27911;
  assign n27915 = ~n27912 & n27914;
  assign n27916 = ~n27913 & n27915;
  assign n27917 = P1_P3_INSTQUEUE_REG_8__2_ & n27679;
  assign n27918 = P1_P3_INSTQUEUE_REG_9__2_ & n27681;
  assign n27919 = P1_P3_INSTQUEUE_REG_10__2_ & n27683;
  assign n27920 = P1_P3_INSTQUEUE_REG_11__2_ & n27685;
  assign n27921 = ~n27917 & ~n27918;
  assign n27922 = ~n27919 & n27921;
  assign n27923 = ~n27920 & n27922;
  assign n27924 = P1_P3_INSTQUEUE_REG_12__2_ & n27691;
  assign n27925 = P1_P3_INSTQUEUE_REG_13__2_ & n27693;
  assign n27926 = P1_P3_INSTQUEUE_REG_14__2_ & n27695;
  assign n27927 = P1_P3_INSTQUEUE_REG_15__2_ & n27697;
  assign n27928 = ~n27924 & ~n27925;
  assign n27929 = ~n27926 & n27928;
  assign n27930 = ~n27927 & n27929;
  assign n27931 = n27909 & n27916;
  assign n27932 = n27923 & n27931;
  assign n27933 = n27930 & n27932;
  assign n27934 = ~n27822 & n27933;
  assign n27935 = n27822 & ~n27933;
  assign n27936 = ~n27934 & ~n27935;
  assign n27937 = ~P1_P3_INSTADDRPOINTER_REG_2_ & ~n27936;
  assign n27938 = P1_P3_INSTADDRPOINTER_REG_2_ & n27936;
  assign n27939 = ~n27937 & ~n27938;
  assign n27940 = n27902 & ~n27939;
  assign n27941 = ~n27902 & n27939;
  assign n27942 = ~n27940 & ~n27941;
  assign n27943 = n27741 & ~n27942;
  assign n27944 = n25938 & ~n27886;
  assign n27945 = n25781 & ~n27886;
  assign n27946 = ~n27944 & ~n27945;
  assign n27947 = P1_P3_INSTADDRPOINTER_REG_1_ & n27754;
  assign n27948 = P1_P3_INSTADDRPOINTER_REG_1_ & n27822;
  assign n27949 = ~n27826 & ~n27947;
  assign n27950 = ~n27948 & n27949;
  assign n27951 = ~n27939 & n27950;
  assign n27952 = ~P1_P3_INSTADDRPOINTER_REG_2_ & n27936;
  assign n27953 = P1_P3_INSTADDRPOINTER_REG_2_ & ~n27936;
  assign n27954 = ~n27952 & ~n27953;
  assign n27955 = ~n27950 & ~n27954;
  assign n27956 = ~n27951 & ~n27955;
  assign n27957 = n27739 & ~n27956;
  assign n27958 = n27946 & ~n27957;
  assign n27959 = n27758 & ~n27886;
  assign n27960 = n27751 & ~n27886;
  assign n27961 = n27747 & ~n27886;
  assign n27962 = n25785 & ~n27886;
  assign n27963 = ~n27959 & ~n27960;
  assign n27964 = ~n27961 & n27963;
  assign n27965 = ~n27962 & n27964;
  assign n27966 = n25641 & ~n27890;
  assign n27967 = n25719 & ~n27890;
  assign n27968 = n25723 & ~n27890;
  assign n27969 = ~P1_P3_INSTADDRPOINTER_REG_2_ & ~n27883;
  assign n27970 = P1_P3_INSTADDRPOINTER_REG_2_ & n27883;
  assign n27971 = ~n27969 & ~n27970;
  assign n27972 = n25739 & ~n27971;
  assign n27973 = n25731 & ~n27971;
  assign n27974 = ~n27966 & ~n27967;
  assign n27975 = ~n27968 & n27974;
  assign n27976 = ~n27972 & n27975;
  assign n27977 = ~n27973 & n27976;
  assign n27978 = ~n27704 & ~n27822;
  assign n27979 = n27933 & ~n27978;
  assign n27980 = ~n27933 & n27978;
  assign n27981 = ~n27979 & ~n27980;
  assign n27982 = ~P1_P3_INSTADDRPOINTER_REG_2_ & ~n27981;
  assign n27983 = P1_P3_INSTADDRPOINTER_REG_2_ & n27981;
  assign n27984 = ~n27982 & ~n27983;
  assign n27985 = ~n27706 & n27852;
  assign n27986 = P1_P3_INSTADDRPOINTER_REG_1_ & ~n27985;
  assign n27987 = ~n27856 & ~n27986;
  assign n27988 = ~n27984 & n27987;
  assign n27989 = ~P1_P3_INSTADDRPOINTER_REG_2_ & n27981;
  assign n27990 = P1_P3_INSTADDRPOINTER_REG_2_ & ~n27981;
  assign n27991 = ~n27989 & ~n27990;
  assign n27992 = ~n27987 & ~n27991;
  assign n27993 = ~n27988 & ~n27992;
  assign n27994 = n25742 & ~n27993;
  assign n27995 = n27965 & n27977;
  assign n27996 = ~n27994 & n27995;
  assign n27997 = ~n27887 & n27899;
  assign n27998 = ~n27943 & n27997;
  assign n27999 = n27958 & n27998;
  assign n28000 = n27996 & n27999;
  assign n28001 = n27634 & ~n28000;
  assign n28002 = ~n27881 & ~n27882;
  assign n4316 = n28001 | ~n28002;
  assign n28004 = P1_P3_INSTADDRPOINTER_REG_3_ & n27633;
  assign n28005 = P1_P3_REIP_REG_3_ & n27778;
  assign n28006 = ~P1_P3_INSTADDRPOINTER_REG_3_ & n27970;
  assign n28007 = P1_P3_INSTADDRPOINTER_REG_3_ & ~n27970;
  assign n28008 = ~n28006 & ~n28007;
  assign n28009 = n25938 & ~n28008;
  assign n28010 = n25781 & ~n28008;
  assign n28011 = ~n28009 & ~n28010;
  assign n28012 = ~n25828 & ~n28008;
  assign n28013 = P1_P3_INSTADDRPOINTER_REG_1_ & P1_P3_INSTADDRPOINTER_REG_2_;
  assign n28014 = ~P1_P3_INSTADDRPOINTER_REG_3_ & n28013;
  assign n28015 = P1_P3_INSTADDRPOINTER_REG_3_ & ~n28013;
  assign n28016 = ~n28014 & ~n28015;
  assign n28017 = n25899 & ~n28016;
  assign n28018 = n25900 & ~n28016;
  assign n28019 = n27642 & ~n28008;
  assign n28020 = n27645 & ~n28008;
  assign n28021 = ~n28019 & ~n28020;
  assign n28022 = n25715 & ~n28016;
  assign n28023 = n28021 & ~n28022;
  assign n28024 = ~n28017 & ~n28018;
  assign n28025 = n28023 & n28024;
  assign n28026 = ~n27950 & ~n27952;
  assign n28027 = ~n27953 & ~n28026;
  assign n28028 = P1_P3_INSTQUEUE_REG_0__3_ & n27652;
  assign n28029 = P1_P3_INSTQUEUE_REG_1__3_ & n27655;
  assign n28030 = P1_P3_INSTQUEUE_REG_2__3_ & n27658;
  assign n28031 = P1_P3_INSTQUEUE_REG_3__3_ & n27661;
  assign n28032 = ~n28028 & ~n28029;
  assign n28033 = ~n28030 & n28032;
  assign n28034 = ~n28031 & n28033;
  assign n28035 = P1_P3_INSTQUEUE_REG_4__3_ & n27667;
  assign n28036 = P1_P3_INSTQUEUE_REG_5__3_ & n27669;
  assign n28037 = P1_P3_INSTQUEUE_REG_6__3_ & n27671;
  assign n28038 = P1_P3_INSTQUEUE_REG_7__3_ & n27673;
  assign n28039 = ~n28035 & ~n28036;
  assign n28040 = ~n28037 & n28039;
  assign n28041 = ~n28038 & n28040;
  assign n28042 = P1_P3_INSTQUEUE_REG_8__3_ & n27679;
  assign n28043 = P1_P3_INSTQUEUE_REG_9__3_ & n27681;
  assign n28044 = P1_P3_INSTQUEUE_REG_10__3_ & n27683;
  assign n28045 = P1_P3_INSTQUEUE_REG_11__3_ & n27685;
  assign n28046 = ~n28042 & ~n28043;
  assign n28047 = ~n28044 & n28046;
  assign n28048 = ~n28045 & n28047;
  assign n28049 = P1_P3_INSTQUEUE_REG_12__3_ & n27691;
  assign n28050 = P1_P3_INSTQUEUE_REG_13__3_ & n27693;
  assign n28051 = P1_P3_INSTQUEUE_REG_14__3_ & n27695;
  assign n28052 = P1_P3_INSTQUEUE_REG_15__3_ & n27697;
  assign n28053 = ~n28049 & ~n28050;
  assign n28054 = ~n28051 & n28053;
  assign n28055 = ~n28052 & n28054;
  assign n28056 = n28034 & n28041;
  assign n28057 = n28048 & n28056;
  assign n28058 = n28055 & n28057;
  assign n28059 = ~n27822 & ~n27933;
  assign n28060 = n28058 & ~n28059;
  assign n28061 = ~n28058 & n28059;
  assign n28062 = ~n28060 & ~n28061;
  assign n28063 = ~P1_P3_INSTADDRPOINTER_REG_3_ & n28062;
  assign n28064 = P1_P3_INSTADDRPOINTER_REG_3_ & ~n28062;
  assign n28065 = ~n28063 & ~n28064;
  assign n28066 = n28027 & ~n28065;
  assign n28067 = P1_P3_INSTADDRPOINTER_REG_3_ & n28062;
  assign n28068 = ~P1_P3_INSTADDRPOINTER_REG_3_ & ~n28062;
  assign n28069 = ~n28067 & ~n28068;
  assign n28070 = ~n28027 & ~n28069;
  assign n28071 = ~n28066 & ~n28070;
  assign n28072 = n27739 & ~n28071;
  assign n28073 = ~n27902 & ~n27952;
  assign n28074 = ~n27953 & ~n28073;
  assign n28075 = n28058 & n28059;
  assign n28076 = ~n28058 & ~n28059;
  assign n28077 = ~n28075 & ~n28076;
  assign n28078 = ~P1_P3_INSTADDRPOINTER_REG_3_ & n28077;
  assign n28079 = ~n28074 & ~n28078;
  assign n28080 = P1_P3_INSTADDRPOINTER_REG_3_ & ~n28077;
  assign n28081 = n28079 & ~n28080;
  assign n28082 = ~P1_P3_INSTADDRPOINTER_REG_3_ & ~n28077;
  assign n28083 = P1_P3_INSTADDRPOINTER_REG_3_ & n28077;
  assign n28084 = ~n28082 & ~n28083;
  assign n28085 = n28074 & n28084;
  assign n28086 = ~n28081 & ~n28085;
  assign n28087 = n27741 & n28086;
  assign n28088 = ~n28072 & ~n28087;
  assign n28089 = n27758 & ~n28008;
  assign n28090 = n27751 & ~n28008;
  assign n28091 = n27747 & ~n28008;
  assign n28092 = n25785 & ~n28008;
  assign n28093 = ~n28089 & ~n28090;
  assign n28094 = ~n28091 & n28093;
  assign n28095 = ~n28092 & n28094;
  assign n28096 = n25641 & ~n28016;
  assign n28097 = n25719 & ~n28016;
  assign n28098 = n25723 & ~n28016;
  assign n28099 = ~P1_P3_INSTADDRPOINTER_REG_3_ & n27969;
  assign n28100 = P1_P3_INSTADDRPOINTER_REG_3_ & ~n27969;
  assign n28101 = ~n28099 & ~n28100;
  assign n28102 = n25739 & n28101;
  assign n28103 = n25731 & n28101;
  assign n28104 = ~n28096 & ~n28097;
  assign n28105 = ~n28098 & n28104;
  assign n28106 = ~n28102 & n28105;
  assign n28107 = ~n28103 & n28106;
  assign n28108 = n27987 & ~n27990;
  assign n28109 = n27979 & n28058;
  assign n28110 = ~n27979 & ~n28058;
  assign n28111 = ~n28109 & ~n28110;
  assign n28112 = P1_P3_INSTADDRPOINTER_REG_3_ & n28111;
  assign n28113 = ~n27989 & n28111;
  assign n28114 = P1_P3_INSTADDRPOINTER_REG_3_ & ~n27989;
  assign n28115 = ~n28113 & ~n28114;
  assign n28116 = ~n28108 & ~n28112;
  assign n28117 = ~n28115 & n28116;
  assign n28118 = ~P1_P3_INSTADDRPOINTER_REG_3_ & n28111;
  assign n28119 = P1_P3_INSTADDRPOINTER_REG_3_ & ~n28111;
  assign n28120 = ~n28118 & ~n28119;
  assign n28121 = ~n27990 & n28120;
  assign n28122 = ~n27987 & ~n27989;
  assign n28123 = n28121 & ~n28122;
  assign n28124 = ~n28117 & ~n28123;
  assign n28125 = n25742 & n28124;
  assign n28126 = n28095 & n28107;
  assign n28127 = ~n28125 & n28126;
  assign n28128 = n28011 & ~n28012;
  assign n28129 = n28025 & n28128;
  assign n28130 = n28088 & n28129;
  assign n28131 = n28127 & n28130;
  assign n28132 = n27634 & ~n28131;
  assign n28133 = ~n28004 & ~n28005;
  assign n4321 = n28132 | ~n28133;
  assign n28135 = P1_P3_INSTADDRPOINTER_REG_4_ & n27633;
  assign n28136 = P1_P3_REIP_REG_4_ & n27778;
  assign n28137 = P1_P3_INSTADDRPOINTER_REG_3_ & n27970;
  assign n28138 = ~P1_P3_INSTADDRPOINTER_REG_4_ & n28137;
  assign n28139 = P1_P3_INSTADDRPOINTER_REG_4_ & ~n28137;
  assign n28140 = ~n28138 & ~n28139;
  assign n28141 = ~n25828 & ~n28140;
  assign n28142 = P1_P3_INSTADDRPOINTER_REG_3_ & n28013;
  assign n28143 = ~P1_P3_INSTADDRPOINTER_REG_4_ & n28142;
  assign n28144 = P1_P3_INSTADDRPOINTER_REG_4_ & ~n28142;
  assign n28145 = ~n28143 & ~n28144;
  assign n28146 = n25899 & ~n28145;
  assign n28147 = n25900 & ~n28145;
  assign n28148 = n27642 & ~n28140;
  assign n28149 = n27645 & ~n28140;
  assign n28150 = ~n28148 & ~n28149;
  assign n28151 = n25715 & ~n28145;
  assign n28152 = n28150 & ~n28151;
  assign n28153 = ~n28146 & ~n28147;
  assign n28154 = n28152 & n28153;
  assign n28155 = P1_P3_INSTQUEUE_REG_0__4_ & n27652;
  assign n28156 = P1_P3_INSTQUEUE_REG_1__4_ & n27655;
  assign n28157 = P1_P3_INSTQUEUE_REG_2__4_ & n27658;
  assign n28158 = P1_P3_INSTQUEUE_REG_3__4_ & n27661;
  assign n28159 = ~n28155 & ~n28156;
  assign n28160 = ~n28157 & n28159;
  assign n28161 = ~n28158 & n28160;
  assign n28162 = P1_P3_INSTQUEUE_REG_4__4_ & n27667;
  assign n28163 = P1_P3_INSTQUEUE_REG_5__4_ & n27669;
  assign n28164 = P1_P3_INSTQUEUE_REG_6__4_ & n27671;
  assign n28165 = P1_P3_INSTQUEUE_REG_7__4_ & n27673;
  assign n28166 = ~n28162 & ~n28163;
  assign n28167 = ~n28164 & n28166;
  assign n28168 = ~n28165 & n28167;
  assign n28169 = P1_P3_INSTQUEUE_REG_8__4_ & n27679;
  assign n28170 = P1_P3_INSTQUEUE_REG_9__4_ & n27681;
  assign n28171 = P1_P3_INSTQUEUE_REG_10__4_ & n27683;
  assign n28172 = P1_P3_INSTQUEUE_REG_11__4_ & n27685;
  assign n28173 = ~n28169 & ~n28170;
  assign n28174 = ~n28171 & n28173;
  assign n28175 = ~n28172 & n28174;
  assign n28176 = P1_P3_INSTQUEUE_REG_12__4_ & n27691;
  assign n28177 = P1_P3_INSTQUEUE_REG_13__4_ & n27693;
  assign n28178 = P1_P3_INSTQUEUE_REG_14__4_ & n27695;
  assign n28179 = P1_P3_INSTQUEUE_REG_15__4_ & n27697;
  assign n28180 = ~n28176 & ~n28177;
  assign n28181 = ~n28178 & n28180;
  assign n28182 = ~n28179 & n28181;
  assign n28183 = n28161 & n28168;
  assign n28184 = n28175 & n28183;
  assign n28185 = n28182 & n28184;
  assign n28186 = n28061 & n28185;
  assign n28187 = ~n28061 & ~n28185;
  assign n28188 = ~n28186 & ~n28187;
  assign n28189 = P1_P3_INSTADDRPOINTER_REG_4_ & ~n28188;
  assign n28190 = ~P1_P3_INSTADDRPOINTER_REG_4_ & n28188;
  assign n28191 = ~n28189 & ~n28190;
  assign n28192 = ~n28079 & ~n28080;
  assign n28193 = n28191 & ~n28192;
  assign n28194 = ~P1_P3_INSTADDRPOINTER_REG_4_ & ~n28188;
  assign n28195 = P1_P3_INSTADDRPOINTER_REG_4_ & n28188;
  assign n28196 = ~n28194 & ~n28195;
  assign n28197 = ~n28080 & n28196;
  assign n28198 = ~n28079 & n28197;
  assign n28199 = ~n28193 & ~n28198;
  assign n28200 = n27741 & n28199;
  assign n28201 = n25938 & ~n28140;
  assign n28202 = n25781 & ~n28140;
  assign n28203 = ~n28201 & ~n28202;
  assign n28204 = ~n27952 & ~n28068;
  assign n28205 = ~n27947 & ~n27948;
  assign n28206 = ~n27953 & n28205;
  assign n28207 = ~n27826 & n28206;
  assign n28208 = n28204 & ~n28207;
  assign n28209 = ~n28067 & ~n28208;
  assign n28210 = n28061 & ~n28185;
  assign n28211 = ~n28061 & n28185;
  assign n28212 = ~n28210 & ~n28211;
  assign n28213 = ~P1_P3_INSTADDRPOINTER_REG_4_ & n28212;
  assign n28214 = P1_P3_INSTADDRPOINTER_REG_4_ & ~n28212;
  assign n28215 = ~n28213 & ~n28214;
  assign n28216 = n28209 & ~n28215;
  assign n28217 = P1_P3_INSTADDRPOINTER_REG_4_ & n28212;
  assign n28218 = ~P1_P3_INSTADDRPOINTER_REG_4_ & ~n28212;
  assign n28219 = ~n28217 & ~n28218;
  assign n28220 = ~n28209 & ~n28219;
  assign n28221 = ~n28216 & ~n28220;
  assign n28222 = n27739 & ~n28221;
  assign n28223 = n28203 & ~n28222;
  assign n28224 = n27758 & ~n28140;
  assign n28225 = n27751 & ~n28140;
  assign n28226 = n27747 & ~n28140;
  assign n28227 = n25785 & ~n28140;
  assign n28228 = ~n28224 & ~n28225;
  assign n28229 = ~n28226 & n28228;
  assign n28230 = ~n28227 & n28229;
  assign n28231 = n25641 & ~n28145;
  assign n28232 = n25719 & ~n28145;
  assign n28233 = n25723 & ~n28145;
  assign n28234 = ~P1_P3_INSTADDRPOINTER_REG_4_ & n28100;
  assign n28235 = P1_P3_INSTADDRPOINTER_REG_4_ & ~n28100;
  assign n28236 = ~n28234 & ~n28235;
  assign n28237 = n25739 & ~n28236;
  assign n28238 = n25731 & ~n28236;
  assign n28239 = ~n28231 & ~n28232;
  assign n28240 = ~n28233 & n28239;
  assign n28241 = ~n28237 & n28240;
  assign n28242 = ~n28238 & n28241;
  assign n28243 = n28110 & n28185;
  assign n28244 = ~n28110 & ~n28185;
  assign n28245 = ~n28243 & ~n28244;
  assign n28246 = ~P1_P3_INSTADDRPOINTER_REG_4_ & ~n28245;
  assign n28247 = P1_P3_INSTADDRPOINTER_REG_4_ & n28245;
  assign n28248 = ~n28246 & ~n28247;
  assign n28249 = n27990 & n28111;
  assign n28250 = ~n27990 & ~n28111;
  assign n28251 = P1_P3_INSTADDRPOINTER_REG_3_ & ~n28250;
  assign n28252 = ~n28249 & ~n28251;
  assign n28253 = ~n27987 & ~n28115;
  assign n28254 = n28252 & ~n28253;
  assign n28255 = ~n28248 & n28254;
  assign n28256 = ~P1_P3_INSTADDRPOINTER_REG_4_ & n28245;
  assign n28257 = P1_P3_INSTADDRPOINTER_REG_4_ & ~n28245;
  assign n28258 = ~n28256 & ~n28257;
  assign n28259 = ~n28254 & ~n28258;
  assign n28260 = ~n28255 & ~n28259;
  assign n28261 = n25742 & ~n28260;
  assign n28262 = n28230 & n28242;
  assign n28263 = ~n28261 & n28262;
  assign n28264 = ~n28141 & n28154;
  assign n28265 = ~n28200 & n28264;
  assign n28266 = n28223 & n28265;
  assign n28267 = n28263 & n28266;
  assign n28268 = n27634 & ~n28267;
  assign n28269 = ~n28135 & ~n28136;
  assign n4326 = n28268 | ~n28269;
  assign n28271 = P1_P3_INSTADDRPOINTER_REG_5_ & n27633;
  assign n28272 = P1_P3_REIP_REG_5_ & n27778;
  assign n28273 = P1_P3_INSTADDRPOINTER_REG_4_ & n28142;
  assign n28274 = ~P1_P3_INSTADDRPOINTER_REG_5_ & n28273;
  assign n28275 = P1_P3_INSTADDRPOINTER_REG_5_ & ~n28273;
  assign n28276 = ~n28274 & ~n28275;
  assign n28277 = n25899 & ~n28276;
  assign n28278 = n25900 & ~n28276;
  assign n28279 = P1_P3_INSTADDRPOINTER_REG_4_ & n28137;
  assign n28280 = ~P1_P3_INSTADDRPOINTER_REG_5_ & n28279;
  assign n28281 = P1_P3_INSTADDRPOINTER_REG_5_ & ~n28279;
  assign n28282 = ~n28280 & ~n28281;
  assign n28283 = n27642 & ~n28282;
  assign n28284 = n27645 & ~n28282;
  assign n28285 = ~n28283 & ~n28284;
  assign n28286 = n25715 & ~n28276;
  assign n28287 = n28285 & ~n28286;
  assign n28288 = ~n28277 & ~n28278;
  assign n28289 = n28287 & n28288;
  assign n28290 = ~n25828 & ~n28282;
  assign n28291 = n28067 & ~n28218;
  assign n28292 = ~n28217 & ~n28291;
  assign n28293 = n28204 & ~n28218;
  assign n28294 = ~n28207 & n28293;
  assign n28295 = n28292 & ~n28294;
  assign n28296 = P1_P3_INSTQUEUE_REG_0__5_ & n27652;
  assign n28297 = P1_P3_INSTQUEUE_REG_1__5_ & n27655;
  assign n28298 = P1_P3_INSTQUEUE_REG_2__5_ & n27658;
  assign n28299 = P1_P3_INSTQUEUE_REG_3__5_ & n27661;
  assign n28300 = ~n28296 & ~n28297;
  assign n28301 = ~n28298 & n28300;
  assign n28302 = ~n28299 & n28301;
  assign n28303 = P1_P3_INSTQUEUE_REG_4__5_ & n27667;
  assign n28304 = P1_P3_INSTQUEUE_REG_5__5_ & n27669;
  assign n28305 = P1_P3_INSTQUEUE_REG_6__5_ & n27671;
  assign n28306 = P1_P3_INSTQUEUE_REG_7__5_ & n27673;
  assign n28307 = ~n28303 & ~n28304;
  assign n28308 = ~n28305 & n28307;
  assign n28309 = ~n28306 & n28308;
  assign n28310 = P1_P3_INSTQUEUE_REG_8__5_ & n27679;
  assign n28311 = P1_P3_INSTQUEUE_REG_9__5_ & n27681;
  assign n28312 = P1_P3_INSTQUEUE_REG_10__5_ & n27683;
  assign n28313 = P1_P3_INSTQUEUE_REG_11__5_ & n27685;
  assign n28314 = ~n28310 & ~n28311;
  assign n28315 = ~n28312 & n28314;
  assign n28316 = ~n28313 & n28315;
  assign n28317 = P1_P3_INSTQUEUE_REG_12__5_ & n27691;
  assign n28318 = P1_P3_INSTQUEUE_REG_13__5_ & n27693;
  assign n28319 = P1_P3_INSTQUEUE_REG_14__5_ & n27695;
  assign n28320 = P1_P3_INSTQUEUE_REG_15__5_ & n27697;
  assign n28321 = ~n28317 & ~n28318;
  assign n28322 = ~n28319 & n28321;
  assign n28323 = ~n28320 & n28322;
  assign n28324 = n28302 & n28309;
  assign n28325 = n28316 & n28324;
  assign n28326 = n28323 & n28325;
  assign n28327 = ~n28210 & n28326;
  assign n28328 = ~n28185 & ~n28326;
  assign n28329 = n28061 & n28328;
  assign n28330 = ~n28327 & ~n28329;
  assign n28331 = ~P1_P3_INSTADDRPOINTER_REG_5_ & n28330;
  assign n28332 = P1_P3_INSTADDRPOINTER_REG_5_ & ~n28330;
  assign n28333 = ~n28331 & ~n28332;
  assign n28334 = n28295 & ~n28333;
  assign n28335 = ~n28295 & n28333;
  assign n28336 = ~n28334 & ~n28335;
  assign n28337 = n27739 & ~n28336;
  assign n28338 = n25938 & ~n28282;
  assign n28339 = n25781 & ~n28282;
  assign n28340 = ~n28338 & ~n28339;
  assign n28341 = n28080 & ~n28190;
  assign n28342 = ~n28189 & ~n28341;
  assign n28343 = ~n28078 & ~n28190;
  assign n28344 = ~n28074 & n28343;
  assign n28345 = n28342 & ~n28344;
  assign n28346 = n28210 & n28326;
  assign n28347 = ~n28210 & ~n28326;
  assign n28348 = ~n28346 & ~n28347;
  assign n28349 = ~P1_P3_INSTADDRPOINTER_REG_5_ & ~n28348;
  assign n28350 = P1_P3_INSTADDRPOINTER_REG_5_ & n28348;
  assign n28351 = ~n28349 & ~n28350;
  assign n28352 = n28345 & ~n28351;
  assign n28353 = ~n28345 & n28351;
  assign n28354 = ~n28352 & ~n28353;
  assign n28355 = n27741 & ~n28354;
  assign n28356 = n28340 & ~n28355;
  assign n28357 = n27758 & ~n28282;
  assign n28358 = n27751 & ~n28282;
  assign n28359 = n27747 & ~n28282;
  assign n28360 = n25785 & ~n28282;
  assign n28361 = ~n28357 & ~n28358;
  assign n28362 = ~n28359 & n28361;
  assign n28363 = ~n28360 & n28362;
  assign n28364 = n25641 & ~n28276;
  assign n28365 = n25719 & ~n28276;
  assign n28366 = n25723 & ~n28276;
  assign n28367 = P1_P3_INSTADDRPOINTER_REG_4_ & n28100;
  assign n28368 = ~P1_P3_INSTADDRPOINTER_REG_5_ & n28367;
  assign n28369 = P1_P3_INSTADDRPOINTER_REG_5_ & ~n28367;
  assign n28370 = ~n28368 & ~n28369;
  assign n28371 = n25739 & ~n28370;
  assign n28372 = n25731 & ~n28370;
  assign n28373 = ~n28364 & ~n28365;
  assign n28374 = ~n28366 & n28373;
  assign n28375 = ~n28371 & n28374;
  assign n28376 = ~n28372 & n28375;
  assign n28377 = n28110 & ~n28185;
  assign n28378 = n28326 & n28377;
  assign n28379 = ~n28326 & ~n28377;
  assign n28380 = ~n28378 & ~n28379;
  assign n28381 = P1_P3_INSTADDRPOINTER_REG_5_ & ~n28380;
  assign n28382 = ~P1_P3_INSTADDRPOINTER_REG_5_ & n28380;
  assign n28383 = ~n28256 & ~n28382;
  assign n28384 = ~n28381 & n28383;
  assign n28385 = n28254 & ~n28257;
  assign n28386 = n28384 & ~n28385;
  assign n28387 = ~P1_P3_INSTADDRPOINTER_REG_5_ & ~n28380;
  assign n28388 = P1_P3_INSTADDRPOINTER_REG_5_ & n28380;
  assign n28389 = ~n28387 & ~n28388;
  assign n28390 = ~n28257 & n28389;
  assign n28391 = ~n28254 & ~n28256;
  assign n28392 = n28390 & ~n28391;
  assign n28393 = ~n28386 & ~n28392;
  assign n28394 = n25742 & n28393;
  assign n28395 = n28363 & n28376;
  assign n28396 = ~n28394 & n28395;
  assign n28397 = n28289 & ~n28290;
  assign n28398 = ~n28337 & n28397;
  assign n28399 = n28356 & n28398;
  assign n28400 = n28396 & n28399;
  assign n28401 = n27634 & ~n28400;
  assign n28402 = ~n28271 & ~n28272;
  assign n4331 = n28401 | ~n28402;
  assign n28404 = P1_P3_INSTADDRPOINTER_REG_6_ & n27633;
  assign n28405 = P1_P3_REIP_REG_6_ & n27778;
  assign n28406 = P1_P3_INSTADDRPOINTER_REG_5_ & n28273;
  assign n28407 = ~P1_P3_INSTADDRPOINTER_REG_6_ & n28406;
  assign n28408 = P1_P3_INSTADDRPOINTER_REG_6_ & ~n28406;
  assign n28409 = ~n28407 & ~n28408;
  assign n28410 = n25899 & ~n28409;
  assign n28411 = n25900 & ~n28409;
  assign n28412 = P1_P3_INSTADDRPOINTER_REG_5_ & n28279;
  assign n28413 = ~P1_P3_INSTADDRPOINTER_REG_6_ & n28412;
  assign n28414 = P1_P3_INSTADDRPOINTER_REG_6_ & ~n28412;
  assign n28415 = ~n28413 & ~n28414;
  assign n28416 = n27642 & ~n28415;
  assign n28417 = n27645 & ~n28415;
  assign n28418 = ~n28416 & ~n28417;
  assign n28419 = n25715 & ~n28409;
  assign n28420 = n28418 & ~n28419;
  assign n28421 = ~n28410 & ~n28411;
  assign n28422 = n28420 & n28421;
  assign n28423 = ~n25828 & ~n28415;
  assign n28424 = ~P1_P3_INSTADDRPOINTER_REG_5_ & ~n28330;
  assign n28425 = ~n28295 & ~n28424;
  assign n28426 = P1_P3_INSTADDRPOINTER_REG_5_ & n28330;
  assign n28427 = ~n28425 & ~n28426;
  assign n28428 = P1_P3_INSTQUEUE_REG_0__6_ & n27652;
  assign n28429 = P1_P3_INSTQUEUE_REG_1__6_ & n27655;
  assign n28430 = P1_P3_INSTQUEUE_REG_2__6_ & n27658;
  assign n28431 = P1_P3_INSTQUEUE_REG_3__6_ & n27661;
  assign n28432 = ~n28428 & ~n28429;
  assign n28433 = ~n28430 & n28432;
  assign n28434 = ~n28431 & n28433;
  assign n28435 = P1_P3_INSTQUEUE_REG_4__6_ & n27667;
  assign n28436 = P1_P3_INSTQUEUE_REG_5__6_ & n27669;
  assign n28437 = P1_P3_INSTQUEUE_REG_6__6_ & n27671;
  assign n28438 = P1_P3_INSTQUEUE_REG_7__6_ & n27673;
  assign n28439 = ~n28435 & ~n28436;
  assign n28440 = ~n28437 & n28439;
  assign n28441 = ~n28438 & n28440;
  assign n28442 = P1_P3_INSTQUEUE_REG_8__6_ & n27679;
  assign n28443 = P1_P3_INSTQUEUE_REG_9__6_ & n27681;
  assign n28444 = P1_P3_INSTQUEUE_REG_10__6_ & n27683;
  assign n28445 = P1_P3_INSTQUEUE_REG_11__6_ & n27685;
  assign n28446 = ~n28442 & ~n28443;
  assign n28447 = ~n28444 & n28446;
  assign n28448 = ~n28445 & n28447;
  assign n28449 = P1_P3_INSTQUEUE_REG_12__6_ & n27691;
  assign n28450 = P1_P3_INSTQUEUE_REG_13__6_ & n27693;
  assign n28451 = P1_P3_INSTQUEUE_REG_14__6_ & n27695;
  assign n28452 = P1_P3_INSTQUEUE_REG_15__6_ & n27697;
  assign n28453 = ~n28449 & ~n28450;
  assign n28454 = ~n28451 & n28453;
  assign n28455 = ~n28452 & n28454;
  assign n28456 = n28434 & n28441;
  assign n28457 = n28448 & n28456;
  assign n28458 = n28455 & n28457;
  assign n28459 = n28329 & ~n28458;
  assign n28460 = ~n28329 & n28458;
  assign n28461 = ~n28459 & ~n28460;
  assign n28462 = ~P1_P3_INSTADDRPOINTER_REG_6_ & n28461;
  assign n28463 = P1_P3_INSTADDRPOINTER_REG_6_ & ~n28461;
  assign n28464 = ~n28462 & ~n28463;
  assign n28465 = n28427 & ~n28464;
  assign n28466 = ~n28427 & n28464;
  assign n28467 = ~n28465 & ~n28466;
  assign n28468 = n27739 & ~n28467;
  assign n28469 = n25938 & ~n28415;
  assign n28470 = n25781 & ~n28415;
  assign n28471 = ~n28469 & ~n28470;
  assign n28472 = ~n28345 & ~n28348;
  assign n28473 = P1_P3_INSTADDRPOINTER_REG_5_ & ~n28345;
  assign n28474 = P1_P3_INSTADDRPOINTER_REG_5_ & ~n28348;
  assign n28475 = ~n28472 & ~n28473;
  assign n28476 = ~n28474 & n28475;
  assign n28477 = n28210 & ~n28326;
  assign n28478 = n28458 & n28477;
  assign n28479 = ~n28458 & ~n28477;
  assign n28480 = ~n28478 & ~n28479;
  assign n28481 = ~P1_P3_INSTADDRPOINTER_REG_6_ & ~n28480;
  assign n28482 = P1_P3_INSTADDRPOINTER_REG_6_ & n28480;
  assign n28483 = ~n28481 & ~n28482;
  assign n28484 = n28476 & ~n28483;
  assign n28485 = ~n28476 & n28483;
  assign n28486 = ~n28484 & ~n28485;
  assign n28487 = n27741 & ~n28486;
  assign n28488 = n28471 & ~n28487;
  assign n28489 = n27758 & ~n28415;
  assign n28490 = n27751 & ~n28415;
  assign n28491 = n27747 & ~n28415;
  assign n28492 = n25785 & ~n28415;
  assign n28493 = ~n28489 & ~n28490;
  assign n28494 = ~n28491 & n28493;
  assign n28495 = ~n28492 & n28494;
  assign n28496 = n25641 & ~n28409;
  assign n28497 = n25719 & ~n28409;
  assign n28498 = n25723 & ~n28409;
  assign n28499 = P1_P3_INSTADDRPOINTER_REG_5_ & n28367;
  assign n28500 = ~P1_P3_INSTADDRPOINTER_REG_6_ & n28499;
  assign n28501 = P1_P3_INSTADDRPOINTER_REG_6_ & ~n28499;
  assign n28502 = ~n28500 & ~n28501;
  assign n28503 = n25739 & ~n28502;
  assign n28504 = n25731 & ~n28502;
  assign n28505 = ~n28496 & ~n28497;
  assign n28506 = ~n28498 & n28505;
  assign n28507 = ~n28503 & n28506;
  assign n28508 = ~n28504 & n28507;
  assign n28509 = n28257 & ~n28380;
  assign n28510 = ~n28257 & n28380;
  assign n28511 = P1_P3_INSTADDRPOINTER_REG_5_ & ~n28510;
  assign n28512 = ~n28509 & ~n28511;
  assign n28513 = ~n28254 & n28383;
  assign n28514 = n28512 & ~n28513;
  assign n28515 = ~n28326 & n28377;
  assign n28516 = n28458 & n28515;
  assign n28517 = ~n28458 & ~n28515;
  assign n28518 = ~n28516 & ~n28517;
  assign n28519 = ~P1_P3_INSTADDRPOINTER_REG_6_ & ~n28518;
  assign n28520 = P1_P3_INSTADDRPOINTER_REG_6_ & n28518;
  assign n28521 = ~n28519 & ~n28520;
  assign n28522 = n28514 & ~n28521;
  assign n28523 = ~n28514 & n28521;
  assign n28524 = ~n28522 & ~n28523;
  assign n28525 = n25742 & ~n28524;
  assign n28526 = n28495 & n28508;
  assign n28527 = ~n28525 & n28526;
  assign n28528 = n28422 & ~n28423;
  assign n28529 = ~n28468 & n28528;
  assign n28530 = n28488 & n28529;
  assign n28531 = n28527 & n28530;
  assign n28532 = n27634 & ~n28531;
  assign n28533 = ~n28404 & ~n28405;
  assign n4336 = n28532 | ~n28533;
  assign n28535 = P1_P3_INSTADDRPOINTER_REG_7_ & n27633;
  assign n28536 = P1_P3_REIP_REG_7_ & n27778;
  assign n28537 = P1_P3_INSTADDRPOINTER_REG_6_ & n28406;
  assign n28538 = ~P1_P3_INSTADDRPOINTER_REG_7_ & n28537;
  assign n28539 = P1_P3_INSTADDRPOINTER_REG_7_ & ~n28537;
  assign n28540 = ~n28538 & ~n28539;
  assign n28541 = n25899 & ~n28540;
  assign n28542 = n25900 & ~n28540;
  assign n28543 = P1_P3_INSTADDRPOINTER_REG_6_ & n28412;
  assign n28544 = ~P1_P3_INSTADDRPOINTER_REG_7_ & n28543;
  assign n28545 = P1_P3_INSTADDRPOINTER_REG_7_ & ~n28543;
  assign n28546 = ~n28544 & ~n28545;
  assign n28547 = n27642 & ~n28546;
  assign n28548 = n27645 & ~n28546;
  assign n28549 = ~n28547 & ~n28548;
  assign n28550 = n25715 & ~n28540;
  assign n28551 = n28549 & ~n28550;
  assign n28552 = ~n28541 & ~n28542;
  assign n28553 = n28551 & n28552;
  assign n28554 = ~n25828 & ~n28546;
  assign n28555 = P1_P3_INSTADDRPOINTER_REG_6_ & n28461;
  assign n28556 = ~P1_P3_INSTADDRPOINTER_REG_6_ & ~n28461;
  assign n28557 = ~n28427 & ~n28556;
  assign n28558 = ~n28555 & ~n28557;
  assign n28559 = n27738 & ~n28459;
  assign n28560 = ~n27738 & ~n28458;
  assign n28561 = n28329 & n28560;
  assign n28562 = ~n28559 & ~n28561;
  assign n28563 = ~P1_P3_INSTADDRPOINTER_REG_7_ & n28562;
  assign n28564 = P1_P3_INSTADDRPOINTER_REG_7_ & ~n28562;
  assign n28565 = ~n28563 & ~n28564;
  assign n28566 = n28558 & ~n28565;
  assign n28567 = ~n28558 & n28565;
  assign n28568 = ~n28566 & ~n28567;
  assign n28569 = n27739 & ~n28568;
  assign n28570 = n25938 & ~n28546;
  assign n28571 = n25781 & ~n28546;
  assign n28572 = ~n28570 & ~n28571;
  assign n28573 = P1_P3_INSTADDRPOINTER_REG_6_ & ~n28480;
  assign n28574 = ~P1_P3_INSTADDRPOINTER_REG_6_ & n28480;
  assign n28575 = ~n28476 & ~n28574;
  assign n28576 = ~n28573 & ~n28575;
  assign n28577 = ~n28458 & n28477;
  assign n28578 = n27738 & n28577;
  assign n28579 = ~n27738 & ~n28577;
  assign n28580 = ~n28578 & ~n28579;
  assign n28581 = ~P1_P3_INSTADDRPOINTER_REG_7_ & ~n28580;
  assign n28582 = P1_P3_INSTADDRPOINTER_REG_7_ & n28580;
  assign n28583 = ~n28581 & ~n28582;
  assign n28584 = n28576 & ~n28583;
  assign n28585 = ~n28576 & n28583;
  assign n28586 = ~n28584 & ~n28585;
  assign n28587 = n27741 & ~n28586;
  assign n28588 = n28572 & ~n28587;
  assign n28589 = n27758 & ~n28546;
  assign n28590 = n27751 & ~n28546;
  assign n28591 = n27747 & ~n28546;
  assign n28592 = n25785 & ~n28546;
  assign n28593 = ~n28589 & ~n28590;
  assign n28594 = ~n28591 & n28593;
  assign n28595 = ~n28592 & n28594;
  assign n28596 = n25641 & ~n28540;
  assign n28597 = n25719 & ~n28540;
  assign n28598 = n25723 & ~n28540;
  assign n28599 = P1_P3_INSTADDRPOINTER_REG_6_ & n28499;
  assign n28600 = ~P1_P3_INSTADDRPOINTER_REG_7_ & n28599;
  assign n28601 = P1_P3_INSTADDRPOINTER_REG_7_ & ~n28599;
  assign n28602 = ~n28600 & ~n28601;
  assign n28603 = n25739 & ~n28602;
  assign n28604 = n25731 & ~n28602;
  assign n28605 = ~n28596 & ~n28597;
  assign n28606 = ~n28598 & n28605;
  assign n28607 = ~n28603 & n28606;
  assign n28608 = ~n28604 & n28607;
  assign n28609 = P1_P3_INSTADDRPOINTER_REG_6_ & ~n28518;
  assign n28610 = ~P1_P3_INSTADDRPOINTER_REG_6_ & n28518;
  assign n28611 = ~n28514 & ~n28610;
  assign n28612 = ~n28609 & ~n28611;
  assign n28613 = ~n28458 & n28515;
  assign n28614 = n27738 & n28613;
  assign n28615 = ~n27738 & ~n28613;
  assign n28616 = ~n28614 & ~n28615;
  assign n28617 = ~P1_P3_INSTADDRPOINTER_REG_7_ & ~n28616;
  assign n28618 = P1_P3_INSTADDRPOINTER_REG_7_ & n28616;
  assign n28619 = ~n28617 & ~n28618;
  assign n28620 = n28612 & ~n28619;
  assign n28621 = ~n28612 & n28619;
  assign n28622 = ~n28620 & ~n28621;
  assign n28623 = n25742 & ~n28622;
  assign n28624 = n28595 & n28608;
  assign n28625 = ~n28623 & n28624;
  assign n28626 = n28553 & ~n28554;
  assign n28627 = ~n28569 & n28626;
  assign n28628 = n28588 & n28627;
  assign n28629 = n28625 & n28628;
  assign n28630 = n27634 & ~n28629;
  assign n28631 = ~n28535 & ~n28536;
  assign n4341 = n28630 | ~n28631;
  assign n28633 = P1_P3_INSTADDRPOINTER_REG_8_ & n27633;
  assign n28634 = P1_P3_REIP_REG_8_ & n27778;
  assign n28635 = P1_P3_INSTADDRPOINTER_REG_7_ & n28537;
  assign n28636 = ~P1_P3_INSTADDRPOINTER_REG_8_ & n28635;
  assign n28637 = P1_P3_INSTADDRPOINTER_REG_8_ & ~n28635;
  assign n28638 = ~n28636 & ~n28637;
  assign n28639 = n25899 & ~n28638;
  assign n28640 = n25900 & ~n28638;
  assign n28641 = n25715 & ~n28638;
  assign n28642 = P1_P3_INSTADDRPOINTER_REG_7_ & n28543;
  assign n28643 = ~P1_P3_INSTADDRPOINTER_REG_8_ & n28642;
  assign n28644 = P1_P3_INSTADDRPOINTER_REG_8_ & ~n28642;
  assign n28645 = ~n28643 & ~n28644;
  assign n28646 = n27645 & ~n28645;
  assign n28647 = n27642 & ~n28645;
  assign n28648 = ~n28641 & ~n28646;
  assign n28649 = ~n28647 & n28648;
  assign n28650 = ~n28639 & ~n28640;
  assign n28651 = n28649 & n28650;
  assign n28652 = ~n25828 & ~n28645;
  assign n28653 = ~P1_P3_INSTADDRPOINTER_REG_7_ & ~n28562;
  assign n28654 = ~n28558 & ~n28653;
  assign n28655 = P1_P3_INSTADDRPOINTER_REG_7_ & n28562;
  assign n28656 = ~n28654 & ~n28655;
  assign n28657 = P1_P3_INSTADDRPOINTER_REG_8_ & n28561;
  assign n28658 = ~P1_P3_INSTADDRPOINTER_REG_8_ & ~n28561;
  assign n28659 = ~n28657 & ~n28658;
  assign n28660 = n28656 & ~n28659;
  assign n28661 = ~n28656 & n28659;
  assign n28662 = ~n28660 & ~n28661;
  assign n28663 = n27739 & ~n28662;
  assign n28664 = n25938 & ~n28645;
  assign n28665 = n25781 & ~n28645;
  assign n28666 = ~n28664 & ~n28665;
  assign n28667 = ~n28576 & ~n28580;
  assign n28668 = P1_P3_INSTADDRPOINTER_REG_7_ & ~n28576;
  assign n28669 = P1_P3_INSTADDRPOINTER_REG_7_ & ~n28580;
  assign n28670 = ~n28667 & ~n28668;
  assign n28671 = ~n28669 & n28670;
  assign n28672 = n28477 & n28560;
  assign n28673 = ~P1_P3_INSTADDRPOINTER_REG_8_ & n28672;
  assign n28674 = P1_P3_INSTADDRPOINTER_REG_8_ & ~n28672;
  assign n28675 = ~n28673 & ~n28674;
  assign n28676 = n28671 & ~n28675;
  assign n28677 = ~n28671 & n28675;
  assign n28678 = ~n28676 & ~n28677;
  assign n28679 = n27741 & ~n28678;
  assign n28680 = n28666 & ~n28679;
  assign n28681 = n27758 & ~n28645;
  assign n28682 = n25785 & ~n28645;
  assign n28683 = n27747 & ~n28645;
  assign n28684 = n27751 & ~n28645;
  assign n28685 = ~n28681 & ~n28682;
  assign n28686 = ~n28683 & n28685;
  assign n28687 = ~n28684 & n28686;
  assign n28688 = n25641 & ~n28638;
  assign n28689 = n25719 & ~n28638;
  assign n28690 = n25723 & ~n28638;
  assign n28691 = P1_P3_INSTADDRPOINTER_REG_7_ & n28599;
  assign n28692 = ~P1_P3_INSTADDRPOINTER_REG_8_ & n28691;
  assign n28693 = P1_P3_INSTADDRPOINTER_REG_8_ & ~n28691;
  assign n28694 = ~n28692 & ~n28693;
  assign n28695 = n25739 & ~n28694;
  assign n28696 = n25731 & ~n28694;
  assign n28697 = ~n28688 & ~n28689;
  assign n28698 = ~n28690 & n28697;
  assign n28699 = ~n28695 & n28698;
  assign n28700 = ~n28696 & n28699;
  assign n28701 = ~n28612 & ~n28616;
  assign n28702 = P1_P3_INSTADDRPOINTER_REG_7_ & ~n28612;
  assign n28703 = P1_P3_INSTADDRPOINTER_REG_7_ & ~n28616;
  assign n28704 = ~n28701 & ~n28702;
  assign n28705 = ~n28703 & n28704;
  assign n28706 = n28515 & n28560;
  assign n28707 = ~P1_P3_INSTADDRPOINTER_REG_8_ & n28706;
  assign n28708 = P1_P3_INSTADDRPOINTER_REG_8_ & ~n28706;
  assign n28709 = ~n28707 & ~n28708;
  assign n28710 = n28705 & ~n28709;
  assign n28711 = ~n28705 & n28709;
  assign n28712 = ~n28710 & ~n28711;
  assign n28713 = n25742 & ~n28712;
  assign n28714 = n28687 & n28700;
  assign n28715 = ~n28713 & n28714;
  assign n28716 = n28651 & ~n28652;
  assign n28717 = ~n28663 & n28716;
  assign n28718 = n28680 & n28717;
  assign n28719 = n28715 & n28718;
  assign n28720 = n27634 & ~n28719;
  assign n28721 = ~n28633 & ~n28634;
  assign n4346 = n28720 | ~n28721;
  assign n28723 = P1_P3_INSTADDRPOINTER_REG_9_ & n27633;
  assign n28724 = P1_P3_REIP_REG_9_ & n27778;
  assign n28725 = P1_P3_INSTADDRPOINTER_REG_8_ & n28635;
  assign n28726 = ~P1_P3_INSTADDRPOINTER_REG_9_ & n28725;
  assign n28727 = P1_P3_INSTADDRPOINTER_REG_9_ & ~n28725;
  assign n28728 = ~n28726 & ~n28727;
  assign n28729 = n25899 & ~n28728;
  assign n28730 = n25900 & ~n28728;
  assign n28731 = P1_P3_INSTADDRPOINTER_REG_8_ & n28642;
  assign n28732 = ~P1_P3_INSTADDRPOINTER_REG_9_ & n28731;
  assign n28733 = P1_P3_INSTADDRPOINTER_REG_9_ & ~n28731;
  assign n28734 = ~n28732 & ~n28733;
  assign n28735 = n27642 & ~n28734;
  assign n28736 = n25715 & ~n28728;
  assign n28737 = n27645 & ~n28734;
  assign n28738 = ~n28736 & ~n28737;
  assign n28739 = ~n28729 & ~n28730;
  assign n28740 = ~n28735 & n28739;
  assign n28741 = n28738 & n28740;
  assign n28742 = ~n25828 & ~n28734;
  assign n28743 = P1_P3_INSTADDRPOINTER_REG_8_ & ~n28656;
  assign n28744 = ~n28561 & ~n28656;
  assign n28745 = P1_P3_INSTADDRPOINTER_REG_8_ & ~n28561;
  assign n28746 = ~n28743 & ~n28744;
  assign n28747 = ~n28745 & n28746;
  assign n28748 = P1_P3_INSTADDRPOINTER_REG_9_ & n28561;
  assign n28749 = ~P1_P3_INSTADDRPOINTER_REG_9_ & ~n28561;
  assign n28750 = ~n28748 & ~n28749;
  assign n28751 = n28747 & ~n28750;
  assign n28752 = P1_P3_INSTADDRPOINTER_REG_9_ & ~n28561;
  assign n28753 = ~P1_P3_INSTADDRPOINTER_REG_9_ & n28561;
  assign n28754 = ~n28752 & ~n28753;
  assign n28755 = ~n28747 & ~n28754;
  assign n28756 = ~n28751 & ~n28755;
  assign n28757 = n27739 & ~n28756;
  assign n28758 = n25938 & ~n28734;
  assign n28759 = n25781 & ~n28734;
  assign n28760 = ~n28758 & ~n28759;
  assign n28761 = P1_P3_INSTADDRPOINTER_REG_8_ & n28672;
  assign n28762 = ~P1_P3_INSTADDRPOINTER_REG_8_ & ~n28672;
  assign n28763 = ~n28671 & ~n28762;
  assign n28764 = ~n28761 & ~n28763;
  assign n28765 = ~P1_P3_INSTADDRPOINTER_REG_9_ & n28764;
  assign n28766 = P1_P3_INSTADDRPOINTER_REG_9_ & ~n28764;
  assign n28767 = ~n28765 & ~n28766;
  assign n28768 = n27741 & n28767;
  assign n28769 = n28760 & ~n28768;
  assign n28770 = n27758 & ~n28734;
  assign n28771 = n25785 & ~n28734;
  assign n28772 = n27747 & ~n28734;
  assign n28773 = n27751 & ~n28734;
  assign n28774 = ~n28770 & ~n28771;
  assign n28775 = ~n28772 & n28774;
  assign n28776 = ~n28773 & n28775;
  assign n28777 = n25641 & ~n28728;
  assign n28778 = n25719 & ~n28728;
  assign n28779 = n25723 & ~n28728;
  assign n28780 = P1_P3_INSTADDRPOINTER_REG_8_ & n28691;
  assign n28781 = ~P1_P3_INSTADDRPOINTER_REG_9_ & n28780;
  assign n28782 = P1_P3_INSTADDRPOINTER_REG_9_ & ~n28780;
  assign n28783 = ~n28781 & ~n28782;
  assign n28784 = n25739 & ~n28783;
  assign n28785 = n25731 & ~n28783;
  assign n28786 = ~n28777 & ~n28778;
  assign n28787 = ~n28779 & n28786;
  assign n28788 = ~n28784 & n28787;
  assign n28789 = ~n28785 & n28788;
  assign n28790 = P1_P3_INSTADDRPOINTER_REG_8_ & n28706;
  assign n28791 = ~P1_P3_INSTADDRPOINTER_REG_8_ & ~n28706;
  assign n28792 = ~n28705 & ~n28791;
  assign n28793 = ~n28790 & ~n28792;
  assign n28794 = ~P1_P3_INSTADDRPOINTER_REG_9_ & n28793;
  assign n28795 = P1_P3_INSTADDRPOINTER_REG_9_ & ~n28793;
  assign n28796 = ~n28794 & ~n28795;
  assign n28797 = n25742 & n28796;
  assign n28798 = n28776 & n28789;
  assign n28799 = ~n28797 & n28798;
  assign n28800 = n28741 & ~n28742;
  assign n28801 = ~n28757 & n28800;
  assign n28802 = n28769 & n28801;
  assign n28803 = n28799 & n28802;
  assign n28804 = n27634 & ~n28803;
  assign n28805 = ~n28723 & ~n28724;
  assign n4351 = n28804 | ~n28805;
  assign n28807 = P1_P3_INSTADDRPOINTER_REG_10_ & n27633;
  assign n28808 = P1_P3_REIP_REG_10_ & n27778;
  assign n28809 = P1_P3_INSTADDRPOINTER_REG_9_ & n28731;
  assign n28810 = ~P1_P3_INSTADDRPOINTER_REG_10_ & n28809;
  assign n28811 = P1_P3_INSTADDRPOINTER_REG_10_ & ~n28809;
  assign n28812 = ~n28810 & ~n28811;
  assign n28813 = ~n25828 & ~n28812;
  assign n28814 = P1_P3_INSTADDRPOINTER_REG_9_ & n28725;
  assign n28815 = ~P1_P3_INSTADDRPOINTER_REG_10_ & n28814;
  assign n28816 = P1_P3_INSTADDRPOINTER_REG_10_ & ~n28814;
  assign n28817 = ~n28815 & ~n28816;
  assign n28818 = n25899 & ~n28817;
  assign n28819 = n25900 & ~n28817;
  assign n28820 = n27642 & ~n28812;
  assign n28821 = n25715 & ~n28817;
  assign n28822 = n27645 & ~n28812;
  assign n28823 = ~n28821 & ~n28822;
  assign n28824 = ~n28818 & ~n28819;
  assign n28825 = ~n28820 & n28824;
  assign n28826 = n28823 & n28825;
  assign n28827 = ~P1_P3_INSTADDRPOINTER_REG_10_ & ~n28766;
  assign n28828 = P1_P3_INSTADDRPOINTER_REG_9_ & P1_P3_INSTADDRPOINTER_REG_10_;
  assign n28829 = ~n28764 & n28828;
  assign n28830 = ~n28827 & ~n28829;
  assign n28831 = n27741 & n28830;
  assign n28832 = n27758 & ~n28812;
  assign n28833 = n25785 & ~n28812;
  assign n28834 = n27747 & ~n28812;
  assign n28835 = n27751 & ~n28812;
  assign n28836 = ~n28832 & ~n28833;
  assign n28837 = ~n28834 & n28836;
  assign n28838 = ~n28835 & n28837;
  assign n28839 = n25641 & ~n28817;
  assign n28840 = n25719 & ~n28817;
  assign n28841 = n25723 & ~n28817;
  assign n28842 = P1_P3_INSTADDRPOINTER_REG_9_ & n28780;
  assign n28843 = ~P1_P3_INSTADDRPOINTER_REG_10_ & n28842;
  assign n28844 = P1_P3_INSTADDRPOINTER_REG_10_ & ~n28842;
  assign n28845 = ~n28843 & ~n28844;
  assign n28846 = n25739 & ~n28845;
  assign n28847 = n25731 & ~n28845;
  assign n28848 = ~n28839 & ~n28840;
  assign n28849 = ~n28841 & n28848;
  assign n28850 = ~n28846 & n28849;
  assign n28851 = ~n28847 & n28850;
  assign n28852 = ~P1_P3_INSTADDRPOINTER_REG_10_ & ~n28795;
  assign n28853 = ~n28793 & n28828;
  assign n28854 = ~n28852 & ~n28853;
  assign n28855 = n25742 & n28854;
  assign n28856 = n28838 & n28851;
  assign n28857 = ~n28855 & n28856;
  assign n28858 = n25938 & ~n28812;
  assign n28859 = n25781 & ~n28812;
  assign n28860 = ~n28858 & ~n28859;
  assign n28861 = ~n28747 & ~n28753;
  assign n28862 = ~n28752 & ~n28861;
  assign n28863 = ~P1_P3_INSTADDRPOINTER_REG_10_ & ~n28561;
  assign n28864 = P1_P3_INSTADDRPOINTER_REG_10_ & n28561;
  assign n28865 = ~n28863 & ~n28864;
  assign n28866 = n28862 & ~n28865;
  assign n28867 = P1_P3_INSTADDRPOINTER_REG_10_ & ~n28561;
  assign n28868 = ~P1_P3_INSTADDRPOINTER_REG_10_ & n28561;
  assign n28869 = ~n28867 & ~n28868;
  assign n28870 = ~n28862 & ~n28869;
  assign n28871 = ~n28866 & ~n28870;
  assign n28872 = n27739 & ~n28871;
  assign n28873 = n28860 & ~n28872;
  assign n28874 = ~n28813 & n28826;
  assign n28875 = ~n28831 & n28874;
  assign n28876 = n28857 & n28875;
  assign n28877 = n28873 & n28876;
  assign n28878 = n27634 & ~n28877;
  assign n28879 = ~n28807 & ~n28808;
  assign n4356 = n28878 | ~n28879;
  assign n28881 = P1_P3_INSTADDRPOINTER_REG_11_ & n27633;
  assign n28882 = P1_P3_REIP_REG_11_ & n27778;
  assign n28883 = P1_P3_INSTADDRPOINTER_REG_10_ & n28809;
  assign n28884 = ~P1_P3_INSTADDRPOINTER_REG_11_ & n28883;
  assign n28885 = P1_P3_INSTADDRPOINTER_REG_11_ & ~n28883;
  assign n28886 = ~n28884 & ~n28885;
  assign n28887 = ~n25828 & ~n28886;
  assign n28888 = P1_P3_INSTADDRPOINTER_REG_10_ & n28814;
  assign n28889 = ~P1_P3_INSTADDRPOINTER_REG_11_ & n28888;
  assign n28890 = P1_P3_INSTADDRPOINTER_REG_11_ & ~n28888;
  assign n28891 = ~n28889 & ~n28890;
  assign n28892 = n25899 & ~n28891;
  assign n28893 = n25900 & ~n28891;
  assign n28894 = n27642 & ~n28886;
  assign n28895 = n25715 & ~n28891;
  assign n28896 = n27645 & ~n28886;
  assign n28897 = ~n28895 & ~n28896;
  assign n28898 = ~n28892 & ~n28893;
  assign n28899 = ~n28894 & n28898;
  assign n28900 = n28897 & n28899;
  assign n28901 = P1_P3_INSTADDRPOINTER_REG_11_ & ~n28829;
  assign n28902 = ~P1_P3_INSTADDRPOINTER_REG_11_ & n28829;
  assign n28903 = ~n28901 & ~n28902;
  assign n28904 = n27741 & ~n28903;
  assign n28905 = n25938 & ~n28886;
  assign n28906 = n25781 & ~n28886;
  assign n28907 = ~n28905 & ~n28906;
  assign n28908 = ~n28753 & ~n28868;
  assign n28909 = ~n28747 & n28908;
  assign n28910 = ~n28752 & ~n28867;
  assign n28911 = ~n28909 & n28910;
  assign n28912 = ~P1_P3_INSTADDRPOINTER_REG_11_ & ~n28561;
  assign n28913 = P1_P3_INSTADDRPOINTER_REG_11_ & n28561;
  assign n28914 = ~n28912 & ~n28913;
  assign n28915 = n28911 & ~n28914;
  assign n28916 = ~n28911 & n28914;
  assign n28917 = ~n28915 & ~n28916;
  assign n28918 = n27739 & ~n28917;
  assign n28919 = n28907 & ~n28918;
  assign n28920 = n27758 & ~n28886;
  assign n28921 = n25785 & ~n28886;
  assign n28922 = n27747 & ~n28886;
  assign n28923 = n27751 & ~n28886;
  assign n28924 = ~n28920 & ~n28921;
  assign n28925 = ~n28922 & n28924;
  assign n28926 = ~n28923 & n28925;
  assign n28927 = n25641 & ~n28891;
  assign n28928 = n25719 & ~n28891;
  assign n28929 = n25723 & ~n28891;
  assign n28930 = P1_P3_INSTADDRPOINTER_REG_10_ & n28842;
  assign n28931 = ~P1_P3_INSTADDRPOINTER_REG_11_ & n28930;
  assign n28932 = P1_P3_INSTADDRPOINTER_REG_11_ & ~n28930;
  assign n28933 = ~n28931 & ~n28932;
  assign n28934 = n25739 & ~n28933;
  assign n28935 = n25731 & ~n28933;
  assign n28936 = ~n28927 & ~n28928;
  assign n28937 = ~n28929 & n28936;
  assign n28938 = ~n28934 & n28937;
  assign n28939 = ~n28935 & n28938;
  assign n28940 = P1_P3_INSTADDRPOINTER_REG_11_ & ~n28853;
  assign n28941 = ~P1_P3_INSTADDRPOINTER_REG_11_ & n28853;
  assign n28942 = ~n28940 & ~n28941;
  assign n28943 = n25742 & ~n28942;
  assign n28944 = n28926 & n28939;
  assign n28945 = ~n28943 & n28944;
  assign n28946 = ~n28887 & n28900;
  assign n28947 = ~n28904 & n28946;
  assign n28948 = n28919 & n28947;
  assign n28949 = n28945 & n28948;
  assign n28950 = n27634 & ~n28949;
  assign n28951 = ~n28881 & ~n28882;
  assign n4361 = n28950 | ~n28951;
  assign n28953 = P1_P3_INSTADDRPOINTER_REG_12_ & n27633;
  assign n28954 = P1_P3_REIP_REG_12_ & n27778;
  assign n28955 = P1_P3_INSTADDRPOINTER_REG_11_ & n28888;
  assign n28956 = ~P1_P3_INSTADDRPOINTER_REG_12_ & n28955;
  assign n28957 = P1_P3_INSTADDRPOINTER_REG_12_ & ~n28955;
  assign n28958 = ~n28956 & ~n28957;
  assign n28959 = n25899 & ~n28958;
  assign n28960 = n25900 & ~n28958;
  assign n28961 = P1_P3_INSTADDRPOINTER_REG_11_ & n28883;
  assign n28962 = ~P1_P3_INSTADDRPOINTER_REG_12_ & n28961;
  assign n28963 = P1_P3_INSTADDRPOINTER_REG_12_ & ~n28961;
  assign n28964 = ~n28962 & ~n28963;
  assign n28965 = n27642 & ~n28964;
  assign n28966 = n25715 & ~n28958;
  assign n28967 = n27645 & ~n28964;
  assign n28968 = ~n28966 & ~n28967;
  assign n28969 = ~n28959 & ~n28960;
  assign n28970 = ~n28965 & n28969;
  assign n28971 = n28968 & n28970;
  assign n28972 = ~n25828 & ~n28964;
  assign n28973 = ~P1_P3_INSTADDRPOINTER_REG_12_ & ~n28561;
  assign n28974 = P1_P3_INSTADDRPOINTER_REG_12_ & n28561;
  assign n28975 = ~n28973 & ~n28974;
  assign n28976 = ~P1_P3_INSTADDRPOINTER_REG_11_ & n28561;
  assign n28977 = n28908 & ~n28976;
  assign n28978 = ~n28747 & n28977;
  assign n28979 = P1_P3_INSTADDRPOINTER_REG_11_ & ~n28561;
  assign n28980 = n28910 & ~n28979;
  assign n28981 = ~n28978 & n28980;
  assign n28982 = ~n28975 & n28981;
  assign n28983 = ~P1_P3_INSTADDRPOINTER_REG_12_ & n28561;
  assign n28984 = P1_P3_INSTADDRPOINTER_REG_12_ & ~n28561;
  assign n28985 = ~n28983 & ~n28984;
  assign n28986 = ~n28981 & ~n28985;
  assign n28987 = ~n28982 & ~n28986;
  assign n28988 = n27739 & ~n28987;
  assign n28989 = n25938 & ~n28964;
  assign n28990 = n25781 & ~n28964;
  assign n28991 = ~n28989 & ~n28990;
  assign n28992 = P1_P3_INSTADDRPOINTER_REG_11_ & n28829;
  assign n28993 = ~P1_P3_INSTADDRPOINTER_REG_12_ & ~n28992;
  assign n28994 = P1_P3_INSTADDRPOINTER_REG_11_ & P1_P3_INSTADDRPOINTER_REG_12_;
  assign n28995 = n28829 & n28994;
  assign n28996 = ~n28993 & ~n28995;
  assign n28997 = n27741 & n28996;
  assign n28998 = n28991 & ~n28997;
  assign n28999 = n27758 & ~n28964;
  assign n29000 = n25785 & ~n28964;
  assign n29001 = n27747 & ~n28964;
  assign n29002 = n27751 & ~n28964;
  assign n29003 = ~n28999 & ~n29000;
  assign n29004 = ~n29001 & n29003;
  assign n29005 = ~n29002 & n29004;
  assign n29006 = n25641 & ~n28958;
  assign n29007 = n25719 & ~n28958;
  assign n29008 = n25723 & ~n28958;
  assign n29009 = P1_P3_INSTADDRPOINTER_REG_11_ & n28930;
  assign n29010 = ~P1_P3_INSTADDRPOINTER_REG_12_ & n29009;
  assign n29011 = P1_P3_INSTADDRPOINTER_REG_12_ & ~n29009;
  assign n29012 = ~n29010 & ~n29011;
  assign n29013 = n25739 & ~n29012;
  assign n29014 = n25731 & ~n29012;
  assign n29015 = ~n29006 & ~n29007;
  assign n29016 = ~n29008 & n29015;
  assign n29017 = ~n29013 & n29016;
  assign n29018 = ~n29014 & n29017;
  assign n29019 = P1_P3_INSTADDRPOINTER_REG_11_ & n28853;
  assign n29020 = ~P1_P3_INSTADDRPOINTER_REG_12_ & ~n29019;
  assign n29021 = n28853 & n28994;
  assign n29022 = ~n29020 & ~n29021;
  assign n29023 = n25742 & n29022;
  assign n29024 = n29005 & n29018;
  assign n29025 = ~n29023 & n29024;
  assign n29026 = n28971 & ~n28972;
  assign n29027 = ~n28988 & n29026;
  assign n29028 = n28998 & n29027;
  assign n29029 = n29025 & n29028;
  assign n29030 = n27634 & ~n29029;
  assign n29031 = ~n28953 & ~n28954;
  assign n4366 = n29030 | ~n29031;
  assign n29033 = P1_P3_INSTADDRPOINTER_REG_13_ & n27633;
  assign n29034 = P1_P3_REIP_REG_13_ & n27778;
  assign n29035 = P1_P3_INSTADDRPOINTER_REG_12_ & n28955;
  assign n29036 = ~P1_P3_INSTADDRPOINTER_REG_13_ & n29035;
  assign n29037 = P1_P3_INSTADDRPOINTER_REG_13_ & ~n29035;
  assign n29038 = ~n29036 & ~n29037;
  assign n29039 = n25899 & ~n29038;
  assign n29040 = n25900 & ~n29038;
  assign n29041 = P1_P3_INSTADDRPOINTER_REG_12_ & n28961;
  assign n29042 = ~P1_P3_INSTADDRPOINTER_REG_13_ & n29041;
  assign n29043 = P1_P3_INSTADDRPOINTER_REG_13_ & ~n29041;
  assign n29044 = ~n29042 & ~n29043;
  assign n29045 = n27642 & ~n29044;
  assign n29046 = n25715 & ~n29038;
  assign n29047 = n27645 & ~n29044;
  assign n29048 = ~n29046 & ~n29047;
  assign n29049 = ~n29039 & ~n29040;
  assign n29050 = ~n29045 & n29049;
  assign n29051 = n29048 & n29050;
  assign n29052 = ~n25828 & ~n29044;
  assign n29053 = P1_P3_INSTADDRPOINTER_REG_13_ & ~n28561;
  assign n29054 = P1_P3_INSTADDRPOINTER_REG_12_ & P1_P3_INSTADDRPOINTER_REG_13_;
  assign n29055 = n28561 & ~n29054;
  assign n29056 = ~n29053 & ~n29055;
  assign n29057 = n28981 & ~n28984;
  assign n29058 = n29056 & ~n29057;
  assign n29059 = ~P1_P3_INSTADDRPOINTER_REG_13_ & ~n28561;
  assign n29060 = P1_P3_INSTADDRPOINTER_REG_13_ & n28561;
  assign n29061 = ~n29059 & ~n29060;
  assign n29062 = ~n28984 & n29061;
  assign n29063 = ~n28981 & ~n28983;
  assign n29064 = n29062 & ~n29063;
  assign n29065 = ~n29058 & ~n29064;
  assign n29066 = n27739 & n29065;
  assign n29067 = n25938 & ~n29044;
  assign n29068 = n25781 & ~n29044;
  assign n29069 = ~n29067 & ~n29068;
  assign n29070 = ~P1_P3_INSTADDRPOINTER_REG_13_ & ~n28995;
  assign n29071 = P1_P3_INSTADDRPOINTER_REG_13_ & n28995;
  assign n29072 = ~n29070 & ~n29071;
  assign n29073 = n27741 & n29072;
  assign n29074 = n29069 & ~n29073;
  assign n29075 = n27758 & ~n29044;
  assign n29076 = n25785 & ~n29044;
  assign n29077 = n27747 & ~n29044;
  assign n29078 = n27751 & ~n29044;
  assign n29079 = ~n29075 & ~n29076;
  assign n29080 = ~n29077 & n29079;
  assign n29081 = ~n29078 & n29080;
  assign n29082 = n25641 & ~n29038;
  assign n29083 = n25719 & ~n29038;
  assign n29084 = n25723 & ~n29038;
  assign n29085 = P1_P3_INSTADDRPOINTER_REG_12_ & n29009;
  assign n29086 = ~P1_P3_INSTADDRPOINTER_REG_13_ & n29085;
  assign n29087 = P1_P3_INSTADDRPOINTER_REG_13_ & ~n29085;
  assign n29088 = ~n29086 & ~n29087;
  assign n29089 = n25739 & ~n29088;
  assign n29090 = n25731 & ~n29088;
  assign n29091 = ~n29082 & ~n29083;
  assign n29092 = ~n29084 & n29091;
  assign n29093 = ~n29089 & n29092;
  assign n29094 = ~n29090 & n29093;
  assign n29095 = ~P1_P3_INSTADDRPOINTER_REG_13_ & ~n29021;
  assign n29096 = P1_P3_INSTADDRPOINTER_REG_13_ & n29021;
  assign n29097 = ~n29095 & ~n29096;
  assign n29098 = n25742 & n29097;
  assign n29099 = n29081 & n29094;
  assign n29100 = ~n29098 & n29099;
  assign n29101 = n29051 & ~n29052;
  assign n29102 = ~n29066 & n29101;
  assign n29103 = n29074 & n29102;
  assign n29104 = n29100 & n29103;
  assign n29105 = n27634 & ~n29104;
  assign n29106 = ~n29033 & ~n29034;
  assign n4371 = n29105 | ~n29106;
  assign n29108 = P1_P3_INSTADDRPOINTER_REG_14_ & n27633;
  assign n29109 = P1_P3_REIP_REG_14_ & n27778;
  assign n29110 = ~n29108 & ~n29109;
  assign n29111 = P1_P3_INSTADDRPOINTER_REG_13_ & n29041;
  assign n29112 = ~P1_P3_INSTADDRPOINTER_REG_14_ & n29111;
  assign n29113 = P1_P3_INSTADDRPOINTER_REG_14_ & ~n29111;
  assign n29114 = ~n29112 & ~n29113;
  assign n29115 = n27758 & ~n29114;
  assign n29116 = n25785 & ~n29114;
  assign n29117 = n27747 & ~n29114;
  assign n29118 = n27751 & ~n29114;
  assign n29119 = ~n29115 & ~n29116;
  assign n29120 = ~n29117 & n29119;
  assign n29121 = ~n29118 & n29120;
  assign n29122 = P1_P3_INSTADDRPOINTER_REG_13_ & n29035;
  assign n29123 = ~P1_P3_INSTADDRPOINTER_REG_14_ & n29122;
  assign n29124 = P1_P3_INSTADDRPOINTER_REG_14_ & ~n29122;
  assign n29125 = ~n29123 & ~n29124;
  assign n29126 = n25641 & ~n29125;
  assign n29127 = n25719 & ~n29125;
  assign n29128 = n25723 & ~n29125;
  assign n29129 = P1_P3_INSTADDRPOINTER_REG_13_ & n29085;
  assign n29130 = ~P1_P3_INSTADDRPOINTER_REG_14_ & n29129;
  assign n29131 = P1_P3_INSTADDRPOINTER_REG_14_ & ~n29129;
  assign n29132 = ~n29130 & ~n29131;
  assign n29133 = n25739 & ~n29132;
  assign n29134 = n25731 & ~n29132;
  assign n29135 = ~n29126 & ~n29127;
  assign n29136 = ~n29128 & n29135;
  assign n29137 = ~n29133 & n29136;
  assign n29138 = ~n29134 & n29137;
  assign n29139 = ~P1_P3_INSTADDRPOINTER_REG_14_ & n29096;
  assign n29140 = P1_P3_INSTADDRPOINTER_REG_14_ & ~n29096;
  assign n29141 = ~n29139 & ~n29140;
  assign n29142 = n25742 & ~n29141;
  assign n29143 = n29121 & n29138;
  assign n29144 = ~n29142 & n29143;
  assign n29145 = n25938 & ~n29114;
  assign n29146 = n25781 & ~n29114;
  assign n29147 = ~n29145 & ~n29146;
  assign n29148 = ~n25828 & ~n29114;
  assign n29149 = n25899 & ~n29125;
  assign n29150 = n25900 & ~n29125;
  assign n29151 = n27642 & ~n29114;
  assign n29152 = n25715 & ~n29125;
  assign n29153 = n27645 & ~n29114;
  assign n29154 = ~n29152 & ~n29153;
  assign n29155 = ~n29149 & ~n29150;
  assign n29156 = ~n29151 & n29155;
  assign n29157 = n29154 & n29156;
  assign n29158 = ~n28984 & ~n29053;
  assign n29159 = n28980 & n29158;
  assign n29160 = n28977 & ~n29055;
  assign n29161 = ~n28747 & n29160;
  assign n29162 = n29159 & ~n29161;
  assign n29163 = ~P1_P3_INSTADDRPOINTER_REG_14_ & ~n28561;
  assign n29164 = P1_P3_INSTADDRPOINTER_REG_14_ & n28561;
  assign n29165 = ~n29163 & ~n29164;
  assign n29166 = n29162 & ~n29165;
  assign n29167 = ~n29162 & n29165;
  assign n29168 = ~n29166 & ~n29167;
  assign n29169 = n27739 & ~n29168;
  assign n29170 = ~P1_P3_INSTADDRPOINTER_REG_14_ & n29071;
  assign n29171 = P1_P3_INSTADDRPOINTER_REG_14_ & ~n29071;
  assign n29172 = ~n29170 & ~n29171;
  assign n29173 = n27741 & ~n29172;
  assign n29174 = n29147 & ~n29148;
  assign n29175 = n29157 & n29174;
  assign n29176 = ~n29169 & n29175;
  assign n29177 = ~n29173 & n29176;
  assign n29178 = n29144 & n29177;
  assign n29179 = n27634 & ~n29178;
  assign n4376 = ~n29110 | n29179;
  assign n29181 = P1_P3_INSTADDRPOINTER_REG_15_ & n27633;
  assign n29182 = P1_P3_REIP_REG_15_ & n27778;
  assign n29183 = ~n29181 & ~n29182;
  assign n29184 = P1_P3_INSTADDRPOINTER_REG_14_ & n29111;
  assign n29185 = ~P1_P3_INSTADDRPOINTER_REG_15_ & n29184;
  assign n29186 = P1_P3_INSTADDRPOINTER_REG_15_ & ~n29184;
  assign n29187 = ~n29185 & ~n29186;
  assign n29188 = n27758 & ~n29187;
  assign n29189 = n25785 & ~n29187;
  assign n29190 = n27747 & ~n29187;
  assign n29191 = n27751 & ~n29187;
  assign n29192 = ~n29188 & ~n29189;
  assign n29193 = ~n29190 & n29192;
  assign n29194 = ~n29191 & n29193;
  assign n29195 = P1_P3_INSTADDRPOINTER_REG_14_ & n29122;
  assign n29196 = ~P1_P3_INSTADDRPOINTER_REG_15_ & n29195;
  assign n29197 = P1_P3_INSTADDRPOINTER_REG_15_ & ~n29195;
  assign n29198 = ~n29196 & ~n29197;
  assign n29199 = n25641 & ~n29198;
  assign n29200 = n25719 & ~n29198;
  assign n29201 = n25723 & ~n29198;
  assign n29202 = P1_P3_INSTADDRPOINTER_REG_14_ & n29129;
  assign n29203 = ~P1_P3_INSTADDRPOINTER_REG_15_ & n29202;
  assign n29204 = P1_P3_INSTADDRPOINTER_REG_15_ & ~n29202;
  assign n29205 = ~n29203 & ~n29204;
  assign n29206 = n25739 & ~n29205;
  assign n29207 = n25731 & ~n29205;
  assign n29208 = ~n29199 & ~n29200;
  assign n29209 = ~n29201 & n29208;
  assign n29210 = ~n29206 & n29209;
  assign n29211 = ~n29207 & n29210;
  assign n29212 = P1_P3_INSTADDRPOINTER_REG_14_ & n29096;
  assign n29213 = ~P1_P3_INSTADDRPOINTER_REG_15_ & ~n29212;
  assign n29214 = P1_P3_INSTADDRPOINTER_REG_14_ & P1_P3_INSTADDRPOINTER_REG_15_;
  assign n29215 = P1_P3_INSTADDRPOINTER_REG_13_ & n29214;
  assign n29216 = n29021 & n29215;
  assign n29217 = ~n29213 & ~n29216;
  assign n29218 = n25742 & n29217;
  assign n29219 = n29194 & n29211;
  assign n29220 = ~n29218 & n29219;
  assign n29221 = n25938 & ~n29187;
  assign n29222 = n25781 & ~n29187;
  assign n29223 = ~n29221 & ~n29222;
  assign n29224 = ~n25828 & ~n29187;
  assign n29225 = n25899 & ~n29198;
  assign n29226 = n25900 & ~n29198;
  assign n29227 = n27642 & ~n29187;
  assign n29228 = n25715 & ~n29198;
  assign n29229 = n27645 & ~n29187;
  assign n29230 = ~n29228 & ~n29229;
  assign n29231 = ~n29225 & ~n29226;
  assign n29232 = ~n29227 & n29231;
  assign n29233 = n29230 & n29232;
  assign n29234 = P1_P3_INSTADDRPOINTER_REG_14_ & ~n28561;
  assign n29235 = ~P1_P3_INSTADDRPOINTER_REG_14_ & n28561;
  assign n29236 = ~n29162 & ~n29235;
  assign n29237 = ~n29234 & ~n29236;
  assign n29238 = ~P1_P3_INSTADDRPOINTER_REG_15_ & ~n28561;
  assign n29239 = P1_P3_INSTADDRPOINTER_REG_15_ & n28561;
  assign n29240 = ~n29238 & ~n29239;
  assign n29241 = n29237 & ~n29240;
  assign n29242 = ~n29237 & n29240;
  assign n29243 = ~n29241 & ~n29242;
  assign n29244 = n27739 & ~n29243;
  assign n29245 = P1_P3_INSTADDRPOINTER_REG_14_ & n29071;
  assign n29246 = ~P1_P3_INSTADDRPOINTER_REG_15_ & ~n29245;
  assign n29247 = n28995 & n29215;
  assign n29248 = ~n29246 & ~n29247;
  assign n29249 = n27741 & n29248;
  assign n29250 = n29223 & ~n29224;
  assign n29251 = n29233 & n29250;
  assign n29252 = ~n29244 & n29251;
  assign n29253 = ~n29249 & n29252;
  assign n29254 = n29220 & n29253;
  assign n29255 = n27634 & ~n29254;
  assign n4381 = ~n29183 | n29255;
  assign n29257 = P1_P3_INSTADDRPOINTER_REG_16_ & n27633;
  assign n29258 = P1_P3_REIP_REG_16_ & n27778;
  assign n29259 = P1_P3_INSTADDRPOINTER_REG_15_ & n29184;
  assign n29260 = ~P1_P3_INSTADDRPOINTER_REG_16_ & n29259;
  assign n29261 = P1_P3_INSTADDRPOINTER_REG_16_ & ~n29259;
  assign n29262 = ~n29260 & ~n29261;
  assign n29263 = ~n25828 & ~n29262;
  assign n29264 = P1_P3_INSTADDRPOINTER_REG_15_ & n29195;
  assign n29265 = ~P1_P3_INSTADDRPOINTER_REG_16_ & n29264;
  assign n29266 = P1_P3_INSTADDRPOINTER_REG_16_ & ~n29264;
  assign n29267 = ~n29265 & ~n29266;
  assign n29268 = n25899 & ~n29267;
  assign n29269 = n25900 & ~n29267;
  assign n29270 = n27642 & ~n29262;
  assign n29271 = n25715 & ~n29267;
  assign n29272 = n27645 & ~n29262;
  assign n29273 = ~n29271 & ~n29272;
  assign n29274 = ~n29268 & ~n29269;
  assign n29275 = ~n29270 & n29274;
  assign n29276 = n29273 & n29275;
  assign n29277 = ~P1_P3_INSTADDRPOINTER_REG_16_ & n29247;
  assign n29278 = P1_P3_INSTADDRPOINTER_REG_16_ & ~n29247;
  assign n29279 = ~n29277 & ~n29278;
  assign n29280 = n27741 & ~n29279;
  assign n29281 = n25938 & ~n29262;
  assign n29282 = n25781 & ~n29262;
  assign n29283 = ~n29281 & ~n29282;
  assign n29284 = P1_P3_INSTADDRPOINTER_REG_15_ & ~n28561;
  assign n29285 = ~P1_P3_INSTADDRPOINTER_REG_15_ & n28561;
  assign n29286 = ~n29237 & ~n29285;
  assign n29287 = ~n29284 & ~n29286;
  assign n29288 = ~P1_P3_INSTADDRPOINTER_REG_16_ & ~n28561;
  assign n29289 = P1_P3_INSTADDRPOINTER_REG_16_ & n28561;
  assign n29290 = ~n29288 & ~n29289;
  assign n29291 = n29287 & ~n29290;
  assign n29292 = ~n29287 & n29290;
  assign n29293 = ~n29291 & ~n29292;
  assign n29294 = n27739 & ~n29293;
  assign n29295 = n29283 & ~n29294;
  assign n29296 = n27758 & ~n29262;
  assign n29297 = n25785 & ~n29262;
  assign n29298 = n27747 & ~n29262;
  assign n29299 = n27751 & ~n29262;
  assign n29300 = ~n29296 & ~n29297;
  assign n29301 = ~n29298 & n29300;
  assign n29302 = ~n29299 & n29301;
  assign n29303 = n25641 & ~n29267;
  assign n29304 = n25719 & ~n29267;
  assign n29305 = n25723 & ~n29267;
  assign n29306 = P1_P3_INSTADDRPOINTER_REG_15_ & n29202;
  assign n29307 = ~P1_P3_INSTADDRPOINTER_REG_16_ & n29306;
  assign n29308 = P1_P3_INSTADDRPOINTER_REG_16_ & ~n29306;
  assign n29309 = ~n29307 & ~n29308;
  assign n29310 = n25739 & ~n29309;
  assign n29311 = n25731 & ~n29309;
  assign n29312 = ~n29303 & ~n29304;
  assign n29313 = ~n29305 & n29312;
  assign n29314 = ~n29310 & n29313;
  assign n29315 = ~n29311 & n29314;
  assign n29316 = ~P1_P3_INSTADDRPOINTER_REG_16_ & n29216;
  assign n29317 = P1_P3_INSTADDRPOINTER_REG_16_ & ~n29216;
  assign n29318 = ~n29316 & ~n29317;
  assign n29319 = n25742 & ~n29318;
  assign n29320 = n29302 & n29315;
  assign n29321 = ~n29319 & n29320;
  assign n29322 = ~n29263 & n29276;
  assign n29323 = ~n29280 & n29322;
  assign n29324 = n29295 & n29323;
  assign n29325 = n29321 & n29324;
  assign n29326 = n27634 & ~n29325;
  assign n29327 = ~n29257 & ~n29258;
  assign n4386 = n29326 | ~n29327;
  assign n29329 = P1_P3_INSTADDRPOINTER_REG_17_ & n27633;
  assign n29330 = P1_P3_REIP_REG_17_ & n27778;
  assign n29331 = P1_P3_INSTADDRPOINTER_REG_16_ & n29259;
  assign n29332 = ~P1_P3_INSTADDRPOINTER_REG_17_ & n29331;
  assign n29333 = P1_P3_INSTADDRPOINTER_REG_17_ & ~n29331;
  assign n29334 = ~n29332 & ~n29333;
  assign n29335 = ~n25828 & ~n29334;
  assign n29336 = n25938 & ~n29334;
  assign n29337 = n25781 & ~n29334;
  assign n29338 = ~n29336 & ~n29337;
  assign n29339 = P1_P3_INSTADDRPOINTER_REG_16_ & n29247;
  assign n29340 = ~P1_P3_INSTADDRPOINTER_REG_17_ & ~n29339;
  assign n29341 = P1_P3_INSTADDRPOINTER_REG_16_ & P1_P3_INSTADDRPOINTER_REG_17_;
  assign n29342 = n29247 & n29341;
  assign n29343 = ~n29340 & ~n29342;
  assign n29344 = n27741 & n29343;
  assign n29345 = n27758 & ~n29334;
  assign n29346 = n25785 & ~n29334;
  assign n29347 = n27747 & ~n29334;
  assign n29348 = n27751 & ~n29334;
  assign n29349 = ~n29345 & ~n29346;
  assign n29350 = ~n29347 & n29349;
  assign n29351 = ~n29348 & n29350;
  assign n29352 = P1_P3_INSTADDRPOINTER_REG_16_ & n29264;
  assign n29353 = ~P1_P3_INSTADDRPOINTER_REG_17_ & n29352;
  assign n29354 = P1_P3_INSTADDRPOINTER_REG_17_ & ~n29352;
  assign n29355 = ~n29353 & ~n29354;
  assign n29356 = n25641 & ~n29355;
  assign n29357 = n25719 & ~n29355;
  assign n29358 = n25723 & ~n29355;
  assign n29359 = P1_P3_INSTADDRPOINTER_REG_16_ & n29306;
  assign n29360 = ~P1_P3_INSTADDRPOINTER_REG_17_ & n29359;
  assign n29361 = P1_P3_INSTADDRPOINTER_REG_17_ & ~n29359;
  assign n29362 = ~n29360 & ~n29361;
  assign n29363 = n25739 & ~n29362;
  assign n29364 = n25731 & ~n29362;
  assign n29365 = ~n29356 & ~n29357;
  assign n29366 = ~n29358 & n29365;
  assign n29367 = ~n29363 & n29366;
  assign n29368 = ~n29364 & n29367;
  assign n29369 = P1_P3_INSTADDRPOINTER_REG_16_ & n29216;
  assign n29370 = ~P1_P3_INSTADDRPOINTER_REG_17_ & ~n29369;
  assign n29371 = n29216 & n29341;
  assign n29372 = ~n29370 & ~n29371;
  assign n29373 = n25742 & n29372;
  assign n29374 = n29351 & n29368;
  assign n29375 = ~n29373 & n29374;
  assign n29376 = n25899 & ~n29355;
  assign n29377 = n25900 & ~n29355;
  assign n29378 = n27642 & ~n29334;
  assign n29379 = n25715 & ~n29355;
  assign n29380 = n27645 & ~n29334;
  assign n29381 = ~n29379 & ~n29380;
  assign n29382 = ~n29287 & n29341;
  assign n29383 = n28561 & ~n29382;
  assign n29384 = P1_P3_INSTADDRPOINTER_REG_17_ & ~n28561;
  assign n29385 = ~P1_P3_INSTADDRPOINTER_REG_16_ & ~n29284;
  assign n29386 = ~n29286 & n29385;
  assign n29387 = ~n29383 & ~n29384;
  assign n29388 = ~n29386 & n29387;
  assign n29389 = P1_P3_INSTADDRPOINTER_REG_17_ & n29386;
  assign n29390 = ~n28561 & ~n29389;
  assign n29391 = P1_P3_INSTADDRPOINTER_REG_17_ & n28561;
  assign n29392 = P1_P3_INSTADDRPOINTER_REG_16_ & ~n29287;
  assign n29393 = ~n29390 & ~n29391;
  assign n29394 = ~n29392 & n29393;
  assign n29395 = ~n29388 & ~n29394;
  assign n29396 = n27739 & n29395;
  assign n29397 = ~n29376 & ~n29377;
  assign n29398 = ~n29378 & n29397;
  assign n29399 = n29381 & n29398;
  assign n29400 = ~n29396 & n29399;
  assign n29401 = ~n29335 & n29338;
  assign n29402 = ~n29344 & n29401;
  assign n29403 = n29375 & n29402;
  assign n29404 = n29400 & n29403;
  assign n29405 = n27634 & ~n29404;
  assign n29406 = ~n29329 & ~n29330;
  assign n4391 = n29405 | ~n29406;
  assign n29408 = P1_P3_INSTADDRPOINTER_REG_18_ & n27633;
  assign n29409 = P1_P3_REIP_REG_18_ & n27778;
  assign n29410 = P1_P3_INSTADDRPOINTER_REG_17_ & n29331;
  assign n29411 = ~P1_P3_INSTADDRPOINTER_REG_18_ & n29410;
  assign n29412 = P1_P3_INSTADDRPOINTER_REG_18_ & ~n29410;
  assign n29413 = ~n29411 & ~n29412;
  assign n29414 = ~n25828 & ~n29413;
  assign n29415 = P1_P3_INSTADDRPOINTER_REG_17_ & n29352;
  assign n29416 = ~P1_P3_INSTADDRPOINTER_REG_18_ & n29415;
  assign n29417 = P1_P3_INSTADDRPOINTER_REG_18_ & ~n29415;
  assign n29418 = ~n29416 & ~n29417;
  assign n29419 = n25899 & ~n29418;
  assign n29420 = n25900 & ~n29418;
  assign n29421 = n27642 & ~n29413;
  assign n29422 = n25715 & ~n29418;
  assign n29423 = n27645 & ~n29413;
  assign n29424 = ~n29422 & ~n29423;
  assign n29425 = ~n29419 & ~n29420;
  assign n29426 = ~n29421 & n29425;
  assign n29427 = n29424 & n29426;
  assign n29428 = ~P1_P3_INSTADDRPOINTER_REG_18_ & n29342;
  assign n29429 = P1_P3_INSTADDRPOINTER_REG_18_ & ~n29342;
  assign n29430 = ~n29428 & ~n29429;
  assign n29431 = n27741 & ~n29430;
  assign n29432 = n25938 & ~n29413;
  assign n29433 = n25781 & ~n29413;
  assign n29434 = ~n29432 & ~n29433;
  assign n29435 = ~n28561 & ~n29386;
  assign n29436 = ~n29382 & ~n29435;
  assign n29437 = ~n29384 & n29436;
  assign n29438 = ~P1_P3_INSTADDRPOINTER_REG_18_ & ~n28561;
  assign n29439 = P1_P3_INSTADDRPOINTER_REG_18_ & n28561;
  assign n29440 = ~n29438 & ~n29439;
  assign n29441 = n29437 & ~n29440;
  assign n29442 = ~n29437 & n29440;
  assign n29443 = ~n29441 & ~n29442;
  assign n29444 = n27739 & ~n29443;
  assign n29445 = n29434 & ~n29444;
  assign n29446 = n27758 & ~n29413;
  assign n29447 = n25785 & ~n29413;
  assign n29448 = n27747 & ~n29413;
  assign n29449 = n27751 & ~n29413;
  assign n29450 = ~n29446 & ~n29447;
  assign n29451 = ~n29448 & n29450;
  assign n29452 = ~n29449 & n29451;
  assign n29453 = n25641 & ~n29418;
  assign n29454 = n25719 & ~n29418;
  assign n29455 = n25723 & ~n29418;
  assign n29456 = P1_P3_INSTADDRPOINTER_REG_17_ & n29359;
  assign n29457 = ~P1_P3_INSTADDRPOINTER_REG_18_ & n29456;
  assign n29458 = P1_P3_INSTADDRPOINTER_REG_18_ & ~n29456;
  assign n29459 = ~n29457 & ~n29458;
  assign n29460 = n25739 & ~n29459;
  assign n29461 = n25731 & ~n29459;
  assign n29462 = ~n29453 & ~n29454;
  assign n29463 = ~n29455 & n29462;
  assign n29464 = ~n29460 & n29463;
  assign n29465 = ~n29461 & n29464;
  assign n29466 = ~P1_P3_INSTADDRPOINTER_REG_18_ & n29371;
  assign n29467 = P1_P3_INSTADDRPOINTER_REG_18_ & ~n29371;
  assign n29468 = ~n29466 & ~n29467;
  assign n29469 = n25742 & ~n29468;
  assign n29470 = n29452 & n29465;
  assign n29471 = ~n29469 & n29470;
  assign n29472 = ~n29414 & n29427;
  assign n29473 = ~n29431 & n29472;
  assign n29474 = n29445 & n29473;
  assign n29475 = n29471 & n29474;
  assign n29476 = n27634 & ~n29475;
  assign n29477 = ~n29408 & ~n29409;
  assign n4396 = n29476 | ~n29477;
  assign n29479 = P1_P3_INSTADDRPOINTER_REG_19_ & n27633;
  assign n29480 = P1_P3_REIP_REG_19_ & n27778;
  assign n29481 = P1_P3_INSTADDRPOINTER_REG_18_ & n29410;
  assign n29482 = ~P1_P3_INSTADDRPOINTER_REG_19_ & n29481;
  assign n29483 = P1_P3_INSTADDRPOINTER_REG_19_ & ~n29481;
  assign n29484 = ~n29482 & ~n29483;
  assign n29485 = ~n25828 & ~n29484;
  assign n29486 = n25938 & ~n29484;
  assign n29487 = n25781 & ~n29484;
  assign n29488 = ~n29486 & ~n29487;
  assign n29489 = P1_P3_INSTADDRPOINTER_REG_18_ & n29342;
  assign n29490 = ~P1_P3_INSTADDRPOINTER_REG_19_ & ~n29489;
  assign n29491 = P1_P3_INSTADDRPOINTER_REG_18_ & P1_P3_INSTADDRPOINTER_REG_19_;
  assign n29492 = n29342 & n29491;
  assign n29493 = ~n29490 & ~n29492;
  assign n29494 = n27741 & n29493;
  assign n29495 = n27758 & ~n29484;
  assign n29496 = n25785 & ~n29484;
  assign n29497 = n27747 & ~n29484;
  assign n29498 = n27751 & ~n29484;
  assign n29499 = ~n29495 & ~n29496;
  assign n29500 = ~n29497 & n29499;
  assign n29501 = ~n29498 & n29500;
  assign n29502 = P1_P3_INSTADDRPOINTER_REG_18_ & n29415;
  assign n29503 = ~P1_P3_INSTADDRPOINTER_REG_19_ & n29502;
  assign n29504 = P1_P3_INSTADDRPOINTER_REG_19_ & ~n29502;
  assign n29505 = ~n29503 & ~n29504;
  assign n29506 = n25641 & ~n29505;
  assign n29507 = n25719 & ~n29505;
  assign n29508 = n25723 & ~n29505;
  assign n29509 = P1_P3_INSTADDRPOINTER_REG_18_ & n29456;
  assign n29510 = ~P1_P3_INSTADDRPOINTER_REG_19_ & n29509;
  assign n29511 = P1_P3_INSTADDRPOINTER_REG_19_ & ~n29509;
  assign n29512 = ~n29510 & ~n29511;
  assign n29513 = n25739 & ~n29512;
  assign n29514 = n25731 & ~n29512;
  assign n29515 = ~n29506 & ~n29507;
  assign n29516 = ~n29508 & n29515;
  assign n29517 = ~n29513 & n29516;
  assign n29518 = ~n29514 & n29517;
  assign n29519 = P1_P3_INSTADDRPOINTER_REG_18_ & n29371;
  assign n29520 = ~P1_P3_INSTADDRPOINTER_REG_19_ & ~n29519;
  assign n29521 = n29371 & n29491;
  assign n29522 = ~n29520 & ~n29521;
  assign n29523 = n25742 & n29522;
  assign n29524 = n29501 & n29518;
  assign n29525 = ~n29523 & n29524;
  assign n29526 = n25899 & ~n29505;
  assign n29527 = n25900 & ~n29505;
  assign n29528 = n27642 & ~n29484;
  assign n29529 = n25715 & ~n29505;
  assign n29530 = n27645 & ~n29484;
  assign n29531 = ~n29529 & ~n29530;
  assign n29532 = ~P1_P3_INSTADDRPOINTER_REG_19_ & ~n28561;
  assign n29533 = P1_P3_INSTADDRPOINTER_REG_19_ & n28561;
  assign n29534 = ~n29532 & ~n29533;
  assign n29535 = ~P1_P3_INSTADDRPOINTER_REG_18_ & n28561;
  assign n29536 = ~n29437 & ~n29535;
  assign n29537 = P1_P3_INSTADDRPOINTER_REG_18_ & ~n28561;
  assign n29538 = ~n29536 & ~n29537;
  assign n29539 = ~n29534 & n29538;
  assign n29540 = ~P1_P3_INSTADDRPOINTER_REG_19_ & n28561;
  assign n29541 = P1_P3_INSTADDRPOINTER_REG_19_ & ~n28561;
  assign n29542 = ~n29540 & ~n29541;
  assign n29543 = ~n29538 & ~n29542;
  assign n29544 = ~n29539 & ~n29543;
  assign n29545 = n27739 & ~n29544;
  assign n29546 = ~n29526 & ~n29527;
  assign n29547 = ~n29528 & n29546;
  assign n29548 = n29531 & n29547;
  assign n29549 = ~n29545 & n29548;
  assign n29550 = ~n29485 & n29488;
  assign n29551 = ~n29494 & n29550;
  assign n29552 = n29525 & n29551;
  assign n29553 = n29549 & n29552;
  assign n29554 = n27634 & ~n29553;
  assign n29555 = ~n29479 & ~n29480;
  assign n4401 = n29554 | ~n29555;
  assign n29557 = P1_P3_INSTADDRPOINTER_REG_20_ & n27633;
  assign n29558 = P1_P3_REIP_REG_20_ & n27778;
  assign n29559 = ~n29557 & ~n29558;
  assign n29560 = P1_P3_INSTADDRPOINTER_REG_19_ & P1_P3_INSTADDRPOINTER_REG_20_;
  assign n29561 = n28561 & ~n29560;
  assign n29562 = P1_P3_INSTADDRPOINTER_REG_20_ & ~n28561;
  assign n29563 = ~n29561 & ~n29562;
  assign n29564 = n29538 & ~n29541;
  assign n29565 = n29563 & ~n29564;
  assign n29566 = ~P1_P3_INSTADDRPOINTER_REG_19_ & n29538;
  assign n29567 = P1_P3_INSTADDRPOINTER_REG_20_ & n29566;
  assign n29568 = ~n28561 & ~n29567;
  assign n29569 = P1_P3_INSTADDRPOINTER_REG_20_ & n28561;
  assign n29570 = P1_P3_INSTADDRPOINTER_REG_19_ & ~n29538;
  assign n29571 = ~n29568 & ~n29569;
  assign n29572 = ~n29570 & n29571;
  assign n29573 = ~n29565 & ~n29572;
  assign n29574 = n27739 & n29573;
  assign n29575 = P1_P3_INSTADDRPOINTER_REG_19_ & n29481;
  assign n29576 = ~P1_P3_INSTADDRPOINTER_REG_20_ & n29575;
  assign n29577 = P1_P3_INSTADDRPOINTER_REG_20_ & ~n29575;
  assign n29578 = ~n29576 & ~n29577;
  assign n29579 = ~n25828 & ~n29578;
  assign n29580 = n25938 & ~n29578;
  assign n29581 = n25781 & ~n29578;
  assign n29582 = ~n29580 & ~n29581;
  assign n29583 = P1_P3_INSTADDRPOINTER_REG_19_ & n29502;
  assign n29584 = ~P1_P3_INSTADDRPOINTER_REG_20_ & n29583;
  assign n29585 = P1_P3_INSTADDRPOINTER_REG_20_ & ~n29583;
  assign n29586 = ~n29584 & ~n29585;
  assign n29587 = n25899 & ~n29586;
  assign n29588 = n25900 & ~n29586;
  assign n29589 = n27642 & ~n29578;
  assign n29590 = n25715 & ~n29586;
  assign n29591 = n27645 & ~n29578;
  assign n29592 = ~n29590 & ~n29591;
  assign n29593 = ~n29587 & ~n29588;
  assign n29594 = ~n29589 & n29593;
  assign n29595 = n29592 & n29594;
  assign n29596 = ~P1_P3_INSTADDRPOINTER_REG_20_ & ~n29492;
  assign n29597 = P1_P3_INSTADDRPOINTER_REG_20_ & n29492;
  assign n29598 = ~n29596 & ~n29597;
  assign n29599 = n27741 & n29598;
  assign n29600 = n27758 & ~n29578;
  assign n29601 = n25785 & ~n29578;
  assign n29602 = n27747 & ~n29578;
  assign n29603 = n27751 & ~n29578;
  assign n29604 = ~n29600 & ~n29601;
  assign n29605 = ~n29602 & n29604;
  assign n29606 = ~n29603 & n29605;
  assign n29607 = n25641 & ~n29586;
  assign n29608 = n25719 & ~n29586;
  assign n29609 = n25723 & ~n29586;
  assign n29610 = P1_P3_INSTADDRPOINTER_REG_19_ & n29509;
  assign n29611 = ~P1_P3_INSTADDRPOINTER_REG_20_ & n29610;
  assign n29612 = P1_P3_INSTADDRPOINTER_REG_20_ & ~n29610;
  assign n29613 = ~n29611 & ~n29612;
  assign n29614 = n25739 & ~n29613;
  assign n29615 = n25731 & ~n29613;
  assign n29616 = ~n29607 & ~n29608;
  assign n29617 = ~n29609 & n29616;
  assign n29618 = ~n29614 & n29617;
  assign n29619 = ~n29615 & n29618;
  assign n29620 = ~P1_P3_INSTADDRPOINTER_REG_20_ & ~n29521;
  assign n29621 = P1_P3_INSTADDRPOINTER_REG_20_ & n29521;
  assign n29622 = ~n29620 & ~n29621;
  assign n29623 = n25742 & n29622;
  assign n29624 = n29606 & n29619;
  assign n29625 = ~n29623 & n29624;
  assign n29626 = ~n29579 & n29582;
  assign n29627 = n29595 & n29626;
  assign n29628 = ~n29599 & n29627;
  assign n29629 = n29625 & n29628;
  assign n29630 = ~n29574 & n29629;
  assign n29631 = n27634 & ~n29630;
  assign n4406 = ~n29559 | n29631;
  assign n29633 = P1_P3_INSTADDRPOINTER_REG_21_ & n27633;
  assign n29634 = P1_P3_REIP_REG_21_ & n27778;
  assign n29635 = ~n29633 & ~n29634;
  assign n29636 = ~n29538 & n29560;
  assign n29637 = ~n29562 & ~n29636;
  assign n29638 = ~n28561 & ~n29566;
  assign n29639 = n29637 & ~n29638;
  assign n29640 = ~P1_P3_INSTADDRPOINTER_REG_21_ & ~n28561;
  assign n29641 = P1_P3_INSTADDRPOINTER_REG_21_ & n28561;
  assign n29642 = ~n29640 & ~n29641;
  assign n29643 = n29639 & ~n29642;
  assign n29644 = ~n29639 & n29642;
  assign n29645 = ~n29643 & ~n29644;
  assign n29646 = n27739 & ~n29645;
  assign n29647 = P1_P3_INSTADDRPOINTER_REG_20_ & n29575;
  assign n29648 = ~P1_P3_INSTADDRPOINTER_REG_21_ & n29647;
  assign n29649 = P1_P3_INSTADDRPOINTER_REG_21_ & ~n29647;
  assign n29650 = ~n29648 & ~n29649;
  assign n29651 = ~n25828 & ~n29650;
  assign n29652 = n25938 & ~n29650;
  assign n29653 = n25781 & ~n29650;
  assign n29654 = ~n29652 & ~n29653;
  assign n29655 = P1_P3_INSTADDRPOINTER_REG_20_ & n29583;
  assign n29656 = ~P1_P3_INSTADDRPOINTER_REG_21_ & n29655;
  assign n29657 = P1_P3_INSTADDRPOINTER_REG_21_ & ~n29655;
  assign n29658 = ~n29656 & ~n29657;
  assign n29659 = n25899 & ~n29658;
  assign n29660 = n25900 & ~n29658;
  assign n29661 = n27642 & ~n29650;
  assign n29662 = n25715 & ~n29658;
  assign n29663 = n27645 & ~n29650;
  assign n29664 = ~n29662 & ~n29663;
  assign n29665 = ~n29659 & ~n29660;
  assign n29666 = ~n29661 & n29665;
  assign n29667 = n29664 & n29666;
  assign n29668 = ~P1_P3_INSTADDRPOINTER_REG_21_ & ~n29597;
  assign n29669 = P1_P3_INSTADDRPOINTER_REG_21_ & n29597;
  assign n29670 = ~n29668 & ~n29669;
  assign n29671 = n27741 & n29670;
  assign n29672 = n25641 & ~n29658;
  assign n29673 = n25719 & ~n29658;
  assign n29674 = n25723 & ~n29658;
  assign n29675 = P1_P3_INSTADDRPOINTER_REG_20_ & n29610;
  assign n29676 = ~P1_P3_INSTADDRPOINTER_REG_21_ & n29675;
  assign n29677 = P1_P3_INSTADDRPOINTER_REG_21_ & ~n29675;
  assign n29678 = ~n29676 & ~n29677;
  assign n29679 = n25739 & ~n29678;
  assign n29680 = n25731 & ~n29678;
  assign n29681 = ~n29672 & ~n29673;
  assign n29682 = ~n29674 & n29681;
  assign n29683 = ~n29679 & n29682;
  assign n29684 = ~n29680 & n29683;
  assign n29685 = n27758 & ~n29650;
  assign n29686 = n25785 & ~n29650;
  assign n29687 = n27747 & ~n29650;
  assign n29688 = n27751 & ~n29650;
  assign n29689 = ~n29685 & ~n29686;
  assign n29690 = ~n29687 & n29689;
  assign n29691 = ~n29688 & n29690;
  assign n29692 = ~P1_P3_INSTADDRPOINTER_REG_21_ & ~n29621;
  assign n29693 = P1_P3_INSTADDRPOINTER_REG_20_ & P1_P3_INSTADDRPOINTER_REG_21_;
  assign n29694 = n29521 & n29693;
  assign n29695 = ~n29692 & ~n29694;
  assign n29696 = n25742 & n29695;
  assign n29697 = n29684 & n29691;
  assign n29698 = ~n29696 & n29697;
  assign n29699 = ~n29651 & n29654;
  assign n29700 = n29667 & n29699;
  assign n29701 = ~n29671 & n29700;
  assign n29702 = n29698 & n29701;
  assign n29703 = ~n29646 & n29702;
  assign n29704 = n27634 & ~n29703;
  assign n4411 = ~n29635 | n29704;
  assign n29706 = P1_P3_INSTADDRPOINTER_REG_22_ & n27633;
  assign n29707 = P1_P3_REIP_REG_22_ & n27778;
  assign n29708 = ~n29706 & ~n29707;
  assign n29709 = P1_P3_INSTADDRPOINTER_REG_21_ & n29675;
  assign n29710 = ~P1_P3_INSTADDRPOINTER_REG_22_ & n29709;
  assign n29711 = P1_P3_INSTADDRPOINTER_REG_22_ & ~n29709;
  assign n29712 = ~n29710 & ~n29711;
  assign n29713 = n25739 & ~n29712;
  assign n29714 = n25731 & ~n29712;
  assign n29715 = ~n29713 & ~n29714;
  assign n29716 = P1_P3_INSTADDRPOINTER_REG_21_ & n29655;
  assign n29717 = ~P1_P3_INSTADDRPOINTER_REG_22_ & n29716;
  assign n29718 = P1_P3_INSTADDRPOINTER_REG_22_ & ~n29716;
  assign n29719 = ~n29717 & ~n29718;
  assign n29720 = n25641 & ~n29719;
  assign n29721 = n25719 & ~n29719;
  assign n29722 = n25723 & ~n29719;
  assign n29723 = ~n29720 & ~n29721;
  assign n29724 = ~n29722 & n29723;
  assign n29725 = P1_P3_INSTADDRPOINTER_REG_21_ & n29647;
  assign n29726 = ~P1_P3_INSTADDRPOINTER_REG_22_ & n29725;
  assign n29727 = P1_P3_INSTADDRPOINTER_REG_22_ & ~n29725;
  assign n29728 = ~n29726 & ~n29727;
  assign n29729 = n27747 & ~n29728;
  assign n29730 = n27751 & ~n29728;
  assign n29731 = n25785 & ~n29728;
  assign n29732 = ~n29729 & ~n29730;
  assign n29733 = ~n29731 & n29732;
  assign n29734 = ~P1_P3_INSTADDRPOINTER_REG_22_ & n29694;
  assign n29735 = P1_P3_INSTADDRPOINTER_REG_22_ & ~n29694;
  assign n29736 = ~n29734 & ~n29735;
  assign n29737 = n25742 & ~n29736;
  assign n29738 = n27758 & ~n29728;
  assign n29739 = ~n29737 & ~n29738;
  assign n29740 = n29715 & n29724;
  assign n29741 = n29733 & n29740;
  assign n29742 = n29739 & n29741;
  assign n29743 = P1_P3_INSTADDRPOINTER_REG_21_ & n29560;
  assign n29744 = n28561 & ~n29743;
  assign n29745 = ~n29535 & ~n29744;
  assign n29746 = ~n29437 & n29745;
  assign n29747 = P1_P3_INSTADDRPOINTER_REG_21_ & ~n28561;
  assign n29748 = ~n29537 & ~n29747;
  assign n29749 = ~n29541 & n29748;
  assign n29750 = ~n29562 & n29749;
  assign n29751 = ~n29746 & n29750;
  assign n29752 = ~P1_P3_INSTADDRPOINTER_REG_22_ & ~n28561;
  assign n29753 = P1_P3_INSTADDRPOINTER_REG_22_ & n28561;
  assign n29754 = ~n29752 & ~n29753;
  assign n29755 = n29751 & ~n29754;
  assign n29756 = ~n29751 & n29754;
  assign n29757 = ~n29755 & ~n29756;
  assign n29758 = n27739 & ~n29757;
  assign n29759 = ~n25828 & ~n29728;
  assign n29760 = n25938 & ~n29728;
  assign n29761 = n25781 & ~n29728;
  assign n29762 = ~n29760 & ~n29761;
  assign n29763 = n25899 & ~n29719;
  assign n29764 = n25900 & ~n29719;
  assign n29765 = n27642 & ~n29728;
  assign n29766 = n25715 & ~n29719;
  assign n29767 = n27645 & ~n29728;
  assign n29768 = ~n29766 & ~n29767;
  assign n29769 = ~n29763 & ~n29764;
  assign n29770 = ~n29765 & n29769;
  assign n29771 = n29768 & n29770;
  assign n29772 = ~P1_P3_INSTADDRPOINTER_REG_22_ & n29669;
  assign n29773 = P1_P3_INSTADDRPOINTER_REG_22_ & ~n29669;
  assign n29774 = ~n29772 & ~n29773;
  assign n29775 = n27741 & ~n29774;
  assign n29776 = ~n29758 & ~n29759;
  assign n29777 = n29762 & n29776;
  assign n29778 = n29771 & n29777;
  assign n29779 = ~n29775 & n29778;
  assign n29780 = n29742 & n29779;
  assign n29781 = n27634 & ~n29780;
  assign n4416 = ~n29708 | n29781;
  assign n29783 = P1_P3_INSTADDRPOINTER_REG_23_ & n27633;
  assign n29784 = P1_P3_REIP_REG_23_ & n27778;
  assign n29785 = ~n29783 & ~n29784;
  assign n29786 = P1_P3_INSTADDRPOINTER_REG_22_ & n29709;
  assign n29787 = ~P1_P3_INSTADDRPOINTER_REG_23_ & n29786;
  assign n29788 = P1_P3_INSTADDRPOINTER_REG_23_ & ~n29786;
  assign n29789 = ~n29787 & ~n29788;
  assign n29790 = n25739 & ~n29789;
  assign n29791 = n25731 & ~n29789;
  assign n29792 = ~n29790 & ~n29791;
  assign n29793 = P1_P3_INSTADDRPOINTER_REG_22_ & n29716;
  assign n29794 = ~P1_P3_INSTADDRPOINTER_REG_23_ & n29793;
  assign n29795 = P1_P3_INSTADDRPOINTER_REG_23_ & ~n29793;
  assign n29796 = ~n29794 & ~n29795;
  assign n29797 = n25641 & ~n29796;
  assign n29798 = n25719 & ~n29796;
  assign n29799 = n25723 & ~n29796;
  assign n29800 = ~n29797 & ~n29798;
  assign n29801 = ~n29799 & n29800;
  assign n29802 = P1_P3_INSTADDRPOINTER_REG_22_ & n29725;
  assign n29803 = ~P1_P3_INSTADDRPOINTER_REG_23_ & n29802;
  assign n29804 = P1_P3_INSTADDRPOINTER_REG_23_ & ~n29802;
  assign n29805 = ~n29803 & ~n29804;
  assign n29806 = n27747 & ~n29805;
  assign n29807 = n27751 & ~n29805;
  assign n29808 = n25785 & ~n29805;
  assign n29809 = ~n29806 & ~n29807;
  assign n29810 = ~n29808 & n29809;
  assign n29811 = P1_P3_INSTADDRPOINTER_REG_22_ & n29694;
  assign n29812 = ~P1_P3_INSTADDRPOINTER_REG_23_ & ~n29811;
  assign n29813 = P1_P3_INSTADDRPOINTER_REG_22_ & P1_P3_INSTADDRPOINTER_REG_23_;
  assign n29814 = n29694 & n29813;
  assign n29815 = ~n29812 & ~n29814;
  assign n29816 = n25742 & n29815;
  assign n29817 = n27758 & ~n29805;
  assign n29818 = ~n29816 & ~n29817;
  assign n29819 = n29792 & n29801;
  assign n29820 = n29810 & n29819;
  assign n29821 = n29818 & n29820;
  assign n29822 = ~P1_P3_INSTADDRPOINTER_REG_22_ & n28561;
  assign n29823 = n29745 & ~n29822;
  assign n29824 = ~n29437 & n29823;
  assign n29825 = P1_P3_INSTADDRPOINTER_REG_22_ & ~n28561;
  assign n29826 = n29750 & ~n29825;
  assign n29827 = ~n29824 & n29826;
  assign n29828 = ~P1_P3_INSTADDRPOINTER_REG_23_ & ~n28561;
  assign n29829 = P1_P3_INSTADDRPOINTER_REG_23_ & n28561;
  assign n29830 = ~n29828 & ~n29829;
  assign n29831 = n29827 & ~n29830;
  assign n29832 = ~n29827 & n29830;
  assign n29833 = ~n29831 & ~n29832;
  assign n29834 = n27739 & ~n29833;
  assign n29835 = ~n25828 & ~n29805;
  assign n29836 = n25938 & ~n29805;
  assign n29837 = n25781 & ~n29805;
  assign n29838 = ~n29836 & ~n29837;
  assign n29839 = n25899 & ~n29796;
  assign n29840 = n25900 & ~n29796;
  assign n29841 = n27642 & ~n29805;
  assign n29842 = n25715 & ~n29796;
  assign n29843 = n27645 & ~n29805;
  assign n29844 = ~n29842 & ~n29843;
  assign n29845 = ~n29839 & ~n29840;
  assign n29846 = ~n29841 & n29845;
  assign n29847 = n29844 & n29846;
  assign n29848 = P1_P3_INSTADDRPOINTER_REG_22_ & n29669;
  assign n29849 = ~P1_P3_INSTADDRPOINTER_REG_23_ & ~n29848;
  assign n29850 = n29669 & n29813;
  assign n29851 = ~n29849 & ~n29850;
  assign n29852 = n27741 & n29851;
  assign n29853 = ~n29834 & ~n29835;
  assign n29854 = n29838 & n29853;
  assign n29855 = n29847 & n29854;
  assign n29856 = ~n29852 & n29855;
  assign n29857 = n29821 & n29856;
  assign n29858 = n27634 & ~n29857;
  assign n4421 = ~n29785 | n29858;
  assign n29860 = P1_P3_INSTADDRPOINTER_REG_24_ & n27633;
  assign n29861 = P1_P3_REIP_REG_24_ & n27778;
  assign n29862 = ~n29860 & ~n29861;
  assign n29863 = P1_P3_INSTADDRPOINTER_REG_23_ & n29786;
  assign n29864 = ~P1_P3_INSTADDRPOINTER_REG_24_ & n29863;
  assign n29865 = P1_P3_INSTADDRPOINTER_REG_24_ & ~n29863;
  assign n29866 = ~n29864 & ~n29865;
  assign n29867 = n25739 & ~n29866;
  assign n29868 = n25731 & ~n29866;
  assign n29869 = ~n29867 & ~n29868;
  assign n29870 = P1_P3_INSTADDRPOINTER_REG_23_ & n29793;
  assign n29871 = ~P1_P3_INSTADDRPOINTER_REG_24_ & n29870;
  assign n29872 = P1_P3_INSTADDRPOINTER_REG_24_ & ~n29870;
  assign n29873 = ~n29871 & ~n29872;
  assign n29874 = n25641 & ~n29873;
  assign n29875 = n25719 & ~n29873;
  assign n29876 = n25723 & ~n29873;
  assign n29877 = ~n29874 & ~n29875;
  assign n29878 = ~n29876 & n29877;
  assign n29879 = ~P1_P3_INSTADDRPOINTER_REG_24_ & n29814;
  assign n29880 = P1_P3_INSTADDRPOINTER_REG_24_ & ~n29814;
  assign n29881 = ~n29879 & ~n29880;
  assign n29882 = n25742 & ~n29881;
  assign n29883 = P1_P3_INSTADDRPOINTER_REG_23_ & n29802;
  assign n29884 = ~P1_P3_INSTADDRPOINTER_REG_24_ & n29883;
  assign n29885 = P1_P3_INSTADDRPOINTER_REG_24_ & ~n29883;
  assign n29886 = ~n29884 & ~n29885;
  assign n29887 = n27758 & ~n29886;
  assign n29888 = ~n29882 & ~n29887;
  assign n29889 = n27747 & ~n29886;
  assign n29890 = n27751 & ~n29886;
  assign n29891 = n25785 & ~n29886;
  assign n29892 = ~n29889 & ~n29890;
  assign n29893 = ~n29891 & n29892;
  assign n29894 = n29869 & n29878;
  assign n29895 = n29888 & n29894;
  assign n29896 = n29893 & n29895;
  assign n29897 = ~P1_P3_INSTADDRPOINTER_REG_23_ & n28561;
  assign n29898 = n29823 & ~n29897;
  assign n29899 = ~n29437 & n29898;
  assign n29900 = P1_P3_INSTADDRPOINTER_REG_23_ & ~n28561;
  assign n29901 = n29826 & ~n29900;
  assign n29902 = ~n29899 & n29901;
  assign n29903 = ~P1_P3_INSTADDRPOINTER_REG_24_ & ~n28561;
  assign n29904 = P1_P3_INSTADDRPOINTER_REG_24_ & n28561;
  assign n29905 = ~n29903 & ~n29904;
  assign n29906 = n29902 & ~n29905;
  assign n29907 = ~n29902 & n29905;
  assign n29908 = ~n29906 & ~n29907;
  assign n29909 = n27739 & ~n29908;
  assign n29910 = ~n25828 & ~n29886;
  assign n29911 = n25938 & ~n29886;
  assign n29912 = n25781 & ~n29886;
  assign n29913 = ~n29911 & ~n29912;
  assign n29914 = ~P1_P3_INSTADDRPOINTER_REG_24_ & n29850;
  assign n29915 = P1_P3_INSTADDRPOINTER_REG_24_ & ~n29850;
  assign n29916 = ~n29914 & ~n29915;
  assign n29917 = n27741 & ~n29916;
  assign n29918 = n25899 & ~n29873;
  assign n29919 = n25900 & ~n29873;
  assign n29920 = n27642 & ~n29886;
  assign n29921 = n25715 & ~n29873;
  assign n29922 = n27645 & ~n29886;
  assign n29923 = ~n29921 & ~n29922;
  assign n29924 = ~n29918 & ~n29919;
  assign n29925 = ~n29920 & n29924;
  assign n29926 = n29923 & n29925;
  assign n29927 = ~n29909 & ~n29910;
  assign n29928 = n29913 & n29927;
  assign n29929 = ~n29917 & n29928;
  assign n29930 = n29926 & n29929;
  assign n29931 = n29896 & n29930;
  assign n29932 = n27634 & ~n29931;
  assign n4426 = ~n29862 | n29932;
  assign n29934 = P1_P3_INSTADDRPOINTER_REG_25_ & n27633;
  assign n29935 = P1_P3_REIP_REG_25_ & n27778;
  assign n29936 = ~n29934 & ~n29935;
  assign n29937 = P1_P3_INSTADDRPOINTER_REG_24_ & n29863;
  assign n29938 = ~P1_P3_INSTADDRPOINTER_REG_25_ & n29937;
  assign n29939 = P1_P3_INSTADDRPOINTER_REG_25_ & ~n29937;
  assign n29940 = ~n29938 & ~n29939;
  assign n29941 = n25739 & ~n29940;
  assign n29942 = n25731 & ~n29940;
  assign n29943 = ~n29941 & ~n29942;
  assign n29944 = P1_P3_INSTADDRPOINTER_REG_24_ & n29870;
  assign n29945 = ~P1_P3_INSTADDRPOINTER_REG_25_ & n29944;
  assign n29946 = P1_P3_INSTADDRPOINTER_REG_25_ & ~n29944;
  assign n29947 = ~n29945 & ~n29946;
  assign n29948 = n25641 & ~n29947;
  assign n29949 = n25719 & ~n29947;
  assign n29950 = n25723 & ~n29947;
  assign n29951 = ~n29948 & ~n29949;
  assign n29952 = ~n29950 & n29951;
  assign n29953 = P1_P3_INSTADDRPOINTER_REG_24_ & n29814;
  assign n29954 = ~P1_P3_INSTADDRPOINTER_REG_25_ & ~n29953;
  assign n29955 = P1_P3_INSTADDRPOINTER_REG_24_ & P1_P3_INSTADDRPOINTER_REG_25_;
  assign n29956 = n29814 & n29955;
  assign n29957 = ~n29954 & ~n29956;
  assign n29958 = n25742 & n29957;
  assign n29959 = P1_P3_INSTADDRPOINTER_REG_24_ & n29883;
  assign n29960 = ~P1_P3_INSTADDRPOINTER_REG_25_ & n29959;
  assign n29961 = P1_P3_INSTADDRPOINTER_REG_25_ & ~n29959;
  assign n29962 = ~n29960 & ~n29961;
  assign n29963 = n27758 & ~n29962;
  assign n29964 = ~n29958 & ~n29963;
  assign n29965 = n27747 & ~n29962;
  assign n29966 = n27751 & ~n29962;
  assign n29967 = n25785 & ~n29962;
  assign n29968 = ~n29965 & ~n29966;
  assign n29969 = ~n29967 & n29968;
  assign n29970 = n29943 & n29952;
  assign n29971 = n29964 & n29970;
  assign n29972 = n29969 & n29971;
  assign n29973 = ~P1_P3_INSTADDRPOINTER_REG_25_ & ~n28561;
  assign n29974 = P1_P3_INSTADDRPOINTER_REG_25_ & n28561;
  assign n29975 = ~n29973 & ~n29974;
  assign n29976 = P1_P3_INSTADDRPOINTER_REG_24_ & ~n28561;
  assign n29977 = n29901 & ~n29976;
  assign n29978 = ~P1_P3_INSTADDRPOINTER_REG_24_ & n28561;
  assign n29979 = n29898 & ~n29978;
  assign n29980 = ~n29437 & n29979;
  assign n29981 = n29977 & ~n29980;
  assign n29982 = ~n29975 & n29981;
  assign n29983 = ~P1_P3_INSTADDRPOINTER_REG_25_ & n28561;
  assign n29984 = P1_P3_INSTADDRPOINTER_REG_25_ & ~n28561;
  assign n29985 = ~n29983 & ~n29984;
  assign n29986 = ~n29981 & ~n29985;
  assign n29987 = ~n29982 & ~n29986;
  assign n29988 = n27739 & ~n29987;
  assign n29989 = ~n25828 & ~n29962;
  assign n29990 = P1_P3_INSTADDRPOINTER_REG_24_ & n29850;
  assign n29991 = ~P1_P3_INSTADDRPOINTER_REG_25_ & ~n29990;
  assign n29992 = n29850 & n29955;
  assign n29993 = ~n29991 & ~n29992;
  assign n29994 = n27741 & n29993;
  assign n29995 = n25938 & ~n29962;
  assign n29996 = n25781 & ~n29962;
  assign n29997 = ~n29995 & ~n29996;
  assign n29998 = n25899 & ~n29947;
  assign n29999 = n25900 & ~n29947;
  assign n30000 = n27642 & ~n29962;
  assign n30001 = n25715 & ~n29947;
  assign n30002 = n27645 & ~n29962;
  assign n30003 = ~n30001 & ~n30002;
  assign n30004 = ~n29998 & ~n29999;
  assign n30005 = ~n30000 & n30004;
  assign n30006 = n30003 & n30005;
  assign n30007 = ~n29988 & ~n29989;
  assign n30008 = ~n29994 & n30007;
  assign n30009 = n29997 & n30008;
  assign n30010 = n30006 & n30009;
  assign n30011 = n29972 & n30010;
  assign n30012 = n27634 & ~n30011;
  assign n4431 = ~n29936 | n30012;
  assign n30014 = P1_P3_INSTADDRPOINTER_REG_26_ & n27633;
  assign n30015 = P1_P3_REIP_REG_26_ & n27778;
  assign n30016 = P1_P3_INSTADDRPOINTER_REG_26_ & ~n28561;
  assign n30017 = P1_P3_INSTADDRPOINTER_REG_25_ & P1_P3_INSTADDRPOINTER_REG_26_;
  assign n30018 = n28561 & ~n30017;
  assign n30019 = ~n30016 & ~n30018;
  assign n30020 = n29981 & ~n29984;
  assign n30021 = n30019 & ~n30020;
  assign n30022 = ~P1_P3_INSTADDRPOINTER_REG_26_ & ~n28561;
  assign n30023 = P1_P3_INSTADDRPOINTER_REG_26_ & n28561;
  assign n30024 = ~n30022 & ~n30023;
  assign n30025 = ~n29984 & n30024;
  assign n30026 = ~n29981 & ~n29983;
  assign n30027 = n30025 & ~n30026;
  assign n30028 = ~n30021 & ~n30027;
  assign n30029 = n27739 & n30028;
  assign n30030 = ~P1_P3_INSTADDRPOINTER_REG_26_ & ~n29992;
  assign n30031 = P1_P3_INSTADDRPOINTER_REG_26_ & n29992;
  assign n30032 = ~n30030 & ~n30031;
  assign n30033 = n27741 & n30032;
  assign n30034 = ~n30029 & ~n30033;
  assign n30035 = P1_P3_INSTADDRPOINTER_REG_25_ & n29959;
  assign n30036 = ~P1_P3_INSTADDRPOINTER_REG_26_ & n30035;
  assign n30037 = P1_P3_INSTADDRPOINTER_REG_26_ & ~n30035;
  assign n30038 = ~n30036 & ~n30037;
  assign n30039 = ~n25828 & ~n30038;
  assign n30040 = n25938 & ~n30038;
  assign n30041 = n25781 & ~n30038;
  assign n30042 = ~n30040 & ~n30041;
  assign n30043 = P1_P3_INSTADDRPOINTER_REG_25_ & n29944;
  assign n30044 = ~P1_P3_INSTADDRPOINTER_REG_26_ & n30043;
  assign n30045 = P1_P3_INSTADDRPOINTER_REG_26_ & ~n30043;
  assign n30046 = ~n30044 & ~n30045;
  assign n30047 = n25899 & ~n30046;
  assign n30048 = n25900 & ~n30046;
  assign n30049 = n27642 & ~n30038;
  assign n30050 = n25715 & ~n30046;
  assign n30051 = n27645 & ~n30038;
  assign n30052 = ~n30050 & ~n30051;
  assign n30053 = ~n30047 & ~n30048;
  assign n30054 = ~n30049 & n30053;
  assign n30055 = n30052 & n30054;
  assign n30056 = P1_P3_INSTADDRPOINTER_REG_25_ & n29937;
  assign n30057 = ~P1_P3_INSTADDRPOINTER_REG_26_ & n30056;
  assign n30058 = P1_P3_INSTADDRPOINTER_REG_26_ & ~n30056;
  assign n30059 = ~n30057 & ~n30058;
  assign n30060 = n25739 & ~n30059;
  assign n30061 = n25731 & ~n30059;
  assign n30062 = ~n30060 & ~n30061;
  assign n30063 = n25641 & ~n30046;
  assign n30064 = n25719 & ~n30046;
  assign n30065 = n25723 & ~n30046;
  assign n30066 = ~n30063 & ~n30064;
  assign n30067 = ~n30065 & n30066;
  assign n30068 = ~P1_P3_INSTADDRPOINTER_REG_26_ & ~n29956;
  assign n30069 = P1_P3_INSTADDRPOINTER_REG_26_ & n29956;
  assign n30070 = ~n30068 & ~n30069;
  assign n30071 = n25742 & n30070;
  assign n30072 = n27758 & ~n30038;
  assign n30073 = ~n30071 & ~n30072;
  assign n30074 = n27747 & ~n30038;
  assign n30075 = n27751 & ~n30038;
  assign n30076 = n25785 & ~n30038;
  assign n30077 = ~n30074 & ~n30075;
  assign n30078 = ~n30076 & n30077;
  assign n30079 = n30062 & n30067;
  assign n30080 = n30073 & n30079;
  assign n30081 = n30078 & n30080;
  assign n30082 = n30034 & ~n30039;
  assign n30083 = n30042 & n30082;
  assign n30084 = n30055 & n30083;
  assign n30085 = n30081 & n30084;
  assign n30086 = n27634 & ~n30085;
  assign n30087 = ~n30014 & ~n30015;
  assign n4436 = n30086 | ~n30087;
  assign n30089 = P1_P3_INSTADDRPOINTER_REG_27_ & n27633;
  assign n30090 = P1_P3_REIP_REG_27_ & n27778;
  assign n30091 = ~n29984 & ~n30016;
  assign n30092 = ~n29981 & ~n30018;
  assign n30093 = n30091 & ~n30092;
  assign n30094 = ~P1_P3_INSTADDRPOINTER_REG_27_ & ~n28561;
  assign n30095 = P1_P3_INSTADDRPOINTER_REG_27_ & n28561;
  assign n30096 = ~n30094 & ~n30095;
  assign n30097 = n30093 & ~n30096;
  assign n30098 = ~n30093 & n30096;
  assign n30099 = ~n30097 & ~n30098;
  assign n30100 = n27739 & ~n30099;
  assign n30101 = ~P1_P3_INSTADDRPOINTER_REG_27_ & n30031;
  assign n30102 = P1_P3_INSTADDRPOINTER_REG_27_ & ~n30031;
  assign n30103 = ~n30101 & ~n30102;
  assign n30104 = n27741 & ~n30103;
  assign n30105 = ~n30100 & ~n30104;
  assign n30106 = P1_P3_INSTADDRPOINTER_REG_26_ & n30035;
  assign n30107 = ~P1_P3_INSTADDRPOINTER_REG_27_ & n30106;
  assign n30108 = P1_P3_INSTADDRPOINTER_REG_27_ & ~n30106;
  assign n30109 = ~n30107 & ~n30108;
  assign n30110 = ~n25828 & ~n30109;
  assign n30111 = n25938 & ~n30109;
  assign n30112 = n25781 & ~n30109;
  assign n30113 = ~n30111 & ~n30112;
  assign n30114 = P1_P3_INSTADDRPOINTER_REG_26_ & n30043;
  assign n30115 = ~P1_P3_INSTADDRPOINTER_REG_27_ & n30114;
  assign n30116 = P1_P3_INSTADDRPOINTER_REG_27_ & ~n30114;
  assign n30117 = ~n30115 & ~n30116;
  assign n30118 = n25899 & ~n30117;
  assign n30119 = n25900 & ~n30117;
  assign n30120 = n27642 & ~n30109;
  assign n30121 = n25715 & ~n30117;
  assign n30122 = n27645 & ~n30109;
  assign n30123 = ~n30121 & ~n30122;
  assign n30124 = ~n30118 & ~n30119;
  assign n30125 = ~n30120 & n30124;
  assign n30126 = n30123 & n30125;
  assign n30127 = P1_P3_INSTADDRPOINTER_REG_26_ & n30056;
  assign n30128 = ~P1_P3_INSTADDRPOINTER_REG_27_ & n30127;
  assign n30129 = P1_P3_INSTADDRPOINTER_REG_27_ & ~n30127;
  assign n30130 = ~n30128 & ~n30129;
  assign n30131 = n25739 & ~n30130;
  assign n30132 = n25731 & ~n30130;
  assign n30133 = ~n30131 & ~n30132;
  assign n30134 = n25641 & ~n30117;
  assign n30135 = n25719 & ~n30117;
  assign n30136 = n25723 & ~n30117;
  assign n30137 = ~n30134 & ~n30135;
  assign n30138 = ~n30136 & n30137;
  assign n30139 = ~P1_P3_INSTADDRPOINTER_REG_27_ & n30069;
  assign n30140 = P1_P3_INSTADDRPOINTER_REG_27_ & ~n30069;
  assign n30141 = ~n30139 & ~n30140;
  assign n30142 = n25742 & ~n30141;
  assign n30143 = n27758 & ~n30109;
  assign n30144 = ~n30142 & ~n30143;
  assign n30145 = n27747 & ~n30109;
  assign n30146 = n27751 & ~n30109;
  assign n30147 = n25785 & ~n30109;
  assign n30148 = ~n30145 & ~n30146;
  assign n30149 = ~n30147 & n30148;
  assign n30150 = n30133 & n30138;
  assign n30151 = n30144 & n30150;
  assign n30152 = n30149 & n30151;
  assign n30153 = n30105 & ~n30110;
  assign n30154 = n30113 & n30153;
  assign n30155 = n30126 & n30154;
  assign n30156 = n30152 & n30155;
  assign n30157 = n27634 & ~n30156;
  assign n30158 = ~n30089 & ~n30090;
  assign n4441 = n30157 | ~n30158;
  assign n30160 = P1_P3_INSTADDRPOINTER_REG_28_ & n27633;
  assign n30161 = P1_P3_REIP_REG_28_ & n27778;
  assign n30162 = P1_P3_INSTADDRPOINTER_REG_27_ & P1_P3_INSTADDRPOINTER_REG_28_;
  assign n30163 = ~n30093 & n30162;
  assign n30164 = n28561 & ~n30163;
  assign n30165 = P1_P3_INSTADDRPOINTER_REG_28_ & ~n28561;
  assign n30166 = ~P1_P3_INSTADDRPOINTER_REG_27_ & ~n29984;
  assign n30167 = ~n30016 & n30166;
  assign n30168 = ~n30092 & n30167;
  assign n30169 = ~n30164 & ~n30165;
  assign n30170 = ~n30168 & n30169;
  assign n30171 = P1_P3_INSTADDRPOINTER_REG_28_ & n30168;
  assign n30172 = ~n28561 & ~n30171;
  assign n30173 = P1_P3_INSTADDRPOINTER_REG_28_ & n28561;
  assign n30174 = P1_P3_INSTADDRPOINTER_REG_27_ & ~n30093;
  assign n30175 = ~n30172 & ~n30173;
  assign n30176 = ~n30174 & n30175;
  assign n30177 = ~n30170 & ~n30176;
  assign n30178 = n27739 & n30177;
  assign n30179 = P1_P3_INSTADDRPOINTER_REG_27_ & n30031;
  assign n30180 = ~P1_P3_INSTADDRPOINTER_REG_28_ & ~n30179;
  assign n30181 = n30031 & n30162;
  assign n30182 = ~n30180 & ~n30181;
  assign n30183 = n27741 & n30182;
  assign n30184 = ~n30178 & ~n30183;
  assign n30185 = P1_P3_INSTADDRPOINTER_REG_27_ & n30106;
  assign n30186 = ~P1_P3_INSTADDRPOINTER_REG_28_ & n30185;
  assign n30187 = P1_P3_INSTADDRPOINTER_REG_28_ & ~n30185;
  assign n30188 = ~n30186 & ~n30187;
  assign n30189 = ~n25828 & ~n30188;
  assign n30190 = n25938 & ~n30188;
  assign n30191 = n25781 & ~n30188;
  assign n30192 = ~n30190 & ~n30191;
  assign n30193 = P1_P3_INSTADDRPOINTER_REG_27_ & n30114;
  assign n30194 = ~P1_P3_INSTADDRPOINTER_REG_28_ & n30193;
  assign n30195 = P1_P3_INSTADDRPOINTER_REG_28_ & ~n30193;
  assign n30196 = ~n30194 & ~n30195;
  assign n30197 = n25899 & ~n30196;
  assign n30198 = n25900 & ~n30196;
  assign n30199 = n27642 & ~n30188;
  assign n30200 = n25715 & ~n30196;
  assign n30201 = n27645 & ~n30188;
  assign n30202 = ~n30200 & ~n30201;
  assign n30203 = ~n30197 & ~n30198;
  assign n30204 = ~n30199 & n30203;
  assign n30205 = n30202 & n30204;
  assign n30206 = P1_P3_INSTADDRPOINTER_REG_27_ & n30127;
  assign n30207 = ~P1_P3_INSTADDRPOINTER_REG_28_ & n30206;
  assign n30208 = P1_P3_INSTADDRPOINTER_REG_28_ & ~n30206;
  assign n30209 = ~n30207 & ~n30208;
  assign n30210 = n25739 & ~n30209;
  assign n30211 = n25731 & ~n30209;
  assign n30212 = ~n30210 & ~n30211;
  assign n30213 = n25641 & ~n30196;
  assign n30214 = n25719 & ~n30196;
  assign n30215 = n25723 & ~n30196;
  assign n30216 = ~n30213 & ~n30214;
  assign n30217 = ~n30215 & n30216;
  assign n30218 = P1_P3_INSTADDRPOINTER_REG_27_ & n30069;
  assign n30219 = ~P1_P3_INSTADDRPOINTER_REG_28_ & ~n30218;
  assign n30220 = n30069 & n30162;
  assign n30221 = ~n30219 & ~n30220;
  assign n30222 = n25742 & n30221;
  assign n30223 = n27758 & ~n30188;
  assign n30224 = ~n30222 & ~n30223;
  assign n30225 = n27747 & ~n30188;
  assign n30226 = n27751 & ~n30188;
  assign n30227 = n25785 & ~n30188;
  assign n30228 = ~n30225 & ~n30226;
  assign n30229 = ~n30227 & n30228;
  assign n30230 = n30212 & n30217;
  assign n30231 = n30224 & n30230;
  assign n30232 = n30229 & n30231;
  assign n30233 = n30184 & ~n30189;
  assign n30234 = n30192 & n30233;
  assign n30235 = n30205 & n30234;
  assign n30236 = n30232 & n30235;
  assign n30237 = n27634 & ~n30236;
  assign n30238 = ~n30160 & ~n30161;
  assign n4446 = n30237 | ~n30238;
  assign n30240 = P1_P3_INSTADDRPOINTER_REG_29_ & n27633;
  assign n30241 = P1_P3_REIP_REG_29_ & n27778;
  assign n30242 = ~n28561 & ~n30168;
  assign n30243 = ~n30165 & ~n30242;
  assign n30244 = ~n30163 & n30243;
  assign n30245 = P1_P3_INSTADDRPOINTER_REG_29_ & n28561;
  assign n30246 = ~P1_P3_INSTADDRPOINTER_REG_29_ & ~n28561;
  assign n30247 = ~n30245 & ~n30246;
  assign n30248 = n30244 & ~n30247;
  assign n30249 = ~n30244 & n30247;
  assign n30250 = ~n30248 & ~n30249;
  assign n30251 = n27739 & ~n30250;
  assign n30252 = ~P1_P3_INSTADDRPOINTER_REG_29_ & ~n30181;
  assign n30253 = P1_P3_INSTADDRPOINTER_REG_29_ & n30181;
  assign n30254 = ~n30252 & ~n30253;
  assign n30255 = n27741 & n30254;
  assign n30256 = ~n30251 & ~n30255;
  assign n30257 = P1_P3_INSTADDRPOINTER_REG_28_ & n30185;
  assign n30258 = ~P1_P3_INSTADDRPOINTER_REG_29_ & n30257;
  assign n30259 = P1_P3_INSTADDRPOINTER_REG_29_ & ~n30257;
  assign n30260 = ~n30258 & ~n30259;
  assign n30261 = ~n25828 & ~n30260;
  assign n30262 = n25938 & ~n30260;
  assign n30263 = n25781 & ~n30260;
  assign n30264 = ~n30262 & ~n30263;
  assign n30265 = P1_P3_INSTADDRPOINTER_REG_28_ & n30193;
  assign n30266 = ~P1_P3_INSTADDRPOINTER_REG_29_ & n30265;
  assign n30267 = P1_P3_INSTADDRPOINTER_REG_29_ & ~n30265;
  assign n30268 = ~n30266 & ~n30267;
  assign n30269 = n25899 & ~n30268;
  assign n30270 = n25900 & ~n30268;
  assign n30271 = n27642 & ~n30260;
  assign n30272 = n25715 & ~n30268;
  assign n30273 = n27645 & ~n30260;
  assign n30274 = ~n30272 & ~n30273;
  assign n30275 = ~n30269 & ~n30270;
  assign n30276 = ~n30271 & n30275;
  assign n30277 = n30274 & n30276;
  assign n30278 = P1_P3_INSTADDRPOINTER_REG_28_ & n30206;
  assign n30279 = ~P1_P3_INSTADDRPOINTER_REG_29_ & n30278;
  assign n30280 = P1_P3_INSTADDRPOINTER_REG_29_ & ~n30278;
  assign n30281 = ~n30279 & ~n30280;
  assign n30282 = n25739 & ~n30281;
  assign n30283 = n25731 & ~n30281;
  assign n30284 = ~n30282 & ~n30283;
  assign n30285 = n25641 & ~n30268;
  assign n30286 = n25719 & ~n30268;
  assign n30287 = n25723 & ~n30268;
  assign n30288 = ~n30285 & ~n30286;
  assign n30289 = ~n30287 & n30288;
  assign n30290 = ~P1_P3_INSTADDRPOINTER_REG_29_ & ~n30220;
  assign n30291 = P1_P3_INSTADDRPOINTER_REG_29_ & n30220;
  assign n30292 = ~n30290 & ~n30291;
  assign n30293 = n25742 & n30292;
  assign n30294 = n27758 & ~n30260;
  assign n30295 = ~n30293 & ~n30294;
  assign n30296 = n27747 & ~n30260;
  assign n30297 = n27751 & ~n30260;
  assign n30298 = n25785 & ~n30260;
  assign n30299 = ~n30296 & ~n30297;
  assign n30300 = ~n30298 & n30299;
  assign n30301 = n30284 & n30289;
  assign n30302 = n30295 & n30301;
  assign n30303 = n30300 & n30302;
  assign n30304 = n30256 & ~n30261;
  assign n30305 = n30264 & n30304;
  assign n30306 = n30277 & n30305;
  assign n30307 = n30303 & n30306;
  assign n30308 = n27634 & ~n30307;
  assign n30309 = ~n30240 & ~n30241;
  assign n4451 = n30308 | ~n30309;
  assign n30311 = P1_P3_INSTADDRPOINTER_REG_30_ & n27633;
  assign n30312 = P1_P3_REIP_REG_30_ & n27778;
  assign n30313 = P1_P3_INSTADDRPOINTER_REG_30_ & n28561;
  assign n30314 = ~P1_P3_INSTADDRPOINTER_REG_30_ & ~n28561;
  assign n30315 = ~n30313 & ~n30314;
  assign n30316 = P1_P3_INSTADDRPOINTER_REG_29_ & ~n30244;
  assign n30317 = ~n28561 & ~n30244;
  assign n30318 = P1_P3_INSTADDRPOINTER_REG_29_ & ~n28561;
  assign n30319 = ~n30316 & ~n30317;
  assign n30320 = ~n30318 & n30319;
  assign n30321 = ~n30315 & n30320;
  assign n30322 = n30315 & ~n30320;
  assign n30323 = ~n30321 & ~n30322;
  assign n30324 = n27739 & ~n30323;
  assign n30325 = ~P1_P3_INSTADDRPOINTER_REG_30_ & n30253;
  assign n30326 = P1_P3_INSTADDRPOINTER_REG_30_ & ~n30253;
  assign n30327 = ~n30325 & ~n30326;
  assign n30328 = n27741 & ~n30327;
  assign n30329 = ~n30324 & ~n30328;
  assign n30330 = P1_P3_INSTADDRPOINTER_REG_29_ & n30257;
  assign n30331 = ~P1_P3_INSTADDRPOINTER_REG_30_ & n30330;
  assign n30332 = P1_P3_INSTADDRPOINTER_REG_30_ & ~n30330;
  assign n30333 = ~n30331 & ~n30332;
  assign n30334 = ~n25828 & ~n30333;
  assign n30335 = n25938 & ~n30333;
  assign n30336 = n25781 & ~n30333;
  assign n30337 = ~n30335 & ~n30336;
  assign n30338 = P1_P3_INSTADDRPOINTER_REG_29_ & n30265;
  assign n30339 = ~P1_P3_INSTADDRPOINTER_REG_30_ & n30338;
  assign n30340 = P1_P3_INSTADDRPOINTER_REG_30_ & ~n30338;
  assign n30341 = ~n30339 & ~n30340;
  assign n30342 = n25899 & ~n30341;
  assign n30343 = n25900 & ~n30341;
  assign n30344 = n27642 & ~n30333;
  assign n30345 = n25715 & ~n30341;
  assign n30346 = n27645 & ~n30333;
  assign n30347 = ~n30345 & ~n30346;
  assign n30348 = ~n30342 & ~n30343;
  assign n30349 = ~n30344 & n30348;
  assign n30350 = n30347 & n30349;
  assign n30351 = P1_P3_INSTADDRPOINTER_REG_29_ & n30278;
  assign n30352 = ~P1_P3_INSTADDRPOINTER_REG_30_ & n30351;
  assign n30353 = P1_P3_INSTADDRPOINTER_REG_30_ & ~n30351;
  assign n30354 = ~n30352 & ~n30353;
  assign n30355 = n25739 & ~n30354;
  assign n30356 = n25731 & ~n30354;
  assign n30357 = ~n30355 & ~n30356;
  assign n30358 = n25641 & ~n30341;
  assign n30359 = n25719 & ~n30341;
  assign n30360 = n25723 & ~n30341;
  assign n30361 = ~n30358 & ~n30359;
  assign n30362 = ~n30360 & n30361;
  assign n30363 = ~P1_P3_INSTADDRPOINTER_REG_30_ & n30291;
  assign n30364 = P1_P3_INSTADDRPOINTER_REG_30_ & ~n30291;
  assign n30365 = ~n30363 & ~n30364;
  assign n30366 = n25742 & ~n30365;
  assign n30367 = n27758 & ~n30333;
  assign n30368 = ~n30366 & ~n30367;
  assign n30369 = n27747 & ~n30333;
  assign n30370 = n27751 & ~n30333;
  assign n30371 = n25785 & ~n30333;
  assign n30372 = ~n30369 & ~n30370;
  assign n30373 = ~n30371 & n30372;
  assign n30374 = n30357 & n30362;
  assign n30375 = n30368 & n30374;
  assign n30376 = n30373 & n30375;
  assign n30377 = n30329 & ~n30334;
  assign n30378 = n30337 & n30377;
  assign n30379 = n30350 & n30378;
  assign n30380 = n30376 & n30379;
  assign n30381 = n27634 & ~n30380;
  assign n30382 = ~n30311 & ~n30312;
  assign n4456 = n30381 | ~n30382;
  assign n30384 = P1_P3_INSTADDRPOINTER_REG_31_ & n27633;
  assign n30385 = P1_P3_REIP_REG_31_ & n27778;
  assign n30386 = P1_P3_INSTADDRPOINTER_REG_30_ & n30291;
  assign n30387 = ~P1_P3_INSTADDRPOINTER_REG_31_ & n30386;
  assign n30388 = P1_P3_INSTADDRPOINTER_REG_31_ & ~n30386;
  assign n30389 = ~n30387 & ~n30388;
  assign n30390 = n25742 & ~n30389;
  assign n30391 = P1_P3_INSTADDRPOINTER_REG_30_ & n30330;
  assign n30392 = ~P1_P3_INSTADDRPOINTER_REG_31_ & n30391;
  assign n30393 = P1_P3_INSTADDRPOINTER_REG_31_ & ~n30391;
  assign n30394 = ~n30392 & ~n30393;
  assign n30395 = n27758 & ~n30394;
  assign n30396 = n25785 & ~n30394;
  assign n30397 = ~n30395 & ~n30396;
  assign n30398 = P1_P3_INSTADDRPOINTER_REG_30_ & n30338;
  assign n30399 = ~P1_P3_INSTADDRPOINTER_REG_31_ & n30398;
  assign n30400 = P1_P3_INSTADDRPOINTER_REG_31_ & ~n30398;
  assign n30401 = ~n30399 & ~n30400;
  assign n30402 = n25723 & ~n30401;
  assign n30403 = n25641 & ~n30401;
  assign n30404 = P1_P3_INSTADDRPOINTER_REG_30_ & n30351;
  assign n30405 = ~P1_P3_INSTADDRPOINTER_REG_31_ & n30404;
  assign n30406 = P1_P3_INSTADDRPOINTER_REG_31_ & ~n30404;
  assign n30407 = ~n30405 & ~n30406;
  assign n30408 = n25731 & ~n30407;
  assign n30409 = ~n30402 & ~n30403;
  assign n30410 = ~n30408 & n30409;
  assign n30411 = n27747 & ~n30394;
  assign n30412 = n27751 & ~n30394;
  assign n30413 = n25739 & ~n30407;
  assign n30414 = ~n30412 & ~n30413;
  assign n30415 = n30410 & ~n30411;
  assign n30416 = n30414 & n30415;
  assign n30417 = ~n30384 & ~n30385;
  assign n30418 = ~n30390 & n30417;
  assign n30419 = n30397 & n30418;
  assign n30420 = n30416 & n30419;
  assign n30421 = P1_P3_INSTADDRPOINTER_REG_30_ & P1_P3_INSTADDRPOINTER_REG_31_;
  assign n30422 = ~n30320 & n30421;
  assign n30423 = n28561 & ~n30422;
  assign n30424 = P1_P3_INSTADDRPOINTER_REG_31_ & ~n28561;
  assign n30425 = ~P1_P3_INSTADDRPOINTER_REG_30_ & n30320;
  assign n30426 = ~n30423 & ~n30424;
  assign n30427 = ~n30425 & n30426;
  assign n30428 = ~P1_P3_INSTADDRPOINTER_REG_30_ & P1_P3_INSTADDRPOINTER_REG_31_;
  assign n30429 = ~n30318 & n30428;
  assign n30430 = ~n30317 & n30429;
  assign n30431 = ~n28561 & ~n30430;
  assign n30432 = P1_P3_INSTADDRPOINTER_REG_31_ & n28561;
  assign n30433 = P1_P3_INSTADDRPOINTER_REG_30_ & ~n30320;
  assign n30434 = ~n30431 & ~n30432;
  assign n30435 = ~n30433 & n30434;
  assign n30436 = ~n30427 & ~n30435;
  assign n30437 = n27739 & n30436;
  assign n30438 = P1_P3_INSTADDRPOINTER_REG_30_ & n30253;
  assign n30439 = ~P1_P3_INSTADDRPOINTER_REG_31_ & n30438;
  assign n30440 = P1_P3_INSTADDRPOINTER_REG_31_ & ~n30438;
  assign n30441 = ~n30439 & ~n30440;
  assign n30442 = n27741 & ~n30441;
  assign n30443 = ~n30437 & ~n30442;
  assign n30444 = ~n25828 & ~n30394;
  assign n30445 = n25938 & ~n30394;
  assign n30446 = n25781 & ~n30394;
  assign n30447 = ~n30445 & ~n30446;
  assign n30448 = n25900 & ~n30401;
  assign n30449 = n30447 & ~n30448;
  assign n30450 = n27642 & ~n30394;
  assign n30451 = n25899 & ~n30401;
  assign n30452 = n25719 & ~n30401;
  assign n30453 = n25715 & ~n30401;
  assign n30454 = n27645 & ~n30394;
  assign n30455 = ~n30452 & ~n30453;
  assign n30456 = ~n30454 & n30455;
  assign n30457 = ~n30450 & ~n30451;
  assign n30458 = n30456 & n30457;
  assign n30459 = n30443 & ~n30444;
  assign n30460 = n30449 & n30459;
  assign n30461 = n30458 & n30460;
  assign n30462 = n30420 & n30461;
  assign n30463 = ~n27634 & ~n30384;
  assign n30464 = ~n30385 & n30463;
  assign n4461 = ~n30462 & ~n30464;
  assign n30466 = P1_P3_STATE2_REG_0_ & ~n25608;
  assign n30467 = ~P1_P3_STATE2_REG_0_ & ~n27601;
  assign n30468 = n25742 & n25745;
  assign n30469 = n25747 & n25751;
  assign n30470 = ~n30468 & ~n30469;
  assign n30471 = n25994 & ~n30470;
  assign n30472 = ~n30467 & ~n30471;
  assign n30473 = n30466 & ~n30472;
  assign n30474 = ~n27738 & n30473;
  assign n30475 = ~n27707 & n30474;
  assign n30476 = n27738 & n30473;
  assign n30477 = ~n27707 & n30476;
  assign n30478 = P1_P3_STATE2_REG_1_ & ~n30472;
  assign n30479 = P1_P3_STATEBS16_REG & n30478;
  assign n30480 = P1_P3_PHYADDRPOINTER_REG_0_ & n30479;
  assign n30481 = ~P1_P3_STATEBS16_REG & n30478;
  assign n30482 = P1_P3_PHYADDRPOINTER_REG_0_ & n30481;
  assign n30483 = P1_P3_PHYADDRPOINTER_REG_0_ & n30472;
  assign n30484 = P1_P3_STATE2_REG_0_ & n25608;
  assign n30485 = ~n30472 & n30484;
  assign n30486 = ~n27755 & n30485;
  assign n30487 = P1_P3_STATE2_REG_2_ & ~P1_P3_STATE2_REG_0_;
  assign n30488 = ~n30472 & n30487;
  assign n30489 = P1_P3_PHYADDRPOINTER_REG_0_ & n30488;
  assign n30490 = n26010 & ~n30472;
  assign n30491 = P1_P3_REIP_REG_0_ & n30490;
  assign n30492 = ~n30483 & ~n30486;
  assign n30493 = ~n30489 & n30492;
  assign n30494 = ~n30491 & n30493;
  assign n30495 = ~n30475 & ~n30477;
  assign n30496 = ~n30480 & n30495;
  assign n30497 = ~n30482 & n30496;
  assign n4466 = ~n30494 | ~n30497;
  assign n30499 = ~n27829 & n30474;
  assign n30500 = ~n27829 & n30476;
  assign n30501 = P1_P3_PHYADDRPOINTER_REG_1_ & n30479;
  assign n30502 = ~P1_P3_PHYADDRPOINTER_REG_1_ & n30481;
  assign n30503 = P1_P3_PHYADDRPOINTER_REG_1_ & n30472;
  assign n30504 = ~n27859 & n30485;
  assign n30505 = ~P1_P3_PHYADDRPOINTER_REG_1_ & n30488;
  assign n30506 = P1_P3_REIP_REG_1_ & n30490;
  assign n30507 = ~n30503 & ~n30504;
  assign n30508 = ~n30505 & n30507;
  assign n30509 = ~n30506 & n30508;
  assign n30510 = ~n30499 & ~n30500;
  assign n30511 = ~n30501 & n30510;
  assign n30512 = ~n30502 & n30511;
  assign n4471 = ~n30509 | ~n30512;
  assign n30514 = ~n27956 & n30474;
  assign n30515 = ~n27942 & n30476;
  assign n30516 = ~P1_P3_PHYADDRPOINTER_REG_2_ & n30479;
  assign n30517 = P1_P3_PHYADDRPOINTER_REG_1_ & ~P1_P3_PHYADDRPOINTER_REG_2_;
  assign n30518 = ~P1_P3_PHYADDRPOINTER_REG_1_ & P1_P3_PHYADDRPOINTER_REG_2_;
  assign n30519 = ~n30517 & ~n30518;
  assign n30520 = n30481 & ~n30519;
  assign n30521 = n30488 & ~n30519;
  assign n30522 = P1_P3_REIP_REG_2_ & n30490;
  assign n30523 = P1_P3_PHYADDRPOINTER_REG_2_ & n30472;
  assign n30524 = ~n27993 & n30485;
  assign n30525 = ~n30521 & ~n30522;
  assign n30526 = ~n30523 & n30525;
  assign n30527 = ~n30524 & n30526;
  assign n30528 = ~n30514 & ~n30515;
  assign n30529 = ~n30516 & n30528;
  assign n30530 = ~n30520 & n30529;
  assign n4476 = ~n30527 | ~n30530;
  assign n30532 = ~n28071 & n30474;
  assign n30533 = n28086 & n30476;
  assign n30534 = P1_P3_PHYADDRPOINTER_REG_2_ & ~P1_P3_PHYADDRPOINTER_REG_3_;
  assign n30535 = ~P1_P3_PHYADDRPOINTER_REG_2_ & P1_P3_PHYADDRPOINTER_REG_3_;
  assign n30536 = ~n30534 & ~n30535;
  assign n30537 = n30479 & ~n30536;
  assign n30538 = P1_P3_PHYADDRPOINTER_REG_1_ & P1_P3_PHYADDRPOINTER_REG_2_;
  assign n30539 = ~P1_P3_PHYADDRPOINTER_REG_3_ & n30538;
  assign n30540 = P1_P3_PHYADDRPOINTER_REG_3_ & ~n30538;
  assign n30541 = ~n30539 & ~n30540;
  assign n30542 = n30481 & ~n30541;
  assign n30543 = n30488 & ~n30541;
  assign n30544 = P1_P3_REIP_REG_3_ & n30490;
  assign n30545 = P1_P3_PHYADDRPOINTER_REG_3_ & n30472;
  assign n30546 = n28124 & n30485;
  assign n30547 = ~n30543 & ~n30544;
  assign n30548 = ~n30545 & n30547;
  assign n30549 = ~n30546 & n30548;
  assign n30550 = ~n30532 & ~n30533;
  assign n30551 = ~n30537 & n30550;
  assign n30552 = ~n30542 & n30551;
  assign n4481 = ~n30549 | ~n30552;
  assign n30554 = P1_P3_PHYADDRPOINTER_REG_2_ & P1_P3_PHYADDRPOINTER_REG_3_;
  assign n30555 = ~P1_P3_PHYADDRPOINTER_REG_4_ & n30554;
  assign n30556 = P1_P3_PHYADDRPOINTER_REG_4_ & ~n30554;
  assign n30557 = ~n30555 & ~n30556;
  assign n30558 = n30479 & ~n30557;
  assign n30559 = P1_P3_PHYADDRPOINTER_REG_3_ & n30538;
  assign n30560 = ~P1_P3_PHYADDRPOINTER_REG_4_ & n30559;
  assign n30561 = P1_P3_PHYADDRPOINTER_REG_4_ & ~n30559;
  assign n30562 = ~n30560 & ~n30561;
  assign n30563 = n30481 & ~n30562;
  assign n30564 = n28199 & n30476;
  assign n30565 = ~n28221 & n30474;
  assign n30566 = n30488 & ~n30562;
  assign n30567 = P1_P3_REIP_REG_4_ & n30490;
  assign n30568 = P1_P3_PHYADDRPOINTER_REG_4_ & n30472;
  assign n30569 = ~n28260 & n30485;
  assign n30570 = ~n30566 & ~n30567;
  assign n30571 = ~n30568 & n30570;
  assign n30572 = ~n30569 & n30571;
  assign n30573 = ~n30558 & ~n30563;
  assign n30574 = ~n30564 & n30573;
  assign n30575 = ~n30565 & n30574;
  assign n4486 = ~n30572 | ~n30575;
  assign n30577 = P1_P3_PHYADDRPOINTER_REG_4_ & n30554;
  assign n30578 = ~P1_P3_PHYADDRPOINTER_REG_5_ & n30577;
  assign n30579 = P1_P3_PHYADDRPOINTER_REG_5_ & ~n30577;
  assign n30580 = ~n30578 & ~n30579;
  assign n30581 = n30479 & ~n30580;
  assign n30582 = P1_P3_PHYADDRPOINTER_REG_4_ & n30559;
  assign n30583 = ~P1_P3_PHYADDRPOINTER_REG_5_ & n30582;
  assign n30584 = P1_P3_PHYADDRPOINTER_REG_5_ & ~n30582;
  assign n30585 = ~n30583 & ~n30584;
  assign n30586 = n30481 & ~n30585;
  assign n30587 = ~n28336 & n30474;
  assign n30588 = ~n28354 & n30476;
  assign n30589 = n30488 & ~n30585;
  assign n30590 = P1_P3_REIP_REG_5_ & n30490;
  assign n30591 = P1_P3_PHYADDRPOINTER_REG_5_ & n30472;
  assign n30592 = n28393 & n30485;
  assign n30593 = ~n30589 & ~n30590;
  assign n30594 = ~n30591 & n30593;
  assign n30595 = ~n30592 & n30594;
  assign n30596 = ~n30581 & ~n30586;
  assign n30597 = ~n30587 & n30596;
  assign n30598 = ~n30588 & n30597;
  assign n4491 = ~n30595 | ~n30598;
  assign n30600 = P1_P3_PHYADDRPOINTER_REG_5_ & n30577;
  assign n30601 = ~P1_P3_PHYADDRPOINTER_REG_6_ & n30600;
  assign n30602 = P1_P3_PHYADDRPOINTER_REG_6_ & ~n30600;
  assign n30603 = ~n30601 & ~n30602;
  assign n30604 = n30479 & ~n30603;
  assign n30605 = P1_P3_PHYADDRPOINTER_REG_5_ & n30582;
  assign n30606 = ~P1_P3_PHYADDRPOINTER_REG_6_ & n30605;
  assign n30607 = P1_P3_PHYADDRPOINTER_REG_6_ & ~n30605;
  assign n30608 = ~n30606 & ~n30607;
  assign n30609 = n30481 & ~n30608;
  assign n30610 = ~n28467 & n30474;
  assign n30611 = ~n28486 & n30476;
  assign n30612 = n30488 & ~n30608;
  assign n30613 = P1_P3_REIP_REG_6_ & n30490;
  assign n30614 = P1_P3_PHYADDRPOINTER_REG_6_ & n30472;
  assign n30615 = ~n28524 & n30485;
  assign n30616 = ~n30612 & ~n30613;
  assign n30617 = ~n30614 & n30616;
  assign n30618 = ~n30615 & n30617;
  assign n30619 = ~n30604 & ~n30609;
  assign n30620 = ~n30610 & n30619;
  assign n30621 = ~n30611 & n30620;
  assign n4496 = ~n30618 | ~n30621;
  assign n30623 = P1_P3_PHYADDRPOINTER_REG_6_ & n30600;
  assign n30624 = ~P1_P3_PHYADDRPOINTER_REG_7_ & n30623;
  assign n30625 = P1_P3_PHYADDRPOINTER_REG_7_ & ~n30623;
  assign n30626 = ~n30624 & ~n30625;
  assign n30627 = n30479 & ~n30626;
  assign n30628 = P1_P3_PHYADDRPOINTER_REG_6_ & n30605;
  assign n30629 = ~P1_P3_PHYADDRPOINTER_REG_7_ & n30628;
  assign n30630 = P1_P3_PHYADDRPOINTER_REG_7_ & ~n30628;
  assign n30631 = ~n30629 & ~n30630;
  assign n30632 = n30481 & ~n30631;
  assign n30633 = ~n28568 & n30474;
  assign n30634 = ~n28586 & n30476;
  assign n30635 = n30488 & ~n30631;
  assign n30636 = P1_P3_REIP_REG_7_ & n30490;
  assign n30637 = P1_P3_PHYADDRPOINTER_REG_7_ & n30472;
  assign n30638 = ~n28622 & n30485;
  assign n30639 = ~n30635 & ~n30636;
  assign n30640 = ~n30637 & n30639;
  assign n30641 = ~n30638 & n30640;
  assign n30642 = ~n30627 & ~n30632;
  assign n30643 = ~n30633 & n30642;
  assign n30644 = ~n30634 & n30643;
  assign n4501 = ~n30641 | ~n30644;
  assign n30646 = P1_P3_PHYADDRPOINTER_REG_7_ & n30623;
  assign n30647 = ~P1_P3_PHYADDRPOINTER_REG_8_ & n30646;
  assign n30648 = P1_P3_PHYADDRPOINTER_REG_8_ & ~n30646;
  assign n30649 = ~n30647 & ~n30648;
  assign n30650 = n30479 & ~n30649;
  assign n30651 = P1_P3_PHYADDRPOINTER_REG_7_ & n30628;
  assign n30652 = ~P1_P3_PHYADDRPOINTER_REG_8_ & n30651;
  assign n30653 = P1_P3_PHYADDRPOINTER_REG_8_ & ~n30651;
  assign n30654 = ~n30652 & ~n30653;
  assign n30655 = n30481 & ~n30654;
  assign n30656 = ~n28662 & n30474;
  assign n30657 = ~n28678 & n30476;
  assign n30658 = n30488 & ~n30654;
  assign n30659 = P1_P3_REIP_REG_8_ & n30490;
  assign n30660 = P1_P3_PHYADDRPOINTER_REG_8_ & n30472;
  assign n30661 = ~n28712 & n30485;
  assign n30662 = ~n30658 & ~n30659;
  assign n30663 = ~n30660 & n30662;
  assign n30664 = ~n30661 & n30663;
  assign n30665 = ~n30650 & ~n30655;
  assign n30666 = ~n30656 & n30665;
  assign n30667 = ~n30657 & n30666;
  assign n4506 = ~n30664 | ~n30667;
  assign n30669 = P1_P3_PHYADDRPOINTER_REG_8_ & n30646;
  assign n30670 = ~P1_P3_PHYADDRPOINTER_REG_9_ & n30669;
  assign n30671 = P1_P3_PHYADDRPOINTER_REG_9_ & ~n30669;
  assign n30672 = ~n30670 & ~n30671;
  assign n30673 = n30479 & ~n30672;
  assign n30674 = P1_P3_PHYADDRPOINTER_REG_8_ & n30651;
  assign n30675 = ~P1_P3_PHYADDRPOINTER_REG_9_ & n30674;
  assign n30676 = P1_P3_PHYADDRPOINTER_REG_9_ & ~n30674;
  assign n30677 = ~n30675 & ~n30676;
  assign n30678 = n30481 & ~n30677;
  assign n30679 = ~n28756 & n30474;
  assign n30680 = n28767 & n30476;
  assign n30681 = n30488 & ~n30677;
  assign n30682 = P1_P3_REIP_REG_9_ & n30490;
  assign n30683 = P1_P3_PHYADDRPOINTER_REG_9_ & n30472;
  assign n30684 = n28796 & n30485;
  assign n30685 = ~n30681 & ~n30682;
  assign n30686 = ~n30683 & n30685;
  assign n30687 = ~n30684 & n30686;
  assign n30688 = ~n30673 & ~n30678;
  assign n30689 = ~n30679 & n30688;
  assign n30690 = ~n30680 & n30689;
  assign n4511 = ~n30687 | ~n30690;
  assign n30692 = P1_P3_PHYADDRPOINTER_REG_9_ & n30669;
  assign n30693 = ~P1_P3_PHYADDRPOINTER_REG_10_ & n30692;
  assign n30694 = P1_P3_PHYADDRPOINTER_REG_10_ & ~n30692;
  assign n30695 = ~n30693 & ~n30694;
  assign n30696 = n30479 & ~n30695;
  assign n30697 = P1_P3_PHYADDRPOINTER_REG_9_ & n30674;
  assign n30698 = ~P1_P3_PHYADDRPOINTER_REG_10_ & n30697;
  assign n30699 = P1_P3_PHYADDRPOINTER_REG_10_ & ~n30697;
  assign n30700 = ~n30698 & ~n30699;
  assign n30701 = n30481 & ~n30700;
  assign n30702 = n28830 & n30476;
  assign n30703 = ~n28871 & n30474;
  assign n30704 = n30488 & ~n30700;
  assign n30705 = P1_P3_REIP_REG_10_ & n30490;
  assign n30706 = P1_P3_PHYADDRPOINTER_REG_10_ & n30472;
  assign n30707 = n28854 & n30485;
  assign n30708 = ~n30704 & ~n30705;
  assign n30709 = ~n30706 & n30708;
  assign n30710 = ~n30707 & n30709;
  assign n30711 = ~n30696 & ~n30701;
  assign n30712 = ~n30702 & n30711;
  assign n30713 = ~n30703 & n30712;
  assign n4516 = ~n30710 | ~n30713;
  assign n30715 = P1_P3_PHYADDRPOINTER_REG_10_ & n30692;
  assign n30716 = ~P1_P3_PHYADDRPOINTER_REG_11_ & n30715;
  assign n30717 = P1_P3_PHYADDRPOINTER_REG_11_ & ~n30715;
  assign n30718 = ~n30716 & ~n30717;
  assign n30719 = n30479 & ~n30718;
  assign n30720 = P1_P3_PHYADDRPOINTER_REG_10_ & n30697;
  assign n30721 = ~P1_P3_PHYADDRPOINTER_REG_11_ & n30720;
  assign n30722 = P1_P3_PHYADDRPOINTER_REG_11_ & ~n30720;
  assign n30723 = ~n30721 & ~n30722;
  assign n30724 = n30481 & ~n30723;
  assign n30725 = ~n28903 & n30476;
  assign n30726 = ~n28917 & n30474;
  assign n30727 = n30488 & ~n30723;
  assign n30728 = P1_P3_REIP_REG_11_ & n30490;
  assign n30729 = P1_P3_PHYADDRPOINTER_REG_11_ & n30472;
  assign n30730 = ~n28942 & n30485;
  assign n30731 = ~n30727 & ~n30728;
  assign n30732 = ~n30729 & n30731;
  assign n30733 = ~n30730 & n30732;
  assign n30734 = ~n30719 & ~n30724;
  assign n30735 = ~n30725 & n30734;
  assign n30736 = ~n30726 & n30735;
  assign n4521 = ~n30733 | ~n30736;
  assign n30738 = P1_P3_PHYADDRPOINTER_REG_11_ & n30715;
  assign n30739 = ~P1_P3_PHYADDRPOINTER_REG_12_ & n30738;
  assign n30740 = P1_P3_PHYADDRPOINTER_REG_12_ & ~n30738;
  assign n30741 = ~n30739 & ~n30740;
  assign n30742 = n30479 & ~n30741;
  assign n30743 = P1_P3_PHYADDRPOINTER_REG_11_ & n30720;
  assign n30744 = ~P1_P3_PHYADDRPOINTER_REG_12_ & n30743;
  assign n30745 = P1_P3_PHYADDRPOINTER_REG_12_ & ~n30743;
  assign n30746 = ~n30744 & ~n30745;
  assign n30747 = n30481 & ~n30746;
  assign n30748 = ~n28987 & n30474;
  assign n30749 = n28996 & n30476;
  assign n30750 = P1_P3_PHYADDRPOINTER_REG_12_ & n30472;
  assign n30751 = P1_P3_REIP_REG_12_ & n30490;
  assign n30752 = n30488 & ~n30746;
  assign n30753 = n29022 & n30485;
  assign n30754 = ~n30750 & ~n30751;
  assign n30755 = ~n30752 & n30754;
  assign n30756 = ~n30753 & n30755;
  assign n30757 = ~n30742 & ~n30747;
  assign n30758 = ~n30748 & n30757;
  assign n30759 = ~n30749 & n30758;
  assign n4526 = ~n30756 | ~n30759;
  assign n30761 = P1_P3_PHYADDRPOINTER_REG_12_ & n30738;
  assign n30762 = ~P1_P3_PHYADDRPOINTER_REG_13_ & n30761;
  assign n30763 = P1_P3_PHYADDRPOINTER_REG_13_ & ~n30761;
  assign n30764 = ~n30762 & ~n30763;
  assign n30765 = n30479 & ~n30764;
  assign n30766 = P1_P3_PHYADDRPOINTER_REG_12_ & n30743;
  assign n30767 = ~P1_P3_PHYADDRPOINTER_REG_13_ & n30766;
  assign n30768 = P1_P3_PHYADDRPOINTER_REG_13_ & ~n30766;
  assign n30769 = ~n30767 & ~n30768;
  assign n30770 = n30481 & ~n30769;
  assign n30771 = n29065 & n30474;
  assign n30772 = n29072 & n30476;
  assign n30773 = P1_P3_PHYADDRPOINTER_REG_13_ & n30472;
  assign n30774 = P1_P3_REIP_REG_13_ & n30490;
  assign n30775 = n30488 & ~n30769;
  assign n30776 = n29097 & n30485;
  assign n30777 = ~n30773 & ~n30774;
  assign n30778 = ~n30775 & n30777;
  assign n30779 = ~n30776 & n30778;
  assign n30780 = ~n30765 & ~n30770;
  assign n30781 = ~n30771 & n30780;
  assign n30782 = ~n30772 & n30781;
  assign n4531 = ~n30779 | ~n30782;
  assign n30784 = P1_P3_PHYADDRPOINTER_REG_13_ & n30761;
  assign n30785 = ~P1_P3_PHYADDRPOINTER_REG_14_ & n30784;
  assign n30786 = P1_P3_PHYADDRPOINTER_REG_14_ & ~n30784;
  assign n30787 = ~n30785 & ~n30786;
  assign n30788 = n30479 & ~n30787;
  assign n30789 = P1_P3_PHYADDRPOINTER_REG_13_ & n30766;
  assign n30790 = ~P1_P3_PHYADDRPOINTER_REG_14_ & n30789;
  assign n30791 = P1_P3_PHYADDRPOINTER_REG_14_ & ~n30789;
  assign n30792 = ~n30790 & ~n30791;
  assign n30793 = n30481 & ~n30792;
  assign n30794 = ~n29168 & n30474;
  assign n30795 = ~n29172 & n30476;
  assign n30796 = P1_P3_PHYADDRPOINTER_REG_14_ & n30472;
  assign n30797 = P1_P3_REIP_REG_14_ & n30490;
  assign n30798 = n30488 & ~n30792;
  assign n30799 = ~n29141 & n30485;
  assign n30800 = ~n30796 & ~n30797;
  assign n30801 = ~n30798 & n30800;
  assign n30802 = ~n30799 & n30801;
  assign n30803 = ~n30788 & ~n30793;
  assign n30804 = ~n30794 & n30803;
  assign n30805 = ~n30795 & n30804;
  assign n4536 = ~n30802 | ~n30805;
  assign n30807 = P1_P3_PHYADDRPOINTER_REG_14_ & n30784;
  assign n30808 = ~P1_P3_PHYADDRPOINTER_REG_15_ & n30807;
  assign n30809 = P1_P3_PHYADDRPOINTER_REG_15_ & ~n30807;
  assign n30810 = ~n30808 & ~n30809;
  assign n30811 = n30479 & ~n30810;
  assign n30812 = P1_P3_PHYADDRPOINTER_REG_14_ & n30789;
  assign n30813 = ~P1_P3_PHYADDRPOINTER_REG_15_ & n30812;
  assign n30814 = P1_P3_PHYADDRPOINTER_REG_15_ & ~n30812;
  assign n30815 = ~n30813 & ~n30814;
  assign n30816 = n30481 & ~n30815;
  assign n30817 = ~n29243 & n30474;
  assign n30818 = n29248 & n30476;
  assign n30819 = P1_P3_PHYADDRPOINTER_REG_15_ & n30472;
  assign n30820 = P1_P3_REIP_REG_15_ & n30490;
  assign n30821 = n30488 & ~n30815;
  assign n30822 = n29217 & n30485;
  assign n30823 = ~n30819 & ~n30820;
  assign n30824 = ~n30821 & n30823;
  assign n30825 = ~n30822 & n30824;
  assign n30826 = ~n30811 & ~n30816;
  assign n30827 = ~n30817 & n30826;
  assign n30828 = ~n30818 & n30827;
  assign n4541 = ~n30825 | ~n30828;
  assign n30830 = P1_P3_PHYADDRPOINTER_REG_15_ & n30807;
  assign n30831 = ~P1_P3_PHYADDRPOINTER_REG_16_ & n30830;
  assign n30832 = P1_P3_PHYADDRPOINTER_REG_16_ & ~n30830;
  assign n30833 = ~n30831 & ~n30832;
  assign n30834 = n30479 & ~n30833;
  assign n30835 = P1_P3_PHYADDRPOINTER_REG_15_ & n30812;
  assign n30836 = ~P1_P3_PHYADDRPOINTER_REG_16_ & n30835;
  assign n30837 = P1_P3_PHYADDRPOINTER_REG_16_ & ~n30835;
  assign n30838 = ~n30836 & ~n30837;
  assign n30839 = n30481 & ~n30838;
  assign n30840 = ~n29279 & n30476;
  assign n30841 = ~n29293 & n30474;
  assign n30842 = P1_P3_PHYADDRPOINTER_REG_16_ & n30472;
  assign n30843 = P1_P3_REIP_REG_16_ & n30490;
  assign n30844 = n30488 & ~n30838;
  assign n30845 = ~n29318 & n30485;
  assign n30846 = ~n30842 & ~n30843;
  assign n30847 = ~n30844 & n30846;
  assign n30848 = ~n30845 & n30847;
  assign n30849 = ~n30834 & ~n30839;
  assign n30850 = ~n30840 & n30849;
  assign n30851 = ~n30841 & n30850;
  assign n4546 = ~n30848 | ~n30851;
  assign n30853 = P1_P3_PHYADDRPOINTER_REG_16_ & n30830;
  assign n30854 = ~P1_P3_PHYADDRPOINTER_REG_17_ & n30853;
  assign n30855 = P1_P3_PHYADDRPOINTER_REG_17_ & ~n30853;
  assign n30856 = ~n30854 & ~n30855;
  assign n30857 = n30479 & ~n30856;
  assign n30858 = P1_P3_PHYADDRPOINTER_REG_16_ & n30835;
  assign n30859 = ~P1_P3_PHYADDRPOINTER_REG_17_ & n30858;
  assign n30860 = P1_P3_PHYADDRPOINTER_REG_17_ & ~n30858;
  assign n30861 = ~n30859 & ~n30860;
  assign n30862 = n30481 & ~n30861;
  assign n30863 = n29343 & n30476;
  assign n30864 = n29395 & n30474;
  assign n30865 = P1_P3_PHYADDRPOINTER_REG_17_ & n30472;
  assign n30866 = P1_P3_REIP_REG_17_ & n30490;
  assign n30867 = n30488 & ~n30861;
  assign n30868 = n29372 & n30485;
  assign n30869 = ~n30865 & ~n30866;
  assign n30870 = ~n30867 & n30869;
  assign n30871 = ~n30868 & n30870;
  assign n30872 = ~n30857 & ~n30862;
  assign n30873 = ~n30863 & n30872;
  assign n30874 = ~n30864 & n30873;
  assign n4551 = ~n30871 | ~n30874;
  assign n30876 = P1_P3_PHYADDRPOINTER_REG_17_ & n30853;
  assign n30877 = ~P1_P3_PHYADDRPOINTER_REG_18_ & n30876;
  assign n30878 = P1_P3_PHYADDRPOINTER_REG_18_ & ~n30876;
  assign n30879 = ~n30877 & ~n30878;
  assign n30880 = n30479 & ~n30879;
  assign n30881 = P1_P3_PHYADDRPOINTER_REG_17_ & n30858;
  assign n30882 = ~P1_P3_PHYADDRPOINTER_REG_18_ & n30881;
  assign n30883 = P1_P3_PHYADDRPOINTER_REG_18_ & ~n30881;
  assign n30884 = ~n30882 & ~n30883;
  assign n30885 = n30481 & ~n30884;
  assign n30886 = ~n29430 & n30476;
  assign n30887 = ~n29443 & n30474;
  assign n30888 = P1_P3_PHYADDRPOINTER_REG_18_ & n30472;
  assign n30889 = P1_P3_REIP_REG_18_ & n30490;
  assign n30890 = n30488 & ~n30884;
  assign n30891 = ~n29468 & n30485;
  assign n30892 = ~n30888 & ~n30889;
  assign n30893 = ~n30890 & n30892;
  assign n30894 = ~n30891 & n30893;
  assign n30895 = ~n30880 & ~n30885;
  assign n30896 = ~n30886 & n30895;
  assign n30897 = ~n30887 & n30896;
  assign n4556 = ~n30894 | ~n30897;
  assign n30899 = P1_P3_PHYADDRPOINTER_REG_18_ & n30876;
  assign n30900 = ~P1_P3_PHYADDRPOINTER_REG_19_ & n30899;
  assign n30901 = P1_P3_PHYADDRPOINTER_REG_19_ & ~n30899;
  assign n30902 = ~n30900 & ~n30901;
  assign n30903 = n30479 & ~n30902;
  assign n30904 = P1_P3_PHYADDRPOINTER_REG_18_ & n30881;
  assign n30905 = ~P1_P3_PHYADDRPOINTER_REG_19_ & n30904;
  assign n30906 = P1_P3_PHYADDRPOINTER_REG_19_ & ~n30904;
  assign n30907 = ~n30905 & ~n30906;
  assign n30908 = n30481 & ~n30907;
  assign n30909 = n29493 & n30476;
  assign n30910 = ~n29544 & n30474;
  assign n30911 = P1_P3_PHYADDRPOINTER_REG_19_ & n30472;
  assign n30912 = P1_P3_REIP_REG_19_ & n30490;
  assign n30913 = n30488 & ~n30907;
  assign n30914 = n29522 & n30485;
  assign n30915 = ~n30911 & ~n30912;
  assign n30916 = ~n30913 & n30915;
  assign n30917 = ~n30914 & n30916;
  assign n30918 = ~n30903 & ~n30908;
  assign n30919 = ~n30909 & n30918;
  assign n30920 = ~n30910 & n30919;
  assign n4561 = ~n30917 | ~n30920;
  assign n30922 = P1_P3_PHYADDRPOINTER_REG_19_ & n30899;
  assign n30923 = ~P1_P3_PHYADDRPOINTER_REG_20_ & n30922;
  assign n30924 = P1_P3_PHYADDRPOINTER_REG_20_ & ~n30922;
  assign n30925 = ~n30923 & ~n30924;
  assign n30926 = n30479 & ~n30925;
  assign n30927 = P1_P3_PHYADDRPOINTER_REG_19_ & n30904;
  assign n30928 = ~P1_P3_PHYADDRPOINTER_REG_20_ & n30927;
  assign n30929 = P1_P3_PHYADDRPOINTER_REG_20_ & ~n30927;
  assign n30930 = ~n30928 & ~n30929;
  assign n30931 = n30481 & ~n30930;
  assign n30932 = n29598 & n30476;
  assign n30933 = P1_P3_PHYADDRPOINTER_REG_20_ & n30472;
  assign n30934 = P1_P3_REIP_REG_20_ & n30490;
  assign n30935 = n30488 & ~n30930;
  assign n30936 = n29622 & n30485;
  assign n30937 = ~n30933 & ~n30934;
  assign n30938 = ~n30935 & n30937;
  assign n30939 = ~n30936 & n30938;
  assign n30940 = n29573 & n30474;
  assign n30941 = ~n30926 & ~n30931;
  assign n30942 = ~n30932 & n30941;
  assign n30943 = n30939 & n30942;
  assign n4566 = n30940 | ~n30943;
  assign n30945 = P1_P3_PHYADDRPOINTER_REG_20_ & n30922;
  assign n30946 = ~P1_P3_PHYADDRPOINTER_REG_21_ & n30945;
  assign n30947 = P1_P3_PHYADDRPOINTER_REG_21_ & ~n30945;
  assign n30948 = ~n30946 & ~n30947;
  assign n30949 = n30479 & ~n30948;
  assign n30950 = P1_P3_PHYADDRPOINTER_REG_20_ & n30927;
  assign n30951 = ~P1_P3_PHYADDRPOINTER_REG_21_ & n30950;
  assign n30952 = P1_P3_PHYADDRPOINTER_REG_21_ & ~n30950;
  assign n30953 = ~n30951 & ~n30952;
  assign n30954 = n30481 & ~n30953;
  assign n30955 = n29670 & n30476;
  assign n30956 = P1_P3_PHYADDRPOINTER_REG_21_ & n30472;
  assign n30957 = P1_P3_REIP_REG_21_ & n30490;
  assign n30958 = n30488 & ~n30953;
  assign n30959 = n29695 & n30485;
  assign n30960 = ~n30956 & ~n30957;
  assign n30961 = ~n30958 & n30960;
  assign n30962 = ~n30959 & n30961;
  assign n30963 = ~n29645 & n30474;
  assign n30964 = ~n30949 & ~n30954;
  assign n30965 = ~n30955 & n30964;
  assign n30966 = n30962 & n30965;
  assign n4571 = n30963 | ~n30966;
  assign n30968 = P1_P3_PHYADDRPOINTER_REG_21_ & n30945;
  assign n30969 = ~P1_P3_PHYADDRPOINTER_REG_22_ & n30968;
  assign n30970 = P1_P3_PHYADDRPOINTER_REG_22_ & ~n30968;
  assign n30971 = ~n30969 & ~n30970;
  assign n30972 = n30479 & ~n30971;
  assign n30973 = P1_P3_PHYADDRPOINTER_REG_21_ & n30950;
  assign n30974 = ~P1_P3_PHYADDRPOINTER_REG_22_ & n30973;
  assign n30975 = P1_P3_PHYADDRPOINTER_REG_22_ & ~n30973;
  assign n30976 = ~n30974 & ~n30975;
  assign n30977 = n30481 & ~n30976;
  assign n30978 = ~n29757 & n30474;
  assign n30979 = ~n29774 & n30476;
  assign n30980 = P1_P3_PHYADDRPOINTER_REG_22_ & n30472;
  assign n30981 = P1_P3_REIP_REG_22_ & n30490;
  assign n30982 = n30488 & ~n30976;
  assign n30983 = ~n29736 & n30485;
  assign n30984 = ~n30980 & ~n30981;
  assign n30985 = ~n30982 & n30984;
  assign n30986 = ~n30983 & n30985;
  assign n30987 = ~n30972 & ~n30977;
  assign n30988 = ~n30978 & n30987;
  assign n30989 = ~n30979 & n30988;
  assign n4576 = ~n30986 | ~n30989;
  assign n30991 = P1_P3_PHYADDRPOINTER_REG_22_ & n30968;
  assign n30992 = ~P1_P3_PHYADDRPOINTER_REG_23_ & n30991;
  assign n30993 = P1_P3_PHYADDRPOINTER_REG_23_ & ~n30991;
  assign n30994 = ~n30992 & ~n30993;
  assign n30995 = n30479 & ~n30994;
  assign n30996 = P1_P3_PHYADDRPOINTER_REG_22_ & n30973;
  assign n30997 = ~P1_P3_PHYADDRPOINTER_REG_23_ & n30996;
  assign n30998 = P1_P3_PHYADDRPOINTER_REG_23_ & ~n30996;
  assign n30999 = ~n30997 & ~n30998;
  assign n31000 = n30481 & ~n30999;
  assign n31001 = ~n29833 & n30474;
  assign n31002 = n29851 & n30476;
  assign n31003 = P1_P3_PHYADDRPOINTER_REG_23_ & n30472;
  assign n31004 = P1_P3_REIP_REG_23_ & n30490;
  assign n31005 = n30488 & ~n30999;
  assign n31006 = n29815 & n30485;
  assign n31007 = ~n31003 & ~n31004;
  assign n31008 = ~n31005 & n31007;
  assign n31009 = ~n31006 & n31008;
  assign n31010 = ~n30995 & ~n31000;
  assign n31011 = ~n31001 & n31010;
  assign n31012 = ~n31002 & n31011;
  assign n4581 = ~n31009 | ~n31012;
  assign n31014 = P1_P3_PHYADDRPOINTER_REG_23_ & n30991;
  assign n31015 = ~P1_P3_PHYADDRPOINTER_REG_24_ & n31014;
  assign n31016 = P1_P3_PHYADDRPOINTER_REG_24_ & ~n31014;
  assign n31017 = ~n31015 & ~n31016;
  assign n31018 = n30479 & ~n31017;
  assign n31019 = ~n29908 & n30474;
  assign n31020 = P1_P3_PHYADDRPOINTER_REG_23_ & n30996;
  assign n31021 = ~P1_P3_PHYADDRPOINTER_REG_24_ & n31020;
  assign n31022 = P1_P3_PHYADDRPOINTER_REG_24_ & ~n31020;
  assign n31023 = ~n31021 & ~n31022;
  assign n31024 = n30481 & ~n31023;
  assign n31025 = ~n29916 & n30476;
  assign n31026 = P1_P3_PHYADDRPOINTER_REG_24_ & n30472;
  assign n31027 = P1_P3_REIP_REG_24_ & n30490;
  assign n31028 = n30488 & ~n31023;
  assign n31029 = ~n29881 & n30485;
  assign n31030 = ~n31026 & ~n31027;
  assign n31031 = ~n31028 & n31030;
  assign n31032 = ~n31029 & n31031;
  assign n31033 = ~n31018 & ~n31019;
  assign n31034 = ~n31024 & n31033;
  assign n31035 = ~n31025 & n31034;
  assign n4586 = ~n31032 | ~n31035;
  assign n31037 = P1_P3_PHYADDRPOINTER_REG_24_ & n31014;
  assign n31038 = ~P1_P3_PHYADDRPOINTER_REG_25_ & n31037;
  assign n31039 = P1_P3_PHYADDRPOINTER_REG_25_ & ~n31037;
  assign n31040 = ~n31038 & ~n31039;
  assign n31041 = n30479 & ~n31040;
  assign n31042 = ~n29987 & n30474;
  assign n31043 = P1_P3_PHYADDRPOINTER_REG_24_ & n31020;
  assign n31044 = ~P1_P3_PHYADDRPOINTER_REG_25_ & n31043;
  assign n31045 = P1_P3_PHYADDRPOINTER_REG_25_ & ~n31043;
  assign n31046 = ~n31044 & ~n31045;
  assign n31047 = n30481 & ~n31046;
  assign n31048 = n29993 & n30476;
  assign n31049 = P1_P3_PHYADDRPOINTER_REG_25_ & n30472;
  assign n31050 = P1_P3_REIP_REG_25_ & n30490;
  assign n31051 = n30488 & ~n31046;
  assign n31052 = n29957 & n30485;
  assign n31053 = ~n31049 & ~n31050;
  assign n31054 = ~n31051 & n31053;
  assign n31055 = ~n31052 & n31054;
  assign n31056 = ~n31041 & ~n31042;
  assign n31057 = ~n31047 & n31056;
  assign n31058 = ~n31048 & n31057;
  assign n4591 = ~n31055 | ~n31058;
  assign n31060 = P1_P3_PHYADDRPOINTER_REG_25_ & n31037;
  assign n31061 = ~P1_P3_PHYADDRPOINTER_REG_26_ & n31060;
  assign n31062 = P1_P3_PHYADDRPOINTER_REG_26_ & ~n31060;
  assign n31063 = ~n31061 & ~n31062;
  assign n31064 = n30479 & ~n31063;
  assign n31065 = n30028 & n30474;
  assign n31066 = P1_P3_PHYADDRPOINTER_REG_25_ & n31043;
  assign n31067 = ~P1_P3_PHYADDRPOINTER_REG_26_ & n31066;
  assign n31068 = P1_P3_PHYADDRPOINTER_REG_26_ & ~n31066;
  assign n31069 = ~n31067 & ~n31068;
  assign n31070 = n30481 & ~n31069;
  assign n31071 = n30032 & n30476;
  assign n31072 = P1_P3_PHYADDRPOINTER_REG_26_ & n30472;
  assign n31073 = n30070 & n30485;
  assign n31074 = n30488 & ~n31069;
  assign n31075 = P1_P3_REIP_REG_26_ & n30490;
  assign n31076 = ~n31072 & ~n31073;
  assign n31077 = ~n31074 & n31076;
  assign n31078 = ~n31075 & n31077;
  assign n31079 = ~n31064 & ~n31065;
  assign n31080 = ~n31070 & n31079;
  assign n31081 = ~n31071 & n31080;
  assign n4596 = ~n31078 | ~n31081;
  assign n31083 = P1_P3_PHYADDRPOINTER_REG_26_ & n31060;
  assign n31084 = ~P1_P3_PHYADDRPOINTER_REG_27_ & n31083;
  assign n31085 = P1_P3_PHYADDRPOINTER_REG_27_ & ~n31083;
  assign n31086 = ~n31084 & ~n31085;
  assign n31087 = n30479 & ~n31086;
  assign n31088 = ~n30099 & n30474;
  assign n31089 = P1_P3_PHYADDRPOINTER_REG_26_ & n31066;
  assign n31090 = ~P1_P3_PHYADDRPOINTER_REG_27_ & n31089;
  assign n31091 = P1_P3_PHYADDRPOINTER_REG_27_ & ~n31089;
  assign n31092 = ~n31090 & ~n31091;
  assign n31093 = n30481 & ~n31092;
  assign n31094 = ~n30103 & n30476;
  assign n31095 = P1_P3_PHYADDRPOINTER_REG_27_ & n30472;
  assign n31096 = ~n30141 & n30485;
  assign n31097 = n30488 & ~n31092;
  assign n31098 = P1_P3_REIP_REG_27_ & n30490;
  assign n31099 = ~n31095 & ~n31096;
  assign n31100 = ~n31097 & n31099;
  assign n31101 = ~n31098 & n31100;
  assign n31102 = ~n31087 & ~n31088;
  assign n31103 = ~n31093 & n31102;
  assign n31104 = ~n31094 & n31103;
  assign n4601 = ~n31101 | ~n31104;
  assign n31106 = n30177 & n30474;
  assign n31107 = n30182 & n30476;
  assign n31108 = P1_P3_PHYADDRPOINTER_REG_27_ & n31083;
  assign n31109 = ~P1_P3_PHYADDRPOINTER_REG_28_ & n31108;
  assign n31110 = P1_P3_PHYADDRPOINTER_REG_28_ & ~n31108;
  assign n31111 = ~n31109 & ~n31110;
  assign n31112 = n30479 & ~n31111;
  assign n31113 = P1_P3_PHYADDRPOINTER_REG_27_ & n31089;
  assign n31114 = ~P1_P3_PHYADDRPOINTER_REG_28_ & n31113;
  assign n31115 = P1_P3_PHYADDRPOINTER_REG_28_ & ~n31113;
  assign n31116 = ~n31114 & ~n31115;
  assign n31117 = n30481 & ~n31116;
  assign n31118 = P1_P3_PHYADDRPOINTER_REG_28_ & n30472;
  assign n31119 = n30221 & n30485;
  assign n31120 = n30488 & ~n31116;
  assign n31121 = P1_P3_REIP_REG_28_ & n30490;
  assign n31122 = ~n31118 & ~n31119;
  assign n31123 = ~n31120 & n31122;
  assign n31124 = ~n31121 & n31123;
  assign n31125 = ~n31106 & ~n31107;
  assign n31126 = ~n31112 & n31125;
  assign n31127 = ~n31117 & n31126;
  assign n4606 = ~n31124 | ~n31127;
  assign n31129 = ~n30250 & n30474;
  assign n31130 = n30254 & n30476;
  assign n31131 = P1_P3_PHYADDRPOINTER_REG_28_ & n31108;
  assign n31132 = ~P1_P3_PHYADDRPOINTER_REG_29_ & n31131;
  assign n31133 = P1_P3_PHYADDRPOINTER_REG_29_ & ~n31131;
  assign n31134 = ~n31132 & ~n31133;
  assign n31135 = n30479 & ~n31134;
  assign n31136 = P1_P3_PHYADDRPOINTER_REG_28_ & n31113;
  assign n31137 = ~P1_P3_PHYADDRPOINTER_REG_29_ & n31136;
  assign n31138 = P1_P3_PHYADDRPOINTER_REG_29_ & ~n31136;
  assign n31139 = ~n31137 & ~n31138;
  assign n31140 = n30481 & ~n31139;
  assign n31141 = P1_P3_PHYADDRPOINTER_REG_29_ & n30472;
  assign n31142 = P1_P3_REIP_REG_29_ & n30490;
  assign n31143 = n30292 & n30485;
  assign n31144 = n30488 & ~n31139;
  assign n31145 = ~n31141 & ~n31142;
  assign n31146 = ~n31143 & n31145;
  assign n31147 = ~n31144 & n31146;
  assign n31148 = ~n31129 & ~n31130;
  assign n31149 = ~n31135 & n31148;
  assign n31150 = ~n31140 & n31149;
  assign n4611 = ~n31147 | ~n31150;
  assign n31152 = ~n30323 & n30474;
  assign n31153 = ~n30327 & n30476;
  assign n31154 = P1_P3_PHYADDRPOINTER_REG_29_ & n31131;
  assign n31155 = ~P1_P3_PHYADDRPOINTER_REG_30_ & n31154;
  assign n31156 = P1_P3_PHYADDRPOINTER_REG_30_ & ~n31154;
  assign n31157 = ~n31155 & ~n31156;
  assign n31158 = n30479 & ~n31157;
  assign n31159 = P1_P3_PHYADDRPOINTER_REG_29_ & n31136;
  assign n31160 = ~P1_P3_PHYADDRPOINTER_REG_30_ & n31159;
  assign n31161 = P1_P3_PHYADDRPOINTER_REG_30_ & ~n31159;
  assign n31162 = ~n31160 & ~n31161;
  assign n31163 = n30481 & ~n31162;
  assign n31164 = P1_P3_PHYADDRPOINTER_REG_30_ & n30472;
  assign n31165 = P1_P3_REIP_REG_30_ & n30490;
  assign n31166 = ~n30365 & n30485;
  assign n31167 = n30488 & ~n31162;
  assign n31168 = ~n31164 & ~n31165;
  assign n31169 = ~n31166 & n31168;
  assign n31170 = ~n31167 & n31169;
  assign n31171 = ~n31152 & ~n31153;
  assign n31172 = ~n31158 & n31171;
  assign n31173 = ~n31163 & n31172;
  assign n4616 = ~n31170 | ~n31173;
  assign n31175 = n30436 & n30474;
  assign n31176 = P1_P3_PHYADDRPOINTER_REG_30_ & n31154;
  assign n31177 = ~P1_P3_PHYADDRPOINTER_REG_31_ & n31176;
  assign n31178 = P1_P3_PHYADDRPOINTER_REG_31_ & ~n31176;
  assign n31179 = ~n31177 & ~n31178;
  assign n31180 = n30479 & ~n31179;
  assign n31181 = ~n30441 & n30476;
  assign n31182 = P1_P3_PHYADDRPOINTER_REG_30_ & n31159;
  assign n31183 = ~P1_P3_PHYADDRPOINTER_REG_31_ & n31182;
  assign n31184 = P1_P3_PHYADDRPOINTER_REG_31_ & ~n31182;
  assign n31185 = ~n31183 & ~n31184;
  assign n31186 = n30481 & ~n31185;
  assign n31187 = P1_P3_PHYADDRPOINTER_REG_31_ & n30472;
  assign n31188 = P1_P3_REIP_REG_31_ & n30490;
  assign n31189 = ~n30389 & n30485;
  assign n31190 = n30488 & ~n31185;
  assign n31191 = ~n31187 & ~n31188;
  assign n31192 = ~n31189 & n31191;
  assign n31193 = ~n31190 & n31192;
  assign n31194 = ~n31175 & ~n31180;
  assign n31195 = ~n31181 & n31194;
  assign n31196 = ~n31186 & n31195;
  assign n4621 = ~n31193 | ~n31196;
  assign n31198 = ~n25267 & n25723;
  assign n31199 = n25692 & n31198;
  assign n31200 = ~n25879 & ~n31199;
  assign n31201 = n25994 & ~n31200;
  assign n31202 = ~n25608 & n31201;
  assign n31203 = P1_BUF2_REG_15_ & n31202;
  assign n31204 = n25608 & n31201;
  assign n31205 = P1_P3_EAX_REG_15_ & n31204;
  assign n31206 = P1_P3_LWORD_REG_15_ & ~n31201;
  assign n31207 = ~n31203 & ~n31205;
  assign n4626 = n31206 | ~n31207;
  assign n31209 = P1_BUF2_REG_14_ & n31202;
  assign n31210 = P1_P3_EAX_REG_14_ & n31204;
  assign n31211 = P1_P3_LWORD_REG_14_ & ~n31201;
  assign n31212 = ~n31209 & ~n31210;
  assign n4631 = n31211 | ~n31212;
  assign n31214 = P1_BUF2_REG_13_ & n31202;
  assign n31215 = P1_P3_EAX_REG_13_ & n31204;
  assign n31216 = P1_P3_LWORD_REG_13_ & ~n31201;
  assign n31217 = ~n31214 & ~n31215;
  assign n4636 = n31216 | ~n31217;
  assign n31219 = P1_BUF2_REG_12_ & n31202;
  assign n31220 = P1_P3_EAX_REG_12_ & n31204;
  assign n31221 = P1_P3_LWORD_REG_12_ & ~n31201;
  assign n31222 = ~n31219 & ~n31220;
  assign n4641 = n31221 | ~n31222;
  assign n31224 = P1_BUF2_REG_11_ & n31202;
  assign n31225 = P1_P3_EAX_REG_11_ & n31204;
  assign n31226 = P1_P3_LWORD_REG_11_ & ~n31201;
  assign n31227 = ~n31224 & ~n31225;
  assign n4646 = n31226 | ~n31227;
  assign n31229 = P1_BUF2_REG_10_ & n31202;
  assign n31230 = P1_P3_EAX_REG_10_ & n31204;
  assign n31231 = P1_P3_LWORD_REG_10_ & ~n31201;
  assign n31232 = ~n31229 & ~n31230;
  assign n4651 = n31231 | ~n31232;
  assign n31234 = P1_BUF2_REG_9_ & n31202;
  assign n31235 = P1_P3_EAX_REG_9_ & n31204;
  assign n31236 = P1_P3_LWORD_REG_9_ & ~n31201;
  assign n31237 = ~n31234 & ~n31235;
  assign n4656 = n31236 | ~n31237;
  assign n31239 = P1_BUF2_REG_8_ & n31202;
  assign n31240 = P1_P3_EAX_REG_8_ & n31204;
  assign n31241 = P1_P3_LWORD_REG_8_ & ~n31201;
  assign n31242 = ~n31239 & ~n31240;
  assign n4661 = n31241 | ~n31242;
  assign n31244 = P1_BUF2_REG_7_ & n31202;
  assign n31245 = P1_P3_EAX_REG_7_ & n31204;
  assign n31246 = P1_P3_LWORD_REG_7_ & ~n31201;
  assign n31247 = ~n31244 & ~n31245;
  assign n4666 = n31246 | ~n31247;
  assign n31249 = P1_BUF2_REG_6_ & n31202;
  assign n31250 = P1_P3_EAX_REG_6_ & n31204;
  assign n31251 = P1_P3_LWORD_REG_6_ & ~n31201;
  assign n31252 = ~n31249 & ~n31250;
  assign n4671 = n31251 | ~n31252;
  assign n31254 = P1_BUF2_REG_5_ & n31202;
  assign n31255 = P1_P3_EAX_REG_5_ & n31204;
  assign n31256 = P1_P3_LWORD_REG_5_ & ~n31201;
  assign n31257 = ~n31254 & ~n31255;
  assign n4676 = n31256 | ~n31257;
  assign n31259 = P1_BUF2_REG_4_ & n31202;
  assign n31260 = P1_P3_EAX_REG_4_ & n31204;
  assign n31261 = P1_P3_LWORD_REG_4_ & ~n31201;
  assign n31262 = ~n31259 & ~n31260;
  assign n4681 = n31261 | ~n31262;
  assign n31264 = P1_BUF2_REG_3_ & n31202;
  assign n31265 = P1_P3_EAX_REG_3_ & n31204;
  assign n31266 = P1_P3_LWORD_REG_3_ & ~n31201;
  assign n31267 = ~n31264 & ~n31265;
  assign n4686 = n31266 | ~n31267;
  assign n31269 = P1_BUF2_REG_2_ & n31202;
  assign n31270 = P1_P3_EAX_REG_2_ & n31204;
  assign n31271 = P1_P3_LWORD_REG_2_ & ~n31201;
  assign n31272 = ~n31269 & ~n31270;
  assign n4691 = n31271 | ~n31272;
  assign n31274 = P1_BUF2_REG_1_ & n31202;
  assign n31275 = P1_P3_EAX_REG_1_ & n31204;
  assign n31276 = P1_P3_LWORD_REG_1_ & ~n31201;
  assign n31277 = ~n31274 & ~n31275;
  assign n4696 = n31276 | ~n31277;
  assign n31279 = P1_BUF2_REG_0_ & n31202;
  assign n31280 = P1_P3_EAX_REG_0_ & n31204;
  assign n31281 = P1_P3_LWORD_REG_0_ & ~n31201;
  assign n31282 = ~n31279 & ~n31280;
  assign n4701 = n31281 | ~n31282;
  assign n31284 = P1_P3_EAX_REG_30_ & n31204;
  assign n31285 = P1_P3_UWORD_REG_14_ & ~n31201;
  assign n31286 = ~n31209 & ~n31284;
  assign n4706 = n31285 | ~n31286;
  assign n31288 = P1_P3_EAX_REG_29_ & n31204;
  assign n31289 = P1_P3_UWORD_REG_13_ & ~n31201;
  assign n31290 = ~n31214 & ~n31288;
  assign n4711 = n31289 | ~n31290;
  assign n31292 = P1_P3_EAX_REG_28_ & n31204;
  assign n31293 = P1_P3_UWORD_REG_12_ & ~n31201;
  assign n31294 = ~n31219 & ~n31292;
  assign n4716 = n31293 | ~n31294;
  assign n31296 = P1_P3_EAX_REG_27_ & n31204;
  assign n31297 = P1_P3_UWORD_REG_11_ & ~n31201;
  assign n31298 = ~n31224 & ~n31296;
  assign n4721 = n31297 | ~n31298;
  assign n31300 = P1_P3_EAX_REG_26_ & n31204;
  assign n31301 = P1_P3_UWORD_REG_10_ & ~n31201;
  assign n31302 = ~n31229 & ~n31300;
  assign n4726 = n31301 | ~n31302;
  assign n31304 = P1_P3_EAX_REG_25_ & n31204;
  assign n31305 = P1_P3_UWORD_REG_9_ & ~n31201;
  assign n31306 = ~n31234 & ~n31304;
  assign n4731 = n31305 | ~n31306;
  assign n31308 = P1_P3_EAX_REG_24_ & n31204;
  assign n31309 = P1_P3_UWORD_REG_8_ & ~n31201;
  assign n31310 = ~n31239 & ~n31308;
  assign n4736 = n31309 | ~n31310;
  assign n31312 = P1_P3_EAX_REG_23_ & n31204;
  assign n31313 = P1_P3_UWORD_REG_7_ & ~n31201;
  assign n31314 = ~n31244 & ~n31312;
  assign n4741 = n31313 | ~n31314;
  assign n31316 = P1_P3_EAX_REG_22_ & n31204;
  assign n31317 = P1_P3_UWORD_REG_6_ & ~n31201;
  assign n31318 = ~n31249 & ~n31316;
  assign n4746 = n31317 | ~n31318;
  assign n31320 = P1_P3_EAX_REG_21_ & n31204;
  assign n31321 = P1_P3_UWORD_REG_5_ & ~n31201;
  assign n31322 = ~n31254 & ~n31320;
  assign n4751 = n31321 | ~n31322;
  assign n31324 = P1_P3_EAX_REG_20_ & n31204;
  assign n31325 = P1_P3_UWORD_REG_4_ & ~n31201;
  assign n31326 = ~n31259 & ~n31324;
  assign n4756 = n31325 | ~n31326;
  assign n31328 = P1_P3_EAX_REG_19_ & n31204;
  assign n31329 = P1_P3_UWORD_REG_3_ & ~n31201;
  assign n31330 = ~n31264 & ~n31328;
  assign n4761 = n31329 | ~n31330;
  assign n31332 = P1_P3_EAX_REG_18_ & n31204;
  assign n31333 = P1_P3_UWORD_REG_2_ & ~n31201;
  assign n31334 = ~n31269 & ~n31332;
  assign n4766 = n31333 | ~n31334;
  assign n31336 = P1_P3_EAX_REG_17_ & n31204;
  assign n31337 = P1_P3_UWORD_REG_1_ & ~n31201;
  assign n31338 = ~n31274 & ~n31336;
  assign n4771 = n31337 | ~n31338;
  assign n31340 = P1_P3_EAX_REG_16_ & n31204;
  assign n31341 = P1_P3_UWORD_REG_0_ & ~n31201;
  assign n31342 = ~n31279 & ~n31340;
  assign n4776 = n31341 | ~n31342;
  assign n31344 = ~P1_P3_STATE2_REG_0_ & n25352;
  assign n31345 = n25358 & n25994;
  assign n31346 = ~n25880 & n31345;
  assign n31347 = ~n31344 & ~n31346;
  assign n31348 = P1_P3_STATE2_REG_0_ & ~n31347;
  assign n31349 = P1_P3_EAX_REG_0_ & n31348;
  assign n31350 = ~P1_P3_STATE2_REG_0_ & ~n31347;
  assign n31351 = P1_P3_LWORD_REG_0_ & n31350;
  assign n31352 = P1_P3_DATAO_REG_0_ & n31347;
  assign n31353 = ~n31349 & ~n31351;
  assign n4781 = n31352 | ~n31353;
  assign n31355 = P1_P3_EAX_REG_1_ & n31348;
  assign n31356 = P1_P3_LWORD_REG_1_ & n31350;
  assign n31357 = P1_P3_DATAO_REG_1_ & n31347;
  assign n31358 = ~n31355 & ~n31356;
  assign n4786 = n31357 | ~n31358;
  assign n31360 = P1_P3_EAX_REG_2_ & n31348;
  assign n31361 = P1_P3_LWORD_REG_2_ & n31350;
  assign n31362 = P1_P3_DATAO_REG_2_ & n31347;
  assign n31363 = ~n31360 & ~n31361;
  assign n4791 = n31362 | ~n31363;
  assign n31365 = P1_P3_EAX_REG_3_ & n31348;
  assign n31366 = P1_P3_LWORD_REG_3_ & n31350;
  assign n31367 = P1_P3_DATAO_REG_3_ & n31347;
  assign n31368 = ~n31365 & ~n31366;
  assign n4796 = n31367 | ~n31368;
  assign n31370 = P1_P3_EAX_REG_4_ & n31348;
  assign n31371 = P1_P3_LWORD_REG_4_ & n31350;
  assign n31372 = P1_P3_DATAO_REG_4_ & n31347;
  assign n31373 = ~n31370 & ~n31371;
  assign n4801 = n31372 | ~n31373;
  assign n31375 = P1_P3_EAX_REG_5_ & n31348;
  assign n31376 = P1_P3_LWORD_REG_5_ & n31350;
  assign n31377 = P1_P3_DATAO_REG_5_ & n31347;
  assign n31378 = ~n31375 & ~n31376;
  assign n4806 = n31377 | ~n31378;
  assign n31380 = P1_P3_EAX_REG_6_ & n31348;
  assign n31381 = P1_P3_LWORD_REG_6_ & n31350;
  assign n31382 = P1_P3_DATAO_REG_6_ & n31347;
  assign n31383 = ~n31380 & ~n31381;
  assign n4811 = n31382 | ~n31383;
  assign n31385 = P1_P3_EAX_REG_7_ & n31348;
  assign n31386 = P1_P3_LWORD_REG_7_ & n31350;
  assign n31387 = P1_P3_DATAO_REG_7_ & n31347;
  assign n31388 = ~n31385 & ~n31386;
  assign n4816 = n31387 | ~n31388;
  assign n31390 = P1_P3_EAX_REG_8_ & n31348;
  assign n31391 = P1_P3_LWORD_REG_8_ & n31350;
  assign n31392 = P1_P3_DATAO_REG_8_ & n31347;
  assign n31393 = ~n31390 & ~n31391;
  assign n4821 = n31392 | ~n31393;
  assign n31395 = P1_P3_EAX_REG_9_ & n31348;
  assign n31396 = P1_P3_LWORD_REG_9_ & n31350;
  assign n31397 = P1_P3_DATAO_REG_9_ & n31347;
  assign n31398 = ~n31395 & ~n31396;
  assign n4826 = n31397 | ~n31398;
  assign n31400 = P1_P3_EAX_REG_10_ & n31348;
  assign n31401 = P1_P3_LWORD_REG_10_ & n31350;
  assign n31402 = P1_P3_DATAO_REG_10_ & n31347;
  assign n31403 = ~n31400 & ~n31401;
  assign n4831 = n31402 | ~n31403;
  assign n31405 = P1_P3_EAX_REG_11_ & n31348;
  assign n31406 = P1_P3_LWORD_REG_11_ & n31350;
  assign n31407 = P1_P3_DATAO_REG_11_ & n31347;
  assign n31408 = ~n31405 & ~n31406;
  assign n4836 = n31407 | ~n31408;
  assign n31410 = P1_P3_EAX_REG_12_ & n31348;
  assign n31411 = P1_P3_LWORD_REG_12_ & n31350;
  assign n31412 = P1_P3_DATAO_REG_12_ & n31347;
  assign n31413 = ~n31410 & ~n31411;
  assign n4841 = n31412 | ~n31413;
  assign n31415 = P1_P3_EAX_REG_13_ & n31348;
  assign n31416 = P1_P3_LWORD_REG_13_ & n31350;
  assign n31417 = P1_P3_DATAO_REG_13_ & n31347;
  assign n31418 = ~n31415 & ~n31416;
  assign n4846 = n31417 | ~n31418;
  assign n31420 = P1_P3_EAX_REG_14_ & n31348;
  assign n31421 = P1_P3_LWORD_REG_14_ & n31350;
  assign n31422 = P1_P3_DATAO_REG_14_ & n31347;
  assign n31423 = ~n31420 & ~n31421;
  assign n4851 = n31422 | ~n31423;
  assign n31425 = P1_P3_EAX_REG_15_ & n31348;
  assign n31426 = P1_P3_LWORD_REG_15_ & n31350;
  assign n31427 = P1_P3_DATAO_REG_15_ & n31347;
  assign n31428 = ~n31425 & ~n31426;
  assign n4856 = n31427 | ~n31428;
  assign n31430 = P1_P3_UWORD_REG_0_ & n31350;
  assign n31431 = P1_P3_DATAO_REG_16_ & n31347;
  assign n31432 = ~n31430 & ~n31431;
  assign n31433 = ~n25639 & n31348;
  assign n31434 = P1_P3_EAX_REG_16_ & n31433;
  assign n4861 = ~n31432 | n31434;
  assign n31436 = P1_P3_UWORD_REG_1_ & n31350;
  assign n31437 = P1_P3_DATAO_REG_17_ & n31347;
  assign n31438 = ~n31436 & ~n31437;
  assign n31439 = P1_P3_EAX_REG_17_ & n31433;
  assign n4866 = ~n31438 | n31439;
  assign n31441 = P1_P3_UWORD_REG_2_ & n31350;
  assign n31442 = P1_P3_DATAO_REG_18_ & n31347;
  assign n31443 = ~n31441 & ~n31442;
  assign n31444 = P1_P3_EAX_REG_18_ & n31433;
  assign n4871 = ~n31443 | n31444;
  assign n31446 = P1_P3_UWORD_REG_3_ & n31350;
  assign n31447 = P1_P3_DATAO_REG_19_ & n31347;
  assign n31448 = ~n31446 & ~n31447;
  assign n31449 = P1_P3_EAX_REG_19_ & n31433;
  assign n4876 = ~n31448 | n31449;
  assign n31451 = P1_P3_UWORD_REG_4_ & n31350;
  assign n31452 = P1_P3_DATAO_REG_20_ & n31347;
  assign n31453 = ~n31451 & ~n31452;
  assign n31454 = P1_P3_EAX_REG_20_ & n31433;
  assign n4881 = ~n31453 | n31454;
  assign n31456 = P1_P3_UWORD_REG_5_ & n31350;
  assign n31457 = P1_P3_DATAO_REG_21_ & n31347;
  assign n31458 = ~n31456 & ~n31457;
  assign n31459 = P1_P3_EAX_REG_21_ & n31433;
  assign n4886 = ~n31458 | n31459;
  assign n31461 = P1_P3_UWORD_REG_6_ & n31350;
  assign n31462 = P1_P3_DATAO_REG_22_ & n31347;
  assign n31463 = ~n31461 & ~n31462;
  assign n31464 = P1_P3_EAX_REG_22_ & n31433;
  assign n4891 = ~n31463 | n31464;
  assign n31466 = P1_P3_UWORD_REG_7_ & n31350;
  assign n31467 = P1_P3_DATAO_REG_23_ & n31347;
  assign n31468 = ~n31466 & ~n31467;
  assign n31469 = P1_P3_EAX_REG_23_ & n31433;
  assign n4896 = ~n31468 | n31469;
  assign n31471 = P1_P3_UWORD_REG_8_ & n31350;
  assign n31472 = P1_P3_DATAO_REG_24_ & n31347;
  assign n31473 = ~n31471 & ~n31472;
  assign n31474 = P1_P3_EAX_REG_24_ & n31433;
  assign n4901 = ~n31473 | n31474;
  assign n31476 = P1_P3_UWORD_REG_9_ & n31350;
  assign n31477 = P1_P3_DATAO_REG_25_ & n31347;
  assign n31478 = ~n31476 & ~n31477;
  assign n31479 = P1_P3_EAX_REG_25_ & n31433;
  assign n4906 = ~n31478 | n31479;
  assign n31481 = P1_P3_UWORD_REG_10_ & n31350;
  assign n31482 = P1_P3_DATAO_REG_26_ & n31347;
  assign n31483 = ~n31481 & ~n31482;
  assign n31484 = P1_P3_EAX_REG_26_ & n31433;
  assign n4911 = ~n31483 | n31484;
  assign n31486 = P1_P3_UWORD_REG_11_ & n31350;
  assign n31487 = P1_P3_DATAO_REG_27_ & n31347;
  assign n31488 = ~n31486 & ~n31487;
  assign n31489 = P1_P3_EAX_REG_27_ & n31433;
  assign n4916 = ~n31488 | n31489;
  assign n31491 = P1_P3_UWORD_REG_12_ & n31350;
  assign n31492 = P1_P3_DATAO_REG_28_ & n31347;
  assign n31493 = ~n31491 & ~n31492;
  assign n31494 = P1_P3_EAX_REG_28_ & n31433;
  assign n4921 = ~n31493 | n31494;
  assign n31496 = P1_P3_UWORD_REG_13_ & n31350;
  assign n31497 = P1_P3_DATAO_REG_29_ & n31347;
  assign n31498 = ~n31496 & ~n31497;
  assign n31499 = P1_P3_EAX_REG_29_ & n31433;
  assign n4926 = ~n31498 | n31499;
  assign n31501 = P1_P3_UWORD_REG_14_ & n31350;
  assign n31502 = P1_P3_DATAO_REG_30_ & n31347;
  assign n31503 = ~n31501 & ~n31502;
  assign n31504 = P1_P3_EAX_REG_30_ & n31433;
  assign n4931 = ~n31503 | n31504;
  assign n4936 = P1_P3_DATAO_REG_31_ & n31347;
  assign n31507 = n25874 & ~n25938;
  assign n31508 = n25994 & ~n31507;
  assign n31509 = n25728 & n31508;
  assign n31510 = ~n27704 & n31509;
  assign n31511 = ~n25511 & n31508;
  assign n31512 = ~n25728 & n31511;
  assign n31513 = P1_BUF2_REG_0_ & n31512;
  assign n31514 = P1_P3_EAX_REG_0_ & ~n31508;
  assign n31515 = n25511 & n31508;
  assign n31516 = ~P1_P3_EAX_REG_0_ & n31515;
  assign n31517 = ~n31514 & ~n31516;
  assign n31518 = ~n31510 & ~n31513;
  assign n4941 = ~n31517 | ~n31518;
  assign n31520 = ~n27822 & n31509;
  assign n31521 = P1_BUF2_REG_1_ & n31512;
  assign n31522 = P1_P3_EAX_REG_1_ & ~n31508;
  assign n31523 = ~P1_P3_EAX_REG_0_ & P1_P3_EAX_REG_1_;
  assign n31524 = P1_P3_EAX_REG_0_ & ~P1_P3_EAX_REG_1_;
  assign n31525 = ~n31523 & ~n31524;
  assign n31526 = n31515 & ~n31525;
  assign n31527 = ~n31522 & ~n31526;
  assign n31528 = ~n31520 & ~n31521;
  assign n4946 = ~n31527 | ~n31528;
  assign n31530 = ~n27933 & n31509;
  assign n31531 = P1_BUF2_REG_2_ & n31512;
  assign n31532 = P1_P3_EAX_REG_2_ & ~n31508;
  assign n31533 = P1_P3_EAX_REG_0_ & P1_P3_EAX_REG_1_;
  assign n31534 = ~P1_P3_EAX_REG_2_ & n31533;
  assign n31535 = P1_P3_EAX_REG_2_ & ~n31533;
  assign n31536 = ~n31534 & ~n31535;
  assign n31537 = n31515 & ~n31536;
  assign n31538 = ~n31532 & ~n31537;
  assign n31539 = ~n31530 & ~n31531;
  assign n4951 = ~n31538 | ~n31539;
  assign n31541 = ~n28058 & n31509;
  assign n31542 = P1_BUF2_REG_3_ & n31512;
  assign n31543 = P1_P3_EAX_REG_3_ & ~n31508;
  assign n31544 = P1_P3_EAX_REG_0_ & P1_P3_EAX_REG_2_;
  assign n31545 = P1_P3_EAX_REG_1_ & n31544;
  assign n31546 = P1_P3_EAX_REG_3_ & ~n31545;
  assign n31547 = ~P1_P3_EAX_REG_3_ & n31545;
  assign n31548 = ~n31546 & ~n31547;
  assign n31549 = n31515 & ~n31548;
  assign n31550 = ~n31543 & ~n31549;
  assign n31551 = ~n31541 & ~n31542;
  assign n4956 = ~n31550 | ~n31551;
  assign n31553 = ~n28185 & n31509;
  assign n31554 = P1_BUF2_REG_4_ & n31512;
  assign n31555 = P1_P3_EAX_REG_4_ & ~n31508;
  assign n31556 = P1_P3_EAX_REG_3_ & n31545;
  assign n31557 = ~P1_P3_EAX_REG_4_ & n31556;
  assign n31558 = P1_P3_EAX_REG_4_ & ~n31556;
  assign n31559 = ~n31557 & ~n31558;
  assign n31560 = n31515 & ~n31559;
  assign n31561 = ~n31555 & ~n31560;
  assign n31562 = ~n31553 & ~n31554;
  assign n4961 = ~n31561 | ~n31562;
  assign n31564 = ~n28326 & n31509;
  assign n31565 = P1_BUF2_REG_5_ & n31512;
  assign n31566 = P1_P3_EAX_REG_5_ & ~n31508;
  assign n31567 = P1_P3_EAX_REG_3_ & P1_P3_EAX_REG_4_;
  assign n31568 = n31545 & n31567;
  assign n31569 = P1_P3_EAX_REG_5_ & ~n31568;
  assign n31570 = ~P1_P3_EAX_REG_5_ & n31568;
  assign n31571 = ~n31569 & ~n31570;
  assign n31572 = n31515 & ~n31571;
  assign n31573 = ~n31566 & ~n31572;
  assign n31574 = ~n31564 & ~n31565;
  assign n4966 = ~n31573 | ~n31574;
  assign n31576 = ~n28458 & n31509;
  assign n31577 = P1_BUF2_REG_6_ & n31512;
  assign n31578 = P1_P3_EAX_REG_6_ & ~n31508;
  assign n31579 = P1_P3_EAX_REG_5_ & n31568;
  assign n31580 = ~P1_P3_EAX_REG_6_ & n31579;
  assign n31581 = P1_P3_EAX_REG_6_ & ~n31579;
  assign n31582 = ~n31580 & ~n31581;
  assign n31583 = n31515 & ~n31582;
  assign n31584 = ~n31578 & ~n31583;
  assign n31585 = ~n31576 & ~n31577;
  assign n4971 = ~n31584 | ~n31585;
  assign n31587 = ~n27738 & n31509;
  assign n31588 = P1_BUF2_REG_7_ & n31512;
  assign n31589 = P1_P3_EAX_REG_7_ & ~n31508;
  assign n31590 = P1_P3_EAX_REG_5_ & P1_P3_EAX_REG_6_;
  assign n31591 = n31568 & n31590;
  assign n31592 = P1_P3_EAX_REG_7_ & ~n31591;
  assign n31593 = ~P1_P3_EAX_REG_7_ & n31591;
  assign n31594 = ~n31592 & ~n31593;
  assign n31595 = n31515 & ~n31594;
  assign n31596 = ~n31589 & ~n31595;
  assign n31597 = ~n31587 & ~n31588;
  assign n4976 = ~n31596 | ~n31597;
  assign n31599 = ~n25888 & ~n25895;
  assign n31600 = ~n25839 & ~n31599;
  assign n31601 = n25369 & n31600;
  assign n31602 = P1_P3_INSTQUEUE_REG_15__0_ & n31601;
  assign n31603 = n25373 & n31600;
  assign n31604 = P1_P3_INSTQUEUE_REG_14__0_ & n31603;
  assign n31605 = n25360 & n31600;
  assign n31606 = P1_P3_INSTQUEUE_REG_13__0_ & n31605;
  assign n31607 = n25364 & n31600;
  assign n31608 = P1_P3_INSTQUEUE_REG_12__0_ & n31607;
  assign n31609 = ~n31602 & ~n31604;
  assign n31610 = ~n31606 & n31609;
  assign n31611 = ~n31608 & n31610;
  assign n31612 = n25839 & ~n31599;
  assign n31613 = n25369 & n31612;
  assign n31614 = P1_P3_INSTQUEUE_REG_11__0_ & n31613;
  assign n31615 = n25373 & n31612;
  assign n31616 = P1_P3_INSTQUEUE_REG_10__0_ & n31615;
  assign n31617 = n25360 & n31612;
  assign n31618 = P1_P3_INSTQUEUE_REG_9__0_ & n31617;
  assign n31619 = n25364 & n31612;
  assign n31620 = P1_P3_INSTQUEUE_REG_8__0_ & n31619;
  assign n31621 = ~n31614 & ~n31616;
  assign n31622 = ~n31618 & n31621;
  assign n31623 = ~n31620 & n31622;
  assign n31624 = ~n25839 & n31599;
  assign n31625 = n25369 & n31624;
  assign n31626 = P1_P3_INSTQUEUE_REG_7__0_ & n31625;
  assign n31627 = n25373 & n31624;
  assign n31628 = P1_P3_INSTQUEUE_REG_6__0_ & n31627;
  assign n31629 = n25360 & n31624;
  assign n31630 = P1_P3_INSTQUEUE_REG_5__0_ & n31629;
  assign n31631 = n25364 & n31624;
  assign n31632 = P1_P3_INSTQUEUE_REG_4__0_ & n31631;
  assign n31633 = ~n31626 & ~n31628;
  assign n31634 = ~n31630 & n31633;
  assign n31635 = ~n31632 & n31634;
  assign n31636 = n25839 & n31599;
  assign n31637 = n25369 & n31636;
  assign n31638 = P1_P3_INSTQUEUE_REG_3__0_ & n31637;
  assign n31639 = n25373 & n31636;
  assign n31640 = P1_P3_INSTQUEUE_REG_2__0_ & n31639;
  assign n31641 = n25360 & n31636;
  assign n31642 = P1_P3_INSTQUEUE_REG_1__0_ & n31641;
  assign n31643 = n25364 & n31636;
  assign n31644 = P1_P3_INSTQUEUE_REG_0__0_ & n31643;
  assign n31645 = ~n31638 & ~n31640;
  assign n31646 = ~n31642 & n31645;
  assign n31647 = ~n31644 & n31646;
  assign n31648 = n31611 & n31623;
  assign n31649 = n31635 & n31648;
  assign n31650 = n31647 & n31649;
  assign n31651 = n31509 & ~n31650;
  assign n31652 = P1_BUF2_REG_8_ & n31512;
  assign n31653 = P1_P3_EAX_REG_8_ & ~n31508;
  assign n31654 = P1_P3_EAX_REG_7_ & n31591;
  assign n31655 = ~P1_P3_EAX_REG_8_ & n31654;
  assign n31656 = P1_P3_EAX_REG_8_ & ~n31654;
  assign n31657 = ~n31655 & ~n31656;
  assign n31658 = n31515 & ~n31657;
  assign n31659 = ~n31653 & ~n31658;
  assign n31660 = ~n31651 & ~n31652;
  assign n4981 = ~n31659 | ~n31660;
  assign n31662 = P1_P3_INSTQUEUE_REG_15__1_ & n31601;
  assign n31663 = P1_P3_INSTQUEUE_REG_14__1_ & n31603;
  assign n31664 = P1_P3_INSTQUEUE_REG_13__1_ & n31605;
  assign n31665 = P1_P3_INSTQUEUE_REG_12__1_ & n31607;
  assign n31666 = ~n31662 & ~n31663;
  assign n31667 = ~n31664 & n31666;
  assign n31668 = ~n31665 & n31667;
  assign n31669 = P1_P3_INSTQUEUE_REG_11__1_ & n31613;
  assign n31670 = P1_P3_INSTQUEUE_REG_10__1_ & n31615;
  assign n31671 = P1_P3_INSTQUEUE_REG_9__1_ & n31617;
  assign n31672 = P1_P3_INSTQUEUE_REG_8__1_ & n31619;
  assign n31673 = ~n31669 & ~n31670;
  assign n31674 = ~n31671 & n31673;
  assign n31675 = ~n31672 & n31674;
  assign n31676 = P1_P3_INSTQUEUE_REG_7__1_ & n31625;
  assign n31677 = P1_P3_INSTQUEUE_REG_6__1_ & n31627;
  assign n31678 = P1_P3_INSTQUEUE_REG_5__1_ & n31629;
  assign n31679 = P1_P3_INSTQUEUE_REG_4__1_ & n31631;
  assign n31680 = ~n31676 & ~n31677;
  assign n31681 = ~n31678 & n31680;
  assign n31682 = ~n31679 & n31681;
  assign n31683 = P1_P3_INSTQUEUE_REG_3__1_ & n31637;
  assign n31684 = P1_P3_INSTQUEUE_REG_2__1_ & n31639;
  assign n31685 = P1_P3_INSTQUEUE_REG_1__1_ & n31641;
  assign n31686 = P1_P3_INSTQUEUE_REG_0__1_ & n31643;
  assign n31687 = ~n31683 & ~n31684;
  assign n31688 = ~n31685 & n31687;
  assign n31689 = ~n31686 & n31688;
  assign n31690 = n31668 & n31675;
  assign n31691 = n31682 & n31690;
  assign n31692 = n31689 & n31691;
  assign n31693 = n31509 & ~n31692;
  assign n31694 = P1_BUF2_REG_9_ & n31512;
  assign n31695 = P1_P3_EAX_REG_9_ & ~n31508;
  assign n31696 = P1_P3_EAX_REG_7_ & P1_P3_EAX_REG_8_;
  assign n31697 = n31591 & n31696;
  assign n31698 = P1_P3_EAX_REG_9_ & ~n31697;
  assign n31699 = ~P1_P3_EAX_REG_9_ & n31697;
  assign n31700 = ~n31698 & ~n31699;
  assign n31701 = n31515 & ~n31700;
  assign n31702 = ~n31695 & ~n31701;
  assign n31703 = ~n31693 & ~n31694;
  assign n4986 = ~n31702 | ~n31703;
  assign n31705 = P1_P3_INSTQUEUE_REG_15__2_ & n31601;
  assign n31706 = P1_P3_INSTQUEUE_REG_14__2_ & n31603;
  assign n31707 = P1_P3_INSTQUEUE_REG_13__2_ & n31605;
  assign n31708 = P1_P3_INSTQUEUE_REG_12__2_ & n31607;
  assign n31709 = ~n31705 & ~n31706;
  assign n31710 = ~n31707 & n31709;
  assign n31711 = ~n31708 & n31710;
  assign n31712 = P1_P3_INSTQUEUE_REG_11__2_ & n31613;
  assign n31713 = P1_P3_INSTQUEUE_REG_10__2_ & n31615;
  assign n31714 = P1_P3_INSTQUEUE_REG_9__2_ & n31617;
  assign n31715 = P1_P3_INSTQUEUE_REG_8__2_ & n31619;
  assign n31716 = ~n31712 & ~n31713;
  assign n31717 = ~n31714 & n31716;
  assign n31718 = ~n31715 & n31717;
  assign n31719 = P1_P3_INSTQUEUE_REG_7__2_ & n31625;
  assign n31720 = P1_P3_INSTQUEUE_REG_6__2_ & n31627;
  assign n31721 = P1_P3_INSTQUEUE_REG_5__2_ & n31629;
  assign n31722 = P1_P3_INSTQUEUE_REG_4__2_ & n31631;
  assign n31723 = ~n31719 & ~n31720;
  assign n31724 = ~n31721 & n31723;
  assign n31725 = ~n31722 & n31724;
  assign n31726 = P1_P3_INSTQUEUE_REG_3__2_ & n31637;
  assign n31727 = P1_P3_INSTQUEUE_REG_2__2_ & n31639;
  assign n31728 = P1_P3_INSTQUEUE_REG_1__2_ & n31641;
  assign n31729 = P1_P3_INSTQUEUE_REG_0__2_ & n31643;
  assign n31730 = ~n31726 & ~n31727;
  assign n31731 = ~n31728 & n31730;
  assign n31732 = ~n31729 & n31731;
  assign n31733 = n31711 & n31718;
  assign n31734 = n31725 & n31733;
  assign n31735 = n31732 & n31734;
  assign n31736 = n31509 & ~n31735;
  assign n31737 = P1_BUF2_REG_10_ & n31512;
  assign n31738 = P1_P3_EAX_REG_10_ & ~n31508;
  assign n31739 = P1_P3_EAX_REG_9_ & n31697;
  assign n31740 = ~P1_P3_EAX_REG_10_ & n31739;
  assign n31741 = P1_P3_EAX_REG_10_ & ~n31739;
  assign n31742 = ~n31740 & ~n31741;
  assign n31743 = n31515 & ~n31742;
  assign n31744 = ~n31738 & ~n31743;
  assign n31745 = ~n31736 & ~n31737;
  assign n4991 = ~n31744 | ~n31745;
  assign n31747 = P1_P3_INSTQUEUE_REG_15__3_ & n31601;
  assign n31748 = P1_P3_INSTQUEUE_REG_14__3_ & n31603;
  assign n31749 = P1_P3_INSTQUEUE_REG_13__3_ & n31605;
  assign n31750 = P1_P3_INSTQUEUE_REG_12__3_ & n31607;
  assign n31751 = ~n31747 & ~n31748;
  assign n31752 = ~n31749 & n31751;
  assign n31753 = ~n31750 & n31752;
  assign n31754 = P1_P3_INSTQUEUE_REG_11__3_ & n31613;
  assign n31755 = P1_P3_INSTQUEUE_REG_10__3_ & n31615;
  assign n31756 = P1_P3_INSTQUEUE_REG_9__3_ & n31617;
  assign n31757 = P1_P3_INSTQUEUE_REG_8__3_ & n31619;
  assign n31758 = ~n31754 & ~n31755;
  assign n31759 = ~n31756 & n31758;
  assign n31760 = ~n31757 & n31759;
  assign n31761 = P1_P3_INSTQUEUE_REG_7__3_ & n31625;
  assign n31762 = P1_P3_INSTQUEUE_REG_6__3_ & n31627;
  assign n31763 = P1_P3_INSTQUEUE_REG_5__3_ & n31629;
  assign n31764 = P1_P3_INSTQUEUE_REG_4__3_ & n31631;
  assign n31765 = ~n31761 & ~n31762;
  assign n31766 = ~n31763 & n31765;
  assign n31767 = ~n31764 & n31766;
  assign n31768 = P1_P3_INSTQUEUE_REG_3__3_ & n31637;
  assign n31769 = P1_P3_INSTQUEUE_REG_2__3_ & n31639;
  assign n31770 = P1_P3_INSTQUEUE_REG_1__3_ & n31641;
  assign n31771 = P1_P3_INSTQUEUE_REG_0__3_ & n31643;
  assign n31772 = ~n31768 & ~n31769;
  assign n31773 = ~n31770 & n31772;
  assign n31774 = ~n31771 & n31773;
  assign n31775 = n31753 & n31760;
  assign n31776 = n31767 & n31775;
  assign n31777 = n31774 & n31776;
  assign n31778 = n31509 & ~n31777;
  assign n31779 = P1_BUF2_REG_11_ & n31512;
  assign n31780 = P1_P3_EAX_REG_11_ & ~n31508;
  assign n31781 = P1_P3_EAX_REG_9_ & P1_P3_EAX_REG_10_;
  assign n31782 = n31697 & n31781;
  assign n31783 = P1_P3_EAX_REG_11_ & ~n31782;
  assign n31784 = ~P1_P3_EAX_REG_11_ & n31782;
  assign n31785 = ~n31783 & ~n31784;
  assign n31786 = n31515 & ~n31785;
  assign n31787 = ~n31780 & ~n31786;
  assign n31788 = ~n31778 & ~n31779;
  assign n4996 = ~n31787 | ~n31788;
  assign n31790 = P1_P3_INSTQUEUE_REG_15__4_ & n31601;
  assign n31791 = P1_P3_INSTQUEUE_REG_14__4_ & n31603;
  assign n31792 = P1_P3_INSTQUEUE_REG_13__4_ & n31605;
  assign n31793 = P1_P3_INSTQUEUE_REG_12__4_ & n31607;
  assign n31794 = ~n31790 & ~n31791;
  assign n31795 = ~n31792 & n31794;
  assign n31796 = ~n31793 & n31795;
  assign n31797 = P1_P3_INSTQUEUE_REG_11__4_ & n31613;
  assign n31798 = P1_P3_INSTQUEUE_REG_10__4_ & n31615;
  assign n31799 = P1_P3_INSTQUEUE_REG_9__4_ & n31617;
  assign n31800 = P1_P3_INSTQUEUE_REG_8__4_ & n31619;
  assign n31801 = ~n31797 & ~n31798;
  assign n31802 = ~n31799 & n31801;
  assign n31803 = ~n31800 & n31802;
  assign n31804 = P1_P3_INSTQUEUE_REG_7__4_ & n31625;
  assign n31805 = P1_P3_INSTQUEUE_REG_6__4_ & n31627;
  assign n31806 = P1_P3_INSTQUEUE_REG_5__4_ & n31629;
  assign n31807 = P1_P3_INSTQUEUE_REG_4__4_ & n31631;
  assign n31808 = ~n31804 & ~n31805;
  assign n31809 = ~n31806 & n31808;
  assign n31810 = ~n31807 & n31809;
  assign n31811 = P1_P3_INSTQUEUE_REG_3__4_ & n31637;
  assign n31812 = P1_P3_INSTQUEUE_REG_2__4_ & n31639;
  assign n31813 = P1_P3_INSTQUEUE_REG_1__4_ & n31641;
  assign n31814 = P1_P3_INSTQUEUE_REG_0__4_ & n31643;
  assign n31815 = ~n31811 & ~n31812;
  assign n31816 = ~n31813 & n31815;
  assign n31817 = ~n31814 & n31816;
  assign n31818 = n31796 & n31803;
  assign n31819 = n31810 & n31818;
  assign n31820 = n31817 & n31819;
  assign n31821 = n31509 & ~n31820;
  assign n31822 = P1_BUF2_REG_12_ & n31512;
  assign n31823 = P1_P3_EAX_REG_12_ & ~n31508;
  assign n31824 = P1_P3_EAX_REG_11_ & n31782;
  assign n31825 = ~P1_P3_EAX_REG_12_ & n31824;
  assign n31826 = P1_P3_EAX_REG_12_ & ~n31824;
  assign n31827 = ~n31825 & ~n31826;
  assign n31828 = n31515 & ~n31827;
  assign n31829 = ~n31823 & ~n31828;
  assign n31830 = ~n31821 & ~n31822;
  assign n5001 = ~n31829 | ~n31830;
  assign n31832 = P1_BUF2_REG_13_ & n31512;
  assign n31833 = P1_P3_INSTQUEUE_REG_15__5_ & n31601;
  assign n31834 = P1_P3_INSTQUEUE_REG_14__5_ & n31603;
  assign n31835 = P1_P3_INSTQUEUE_REG_13__5_ & n31605;
  assign n31836 = P1_P3_INSTQUEUE_REG_12__5_ & n31607;
  assign n31837 = ~n31833 & ~n31834;
  assign n31838 = ~n31835 & n31837;
  assign n31839 = ~n31836 & n31838;
  assign n31840 = P1_P3_INSTQUEUE_REG_11__5_ & n31613;
  assign n31841 = P1_P3_INSTQUEUE_REG_10__5_ & n31615;
  assign n31842 = P1_P3_INSTQUEUE_REG_9__5_ & n31617;
  assign n31843 = P1_P3_INSTQUEUE_REG_8__5_ & n31619;
  assign n31844 = ~n31840 & ~n31841;
  assign n31845 = ~n31842 & n31844;
  assign n31846 = ~n31843 & n31845;
  assign n31847 = P1_P3_INSTQUEUE_REG_7__5_ & n31625;
  assign n31848 = P1_P3_INSTQUEUE_REG_6__5_ & n31627;
  assign n31849 = P1_P3_INSTQUEUE_REG_5__5_ & n31629;
  assign n31850 = P1_P3_INSTQUEUE_REG_4__5_ & n31631;
  assign n31851 = ~n31847 & ~n31848;
  assign n31852 = ~n31849 & n31851;
  assign n31853 = ~n31850 & n31852;
  assign n31854 = P1_P3_INSTQUEUE_REG_3__5_ & n31637;
  assign n31855 = P1_P3_INSTQUEUE_REG_2__5_ & n31639;
  assign n31856 = P1_P3_INSTQUEUE_REG_1__5_ & n31641;
  assign n31857 = P1_P3_INSTQUEUE_REG_0__5_ & n31643;
  assign n31858 = ~n31854 & ~n31855;
  assign n31859 = ~n31856 & n31858;
  assign n31860 = ~n31857 & n31859;
  assign n31861 = n31839 & n31846;
  assign n31862 = n31853 & n31861;
  assign n31863 = n31860 & n31862;
  assign n31864 = n31509 & ~n31863;
  assign n31865 = P1_P3_EAX_REG_13_ & ~n31508;
  assign n31866 = ~n31864 & ~n31865;
  assign n31867 = P1_P3_EAX_REG_11_ & P1_P3_EAX_REG_12_;
  assign n31868 = n31782 & n31867;
  assign n31869 = P1_P3_EAX_REG_13_ & ~n31868;
  assign n31870 = ~P1_P3_EAX_REG_13_ & n31868;
  assign n31871 = ~n31869 & ~n31870;
  assign n31872 = n31515 & ~n31871;
  assign n31873 = ~n31832 & n31866;
  assign n5006 = n31872 | ~n31873;
  assign n31875 = P1_BUF2_REG_14_ & n31512;
  assign n31876 = P1_P3_INSTQUEUE_REG_15__6_ & n31601;
  assign n31877 = P1_P3_INSTQUEUE_REG_14__6_ & n31603;
  assign n31878 = P1_P3_INSTQUEUE_REG_13__6_ & n31605;
  assign n31879 = P1_P3_INSTQUEUE_REG_12__6_ & n31607;
  assign n31880 = ~n31876 & ~n31877;
  assign n31881 = ~n31878 & n31880;
  assign n31882 = ~n31879 & n31881;
  assign n31883 = P1_P3_INSTQUEUE_REG_11__6_ & n31613;
  assign n31884 = P1_P3_INSTQUEUE_REG_10__6_ & n31615;
  assign n31885 = P1_P3_INSTQUEUE_REG_9__6_ & n31617;
  assign n31886 = P1_P3_INSTQUEUE_REG_8__6_ & n31619;
  assign n31887 = ~n31883 & ~n31884;
  assign n31888 = ~n31885 & n31887;
  assign n31889 = ~n31886 & n31888;
  assign n31890 = P1_P3_INSTQUEUE_REG_7__6_ & n31625;
  assign n31891 = P1_P3_INSTQUEUE_REG_6__6_ & n31627;
  assign n31892 = P1_P3_INSTQUEUE_REG_5__6_ & n31629;
  assign n31893 = P1_P3_INSTQUEUE_REG_4__6_ & n31631;
  assign n31894 = ~n31890 & ~n31891;
  assign n31895 = ~n31892 & n31894;
  assign n31896 = ~n31893 & n31895;
  assign n31897 = P1_P3_INSTQUEUE_REG_3__6_ & n31637;
  assign n31898 = P1_P3_INSTQUEUE_REG_2__6_ & n31639;
  assign n31899 = P1_P3_INSTQUEUE_REG_1__6_ & n31641;
  assign n31900 = P1_P3_INSTQUEUE_REG_0__6_ & n31643;
  assign n31901 = ~n31897 & ~n31898;
  assign n31902 = ~n31899 & n31901;
  assign n31903 = ~n31900 & n31902;
  assign n31904 = n31882 & n31889;
  assign n31905 = n31896 & n31904;
  assign n31906 = n31903 & n31905;
  assign n31907 = n31509 & ~n31906;
  assign n31908 = P1_P3_EAX_REG_14_ & ~n31508;
  assign n31909 = ~n31907 & ~n31908;
  assign n31910 = P1_P3_EAX_REG_13_ & n31868;
  assign n31911 = ~P1_P3_EAX_REG_14_ & n31910;
  assign n31912 = P1_P3_EAX_REG_14_ & ~n31910;
  assign n31913 = ~n31911 & ~n31912;
  assign n31914 = n31515 & ~n31913;
  assign n31915 = ~n31875 & n31909;
  assign n5011 = n31914 | ~n31915;
  assign n31917 = P1_BUF2_REG_15_ & n31512;
  assign n31918 = P1_P3_INSTQUEUE_REG_15__7_ & n31601;
  assign n31919 = P1_P3_INSTQUEUE_REG_14__7_ & n31603;
  assign n31920 = P1_P3_INSTQUEUE_REG_13__7_ & n31605;
  assign n31921 = P1_P3_INSTQUEUE_REG_12__7_ & n31607;
  assign n31922 = ~n31918 & ~n31919;
  assign n31923 = ~n31920 & n31922;
  assign n31924 = ~n31921 & n31923;
  assign n31925 = P1_P3_INSTQUEUE_REG_11__7_ & n31613;
  assign n31926 = P1_P3_INSTQUEUE_REG_10__7_ & n31615;
  assign n31927 = P1_P3_INSTQUEUE_REG_9__7_ & n31617;
  assign n31928 = P1_P3_INSTQUEUE_REG_8__7_ & n31619;
  assign n31929 = ~n31925 & ~n31926;
  assign n31930 = ~n31927 & n31929;
  assign n31931 = ~n31928 & n31930;
  assign n31932 = P1_P3_INSTQUEUE_REG_7__7_ & n31625;
  assign n31933 = P1_P3_INSTQUEUE_REG_6__7_ & n31627;
  assign n31934 = P1_P3_INSTQUEUE_REG_5__7_ & n31629;
  assign n31935 = P1_P3_INSTQUEUE_REG_4__7_ & n31631;
  assign n31936 = ~n31932 & ~n31933;
  assign n31937 = ~n31934 & n31936;
  assign n31938 = ~n31935 & n31937;
  assign n31939 = P1_P3_INSTQUEUE_REG_3__7_ & n31637;
  assign n31940 = P1_P3_INSTQUEUE_REG_2__7_ & n31639;
  assign n31941 = P1_P3_INSTQUEUE_REG_1__7_ & n31641;
  assign n31942 = P1_P3_INSTQUEUE_REG_0__7_ & n31643;
  assign n31943 = ~n31939 & ~n31940;
  assign n31944 = ~n31941 & n31943;
  assign n31945 = ~n31942 & n31944;
  assign n31946 = n31924 & n31931;
  assign n31947 = n31938 & n31946;
  assign n31948 = n31945 & n31947;
  assign n31949 = n31509 & ~n31948;
  assign n31950 = P1_P3_EAX_REG_15_ & ~n31508;
  assign n31951 = ~n31949 & ~n31950;
  assign n31952 = P1_P3_EAX_REG_13_ & P1_P3_EAX_REG_14_;
  assign n31953 = n31868 & n31952;
  assign n31954 = P1_P3_EAX_REG_15_ & ~n31953;
  assign n31955 = ~P1_P3_EAX_REG_15_ & n31953;
  assign n31956 = ~n31954 & ~n31955;
  assign n31957 = n31515 & ~n31956;
  assign n31958 = ~n31917 & n31951;
  assign n5016 = n31957 | ~n31958;
  assign n31960 = ~n25448 & n31511;
  assign n31961 = P1_BUF2_REG_16_ & n31960;
  assign n31962 = n25417 & n31511;
  assign n31963 = P1_BUF2_REG_0_ & n31962;
  assign n31964 = P1_P3_EAX_REG_16_ & ~n31508;
  assign n31965 = P1_P3_INSTQUEUERD_ADDR_REG_2_ & ~n25373;
  assign n31966 = ~P1_P3_INSTQUEUERD_ADDR_REG_3_ & n31965;
  assign n31967 = P1_P3_INSTQUEUERD_ADDR_REG_3_ & ~n31965;
  assign n31968 = ~n31966 & ~n31967;
  assign n31969 = ~n25374 & ~n31965;
  assign n31970 = n31968 & n31969;
  assign n31971 = n27654 & n31970;
  assign n31972 = P1_P3_INSTQUEUE_REG_7__0_ & n31971;
  assign n31973 = n27651 & n31970;
  assign n31974 = P1_P3_INSTQUEUE_REG_6__0_ & n31973;
  assign n31975 = n27660 & n31970;
  assign n31976 = P1_P3_INSTQUEUE_REG_5__0_ & n31975;
  assign n31977 = n27657 & n31970;
  assign n31978 = P1_P3_INSTQUEUE_REG_4__0_ & n31977;
  assign n31979 = ~n31972 & ~n31974;
  assign n31980 = ~n31976 & n31979;
  assign n31981 = ~n31978 & n31980;
  assign n31982 = n31968 & ~n31969;
  assign n31983 = n27654 & n31982;
  assign n31984 = P1_P3_INSTQUEUE_REG_3__0_ & n31983;
  assign n31985 = n27651 & n31982;
  assign n31986 = P1_P3_INSTQUEUE_REG_2__0_ & n31985;
  assign n31987 = n27660 & n31982;
  assign n31988 = P1_P3_INSTQUEUE_REG_1__0_ & n31987;
  assign n31989 = n27657 & n31982;
  assign n31990 = P1_P3_INSTQUEUE_REG_0__0_ & n31989;
  assign n31991 = ~n31984 & ~n31986;
  assign n31992 = ~n31988 & n31991;
  assign n31993 = ~n31990 & n31992;
  assign n31994 = ~n31968 & n31969;
  assign n31995 = n27654 & n31994;
  assign n31996 = P1_P3_INSTQUEUE_REG_15__0_ & n31995;
  assign n31997 = n27651 & n31994;
  assign n31998 = P1_P3_INSTQUEUE_REG_14__0_ & n31997;
  assign n31999 = n27660 & n31994;
  assign n32000 = P1_P3_INSTQUEUE_REG_13__0_ & n31999;
  assign n32001 = n27657 & n31994;
  assign n32002 = P1_P3_INSTQUEUE_REG_12__0_ & n32001;
  assign n32003 = ~n31996 & ~n31998;
  assign n32004 = ~n32000 & n32003;
  assign n32005 = ~n32002 & n32004;
  assign n32006 = ~n31968 & ~n31969;
  assign n32007 = n27654 & n32006;
  assign n32008 = P1_P3_INSTQUEUE_REG_11__0_ & n32007;
  assign n32009 = n27651 & n32006;
  assign n32010 = P1_P3_INSTQUEUE_REG_10__0_ & n32009;
  assign n32011 = n27660 & n32006;
  assign n32012 = P1_P3_INSTQUEUE_REG_9__0_ & n32011;
  assign n32013 = n27657 & n32006;
  assign n32014 = P1_P3_INSTQUEUE_REG_8__0_ & n32013;
  assign n32015 = ~n32008 & ~n32010;
  assign n32016 = ~n32012 & n32015;
  assign n32017 = ~n32014 & n32016;
  assign n32018 = n31981 & n31993;
  assign n32019 = n32005 & n32018;
  assign n32020 = n32017 & n32019;
  assign n32021 = n31509 & ~n32020;
  assign n32022 = ~n31964 & ~n32021;
  assign n32023 = P1_P3_EAX_REG_15_ & n31953;
  assign n32024 = ~P1_P3_EAX_REG_16_ & n32023;
  assign n32025 = P1_P3_EAX_REG_16_ & ~n32023;
  assign n32026 = ~n32024 & ~n32025;
  assign n32027 = n31515 & ~n32026;
  assign n32028 = ~n31961 & ~n31963;
  assign n32029 = n32022 & n32028;
  assign n5021 = n32027 | ~n32029;
  assign n32031 = P1_BUF2_REG_17_ & n31960;
  assign n32032 = P1_BUF2_REG_1_ & n31962;
  assign n32033 = P1_P3_EAX_REG_17_ & ~n31508;
  assign n32034 = P1_P3_INSTQUEUE_REG_7__1_ & n31971;
  assign n32035 = P1_P3_INSTQUEUE_REG_6__1_ & n31973;
  assign n32036 = P1_P3_INSTQUEUE_REG_5__1_ & n31975;
  assign n32037 = P1_P3_INSTQUEUE_REG_4__1_ & n31977;
  assign n32038 = ~n32034 & ~n32035;
  assign n32039 = ~n32036 & n32038;
  assign n32040 = ~n32037 & n32039;
  assign n32041 = P1_P3_INSTQUEUE_REG_3__1_ & n31983;
  assign n32042 = P1_P3_INSTQUEUE_REG_2__1_ & n31985;
  assign n32043 = P1_P3_INSTQUEUE_REG_1__1_ & n31987;
  assign n32044 = P1_P3_INSTQUEUE_REG_0__1_ & n31989;
  assign n32045 = ~n32041 & ~n32042;
  assign n32046 = ~n32043 & n32045;
  assign n32047 = ~n32044 & n32046;
  assign n32048 = P1_P3_INSTQUEUE_REG_15__1_ & n31995;
  assign n32049 = P1_P3_INSTQUEUE_REG_14__1_ & n31997;
  assign n32050 = P1_P3_INSTQUEUE_REG_13__1_ & n31999;
  assign n32051 = P1_P3_INSTQUEUE_REG_12__1_ & n32001;
  assign n32052 = ~n32048 & ~n32049;
  assign n32053 = ~n32050 & n32052;
  assign n32054 = ~n32051 & n32053;
  assign n32055 = P1_P3_INSTQUEUE_REG_11__1_ & n32007;
  assign n32056 = P1_P3_INSTQUEUE_REG_10__1_ & n32009;
  assign n32057 = P1_P3_INSTQUEUE_REG_9__1_ & n32011;
  assign n32058 = P1_P3_INSTQUEUE_REG_8__1_ & n32013;
  assign n32059 = ~n32055 & ~n32056;
  assign n32060 = ~n32057 & n32059;
  assign n32061 = ~n32058 & n32060;
  assign n32062 = n32040 & n32047;
  assign n32063 = n32054 & n32062;
  assign n32064 = n32061 & n32063;
  assign n32065 = n31509 & ~n32064;
  assign n32066 = ~n32033 & ~n32065;
  assign n32067 = P1_P3_EAX_REG_15_ & P1_P3_EAX_REG_16_;
  assign n32068 = n31953 & n32067;
  assign n32069 = P1_P3_EAX_REG_17_ & ~n32068;
  assign n32070 = ~P1_P3_EAX_REG_17_ & n32068;
  assign n32071 = ~n32069 & ~n32070;
  assign n32072 = n31515 & ~n32071;
  assign n32073 = ~n32031 & ~n32032;
  assign n32074 = n32066 & n32073;
  assign n5026 = n32072 | ~n32074;
  assign n32076 = P1_BUF2_REG_18_ & n31960;
  assign n32077 = P1_BUF2_REG_2_ & n31962;
  assign n32078 = P1_P3_EAX_REG_18_ & ~n31508;
  assign n32079 = P1_P3_INSTQUEUE_REG_7__2_ & n31971;
  assign n32080 = P1_P3_INSTQUEUE_REG_6__2_ & n31973;
  assign n32081 = P1_P3_INSTQUEUE_REG_5__2_ & n31975;
  assign n32082 = P1_P3_INSTQUEUE_REG_4__2_ & n31977;
  assign n32083 = ~n32079 & ~n32080;
  assign n32084 = ~n32081 & n32083;
  assign n32085 = ~n32082 & n32084;
  assign n32086 = P1_P3_INSTQUEUE_REG_3__2_ & n31983;
  assign n32087 = P1_P3_INSTQUEUE_REG_2__2_ & n31985;
  assign n32088 = P1_P3_INSTQUEUE_REG_1__2_ & n31987;
  assign n32089 = P1_P3_INSTQUEUE_REG_0__2_ & n31989;
  assign n32090 = ~n32086 & ~n32087;
  assign n32091 = ~n32088 & n32090;
  assign n32092 = ~n32089 & n32091;
  assign n32093 = P1_P3_INSTQUEUE_REG_15__2_ & n31995;
  assign n32094 = P1_P3_INSTQUEUE_REG_14__2_ & n31997;
  assign n32095 = P1_P3_INSTQUEUE_REG_13__2_ & n31999;
  assign n32096 = P1_P3_INSTQUEUE_REG_12__2_ & n32001;
  assign n32097 = ~n32093 & ~n32094;
  assign n32098 = ~n32095 & n32097;
  assign n32099 = ~n32096 & n32098;
  assign n32100 = P1_P3_INSTQUEUE_REG_11__2_ & n32007;
  assign n32101 = P1_P3_INSTQUEUE_REG_10__2_ & n32009;
  assign n32102 = P1_P3_INSTQUEUE_REG_9__2_ & n32011;
  assign n32103 = P1_P3_INSTQUEUE_REG_8__2_ & n32013;
  assign n32104 = ~n32100 & ~n32101;
  assign n32105 = ~n32102 & n32104;
  assign n32106 = ~n32103 & n32105;
  assign n32107 = n32085 & n32092;
  assign n32108 = n32099 & n32107;
  assign n32109 = n32106 & n32108;
  assign n32110 = n31509 & ~n32109;
  assign n32111 = ~n32078 & ~n32110;
  assign n32112 = P1_P3_EAX_REG_17_ & n32068;
  assign n32113 = ~P1_P3_EAX_REG_18_ & n32112;
  assign n32114 = P1_P3_EAX_REG_18_ & ~n32112;
  assign n32115 = ~n32113 & ~n32114;
  assign n32116 = n31515 & ~n32115;
  assign n32117 = ~n32076 & ~n32077;
  assign n32118 = n32111 & n32117;
  assign n5031 = n32116 | ~n32118;
  assign n32120 = P1_BUF2_REG_19_ & n31960;
  assign n32121 = P1_BUF2_REG_3_ & n31962;
  assign n32122 = P1_P3_EAX_REG_19_ & ~n31508;
  assign n32123 = P1_P3_INSTQUEUE_REG_7__3_ & n31971;
  assign n32124 = P1_P3_INSTQUEUE_REG_6__3_ & n31973;
  assign n32125 = P1_P3_INSTQUEUE_REG_5__3_ & n31975;
  assign n32126 = P1_P3_INSTQUEUE_REG_4__3_ & n31977;
  assign n32127 = ~n32123 & ~n32124;
  assign n32128 = ~n32125 & n32127;
  assign n32129 = ~n32126 & n32128;
  assign n32130 = P1_P3_INSTQUEUE_REG_3__3_ & n31983;
  assign n32131 = P1_P3_INSTQUEUE_REG_2__3_ & n31985;
  assign n32132 = P1_P3_INSTQUEUE_REG_1__3_ & n31987;
  assign n32133 = P1_P3_INSTQUEUE_REG_0__3_ & n31989;
  assign n32134 = ~n32130 & ~n32131;
  assign n32135 = ~n32132 & n32134;
  assign n32136 = ~n32133 & n32135;
  assign n32137 = P1_P3_INSTQUEUE_REG_15__3_ & n31995;
  assign n32138 = P1_P3_INSTQUEUE_REG_14__3_ & n31997;
  assign n32139 = P1_P3_INSTQUEUE_REG_13__3_ & n31999;
  assign n32140 = P1_P3_INSTQUEUE_REG_12__3_ & n32001;
  assign n32141 = ~n32137 & ~n32138;
  assign n32142 = ~n32139 & n32141;
  assign n32143 = ~n32140 & n32142;
  assign n32144 = P1_P3_INSTQUEUE_REG_11__3_ & n32007;
  assign n32145 = P1_P3_INSTQUEUE_REG_10__3_ & n32009;
  assign n32146 = P1_P3_INSTQUEUE_REG_9__3_ & n32011;
  assign n32147 = P1_P3_INSTQUEUE_REG_8__3_ & n32013;
  assign n32148 = ~n32144 & ~n32145;
  assign n32149 = ~n32146 & n32148;
  assign n32150 = ~n32147 & n32149;
  assign n32151 = n32129 & n32136;
  assign n32152 = n32143 & n32151;
  assign n32153 = n32150 & n32152;
  assign n32154 = n31509 & ~n32153;
  assign n32155 = ~n32122 & ~n32154;
  assign n32156 = P1_P3_EAX_REG_17_ & P1_P3_EAX_REG_18_;
  assign n32157 = n32068 & n32156;
  assign n32158 = P1_P3_EAX_REG_19_ & ~n32157;
  assign n32159 = ~P1_P3_EAX_REG_19_ & n32157;
  assign n32160 = ~n32158 & ~n32159;
  assign n32161 = n31515 & ~n32160;
  assign n32162 = ~n32120 & ~n32121;
  assign n32163 = n32155 & n32162;
  assign n5036 = n32161 | ~n32163;
  assign n32165 = P1_BUF2_REG_20_ & n31960;
  assign n32166 = P1_BUF2_REG_4_ & n31962;
  assign n32167 = P1_P3_EAX_REG_20_ & ~n31508;
  assign n32168 = P1_P3_INSTQUEUE_REG_7__4_ & n31971;
  assign n32169 = P1_P3_INSTQUEUE_REG_6__4_ & n31973;
  assign n32170 = P1_P3_INSTQUEUE_REG_5__4_ & n31975;
  assign n32171 = P1_P3_INSTQUEUE_REG_4__4_ & n31977;
  assign n32172 = ~n32168 & ~n32169;
  assign n32173 = ~n32170 & n32172;
  assign n32174 = ~n32171 & n32173;
  assign n32175 = P1_P3_INSTQUEUE_REG_3__4_ & n31983;
  assign n32176 = P1_P3_INSTQUEUE_REG_2__4_ & n31985;
  assign n32177 = P1_P3_INSTQUEUE_REG_1__4_ & n31987;
  assign n32178 = P1_P3_INSTQUEUE_REG_0__4_ & n31989;
  assign n32179 = ~n32175 & ~n32176;
  assign n32180 = ~n32177 & n32179;
  assign n32181 = ~n32178 & n32180;
  assign n32182 = P1_P3_INSTQUEUE_REG_15__4_ & n31995;
  assign n32183 = P1_P3_INSTQUEUE_REG_14__4_ & n31997;
  assign n32184 = P1_P3_INSTQUEUE_REG_13__4_ & n31999;
  assign n32185 = P1_P3_INSTQUEUE_REG_12__4_ & n32001;
  assign n32186 = ~n32182 & ~n32183;
  assign n32187 = ~n32184 & n32186;
  assign n32188 = ~n32185 & n32187;
  assign n32189 = P1_P3_INSTQUEUE_REG_11__4_ & n32007;
  assign n32190 = P1_P3_INSTQUEUE_REG_10__4_ & n32009;
  assign n32191 = P1_P3_INSTQUEUE_REG_9__4_ & n32011;
  assign n32192 = P1_P3_INSTQUEUE_REG_8__4_ & n32013;
  assign n32193 = ~n32189 & ~n32190;
  assign n32194 = ~n32191 & n32193;
  assign n32195 = ~n32192 & n32194;
  assign n32196 = n32174 & n32181;
  assign n32197 = n32188 & n32196;
  assign n32198 = n32195 & n32197;
  assign n32199 = n31509 & ~n32198;
  assign n32200 = ~n32167 & ~n32199;
  assign n32201 = P1_P3_EAX_REG_19_ & n32157;
  assign n32202 = ~P1_P3_EAX_REG_20_ & n32201;
  assign n32203 = P1_P3_EAX_REG_20_ & ~n32201;
  assign n32204 = ~n32202 & ~n32203;
  assign n32205 = n31515 & ~n32204;
  assign n32206 = ~n32165 & ~n32166;
  assign n32207 = n32200 & n32206;
  assign n5041 = n32205 | ~n32207;
  assign n32209 = P1_BUF2_REG_21_ & n31960;
  assign n32210 = P1_BUF2_REG_5_ & n31962;
  assign n32211 = P1_P3_EAX_REG_21_ & ~n31508;
  assign n32212 = P1_P3_INSTQUEUE_REG_7__5_ & n31971;
  assign n32213 = P1_P3_INSTQUEUE_REG_6__5_ & n31973;
  assign n32214 = P1_P3_INSTQUEUE_REG_5__5_ & n31975;
  assign n32215 = P1_P3_INSTQUEUE_REG_4__5_ & n31977;
  assign n32216 = ~n32212 & ~n32213;
  assign n32217 = ~n32214 & n32216;
  assign n32218 = ~n32215 & n32217;
  assign n32219 = P1_P3_INSTQUEUE_REG_3__5_ & n31983;
  assign n32220 = P1_P3_INSTQUEUE_REG_2__5_ & n31985;
  assign n32221 = P1_P3_INSTQUEUE_REG_1__5_ & n31987;
  assign n32222 = P1_P3_INSTQUEUE_REG_0__5_ & n31989;
  assign n32223 = ~n32219 & ~n32220;
  assign n32224 = ~n32221 & n32223;
  assign n32225 = ~n32222 & n32224;
  assign n32226 = P1_P3_INSTQUEUE_REG_15__5_ & n31995;
  assign n32227 = P1_P3_INSTQUEUE_REG_14__5_ & n31997;
  assign n32228 = P1_P3_INSTQUEUE_REG_13__5_ & n31999;
  assign n32229 = P1_P3_INSTQUEUE_REG_12__5_ & n32001;
  assign n32230 = ~n32226 & ~n32227;
  assign n32231 = ~n32228 & n32230;
  assign n32232 = ~n32229 & n32231;
  assign n32233 = P1_P3_INSTQUEUE_REG_11__5_ & n32007;
  assign n32234 = P1_P3_INSTQUEUE_REG_10__5_ & n32009;
  assign n32235 = P1_P3_INSTQUEUE_REG_9__5_ & n32011;
  assign n32236 = P1_P3_INSTQUEUE_REG_8__5_ & n32013;
  assign n32237 = ~n32233 & ~n32234;
  assign n32238 = ~n32235 & n32237;
  assign n32239 = ~n32236 & n32238;
  assign n32240 = n32218 & n32225;
  assign n32241 = n32232 & n32240;
  assign n32242 = n32239 & n32241;
  assign n32243 = n31509 & ~n32242;
  assign n32244 = ~n32211 & ~n32243;
  assign n32245 = P1_P3_EAX_REG_19_ & P1_P3_EAX_REG_20_;
  assign n32246 = n32157 & n32245;
  assign n32247 = P1_P3_EAX_REG_21_ & ~n32246;
  assign n32248 = ~P1_P3_EAX_REG_21_ & n32246;
  assign n32249 = ~n32247 & ~n32248;
  assign n32250 = n31515 & ~n32249;
  assign n32251 = ~n32209 & ~n32210;
  assign n32252 = n32244 & n32251;
  assign n5046 = n32250 | ~n32252;
  assign n32254 = P1_BUF2_REG_22_ & n31960;
  assign n32255 = P1_BUF2_REG_6_ & n31962;
  assign n32256 = P1_P3_EAX_REG_22_ & ~n31508;
  assign n32257 = P1_P3_INSTQUEUE_REG_7__6_ & n31971;
  assign n32258 = P1_P3_INSTQUEUE_REG_6__6_ & n31973;
  assign n32259 = P1_P3_INSTQUEUE_REG_5__6_ & n31975;
  assign n32260 = P1_P3_INSTQUEUE_REG_4__6_ & n31977;
  assign n32261 = ~n32257 & ~n32258;
  assign n32262 = ~n32259 & n32261;
  assign n32263 = ~n32260 & n32262;
  assign n32264 = P1_P3_INSTQUEUE_REG_3__6_ & n31983;
  assign n32265 = P1_P3_INSTQUEUE_REG_2__6_ & n31985;
  assign n32266 = P1_P3_INSTQUEUE_REG_1__6_ & n31987;
  assign n32267 = P1_P3_INSTQUEUE_REG_0__6_ & n31989;
  assign n32268 = ~n32264 & ~n32265;
  assign n32269 = ~n32266 & n32268;
  assign n32270 = ~n32267 & n32269;
  assign n32271 = P1_P3_INSTQUEUE_REG_15__6_ & n31995;
  assign n32272 = P1_P3_INSTQUEUE_REG_14__6_ & n31997;
  assign n32273 = P1_P3_INSTQUEUE_REG_13__6_ & n31999;
  assign n32274 = P1_P3_INSTQUEUE_REG_12__6_ & n32001;
  assign n32275 = ~n32271 & ~n32272;
  assign n32276 = ~n32273 & n32275;
  assign n32277 = ~n32274 & n32276;
  assign n32278 = P1_P3_INSTQUEUE_REG_11__6_ & n32007;
  assign n32279 = P1_P3_INSTQUEUE_REG_10__6_ & n32009;
  assign n32280 = P1_P3_INSTQUEUE_REG_9__6_ & n32011;
  assign n32281 = P1_P3_INSTQUEUE_REG_8__6_ & n32013;
  assign n32282 = ~n32278 & ~n32279;
  assign n32283 = ~n32280 & n32282;
  assign n32284 = ~n32281 & n32283;
  assign n32285 = n32263 & n32270;
  assign n32286 = n32277 & n32285;
  assign n32287 = n32284 & n32286;
  assign n32288 = n31509 & ~n32287;
  assign n32289 = ~n32256 & ~n32288;
  assign n32290 = P1_P3_EAX_REG_21_ & n32246;
  assign n32291 = ~P1_P3_EAX_REG_22_ & n32290;
  assign n32292 = P1_P3_EAX_REG_22_ & ~n32290;
  assign n32293 = ~n32291 & ~n32292;
  assign n32294 = n31515 & ~n32293;
  assign n32295 = ~n32254 & ~n32255;
  assign n32296 = n32289 & n32295;
  assign n5051 = n32294 | ~n32296;
  assign n32298 = P1_BUF2_REG_23_ & n31960;
  assign n32299 = P1_BUF2_REG_7_ & n31962;
  assign n32300 = P1_P3_EAX_REG_23_ & ~n31508;
  assign n32301 = P1_P3_INSTQUEUERD_ADDR_REG_3_ & ~P1_P3_INSTQUEUERD_ADDR_REG_2_;
  assign n32302 = ~n25390 & ~n32301;
  assign n32303 = n25361 & n32302;
  assign n32304 = P1_P3_INSTQUEUE_REG_7__0_ & n32303;
  assign n32305 = n25365 & n32302;
  assign n32306 = P1_P3_INSTQUEUE_REG_6__0_ & n32305;
  assign n32307 = n25370 & n32302;
  assign n32308 = P1_P3_INSTQUEUE_REG_5__0_ & n32307;
  assign n32309 = n25374 & n32302;
  assign n32310 = P1_P3_INSTQUEUE_REG_4__0_ & n32309;
  assign n32311 = ~n32304 & ~n32306;
  assign n32312 = ~n32308 & n32311;
  assign n32313 = ~n32310 & n32312;
  assign n32314 = P1_P3_INSTQUEUERD_ADDR_REG_2_ & n32302;
  assign n32315 = n25360 & n32314;
  assign n32316 = P1_P3_INSTQUEUE_REG_3__0_ & n32315;
  assign n32317 = n25364 & n32314;
  assign n32318 = P1_P3_INSTQUEUE_REG_2__0_ & n32317;
  assign n32319 = n25369 & n32314;
  assign n32320 = P1_P3_INSTQUEUE_REG_1__0_ & n32319;
  assign n32321 = n25373 & n32314;
  assign n32322 = P1_P3_INSTQUEUE_REG_0__0_ & n32321;
  assign n32323 = ~n32316 & ~n32318;
  assign n32324 = ~n32320 & n32323;
  assign n32325 = ~n32322 & n32324;
  assign n32326 = n25361 & ~n32302;
  assign n32327 = P1_P3_INSTQUEUE_REG_15__0_ & n32326;
  assign n32328 = n25365 & ~n32302;
  assign n32329 = P1_P3_INSTQUEUE_REG_14__0_ & n32328;
  assign n32330 = n25370 & ~n32302;
  assign n32331 = P1_P3_INSTQUEUE_REG_13__0_ & n32330;
  assign n32332 = n25374 & ~n32302;
  assign n32333 = P1_P3_INSTQUEUE_REG_12__0_ & n32332;
  assign n32334 = ~n32327 & ~n32329;
  assign n32335 = ~n32331 & n32334;
  assign n32336 = ~n32333 & n32335;
  assign n32337 = P1_P3_INSTQUEUERD_ADDR_REG_2_ & ~n32302;
  assign n32338 = n25360 & n32337;
  assign n32339 = P1_P3_INSTQUEUE_REG_11__0_ & n32338;
  assign n32340 = n25364 & n32337;
  assign n32341 = P1_P3_INSTQUEUE_REG_10__0_ & n32340;
  assign n32342 = n25369 & n32337;
  assign n32343 = P1_P3_INSTQUEUE_REG_9__0_ & n32342;
  assign n32344 = n25373 & n32337;
  assign n32345 = P1_P3_INSTQUEUE_REG_8__0_ & n32344;
  assign n32346 = ~n32339 & ~n32341;
  assign n32347 = ~n32343 & n32346;
  assign n32348 = ~n32345 & n32347;
  assign n32349 = n32313 & n32325;
  assign n32350 = n32336 & n32349;
  assign n32351 = n32348 & n32350;
  assign n32352 = P1_P3_INSTQUEUE_REG_7__7_ & n31971;
  assign n32353 = P1_P3_INSTQUEUE_REG_6__7_ & n31973;
  assign n32354 = P1_P3_INSTQUEUE_REG_5__7_ & n31975;
  assign n32355 = P1_P3_INSTQUEUE_REG_4__7_ & n31977;
  assign n32356 = ~n32352 & ~n32353;
  assign n32357 = ~n32354 & n32356;
  assign n32358 = ~n32355 & n32357;
  assign n32359 = P1_P3_INSTQUEUE_REG_3__7_ & n31983;
  assign n32360 = P1_P3_INSTQUEUE_REG_2__7_ & n31985;
  assign n32361 = P1_P3_INSTQUEUE_REG_1__7_ & n31987;
  assign n32362 = P1_P3_INSTQUEUE_REG_0__7_ & n31989;
  assign n32363 = ~n32359 & ~n32360;
  assign n32364 = ~n32361 & n32363;
  assign n32365 = ~n32362 & n32364;
  assign n32366 = P1_P3_INSTQUEUE_REG_15__7_ & n31995;
  assign n32367 = P1_P3_INSTQUEUE_REG_14__7_ & n31997;
  assign n32368 = P1_P3_INSTQUEUE_REG_13__7_ & n31999;
  assign n32369 = P1_P3_INSTQUEUE_REG_12__7_ & n32001;
  assign n32370 = ~n32366 & ~n32367;
  assign n32371 = ~n32368 & n32370;
  assign n32372 = ~n32369 & n32371;
  assign n32373 = P1_P3_INSTQUEUE_REG_11__7_ & n32007;
  assign n32374 = P1_P3_INSTQUEUE_REG_10__7_ & n32009;
  assign n32375 = P1_P3_INSTQUEUE_REG_9__7_ & n32011;
  assign n32376 = P1_P3_INSTQUEUE_REG_8__7_ & n32013;
  assign n32377 = ~n32373 & ~n32374;
  assign n32378 = ~n32375 & n32377;
  assign n32379 = ~n32376 & n32378;
  assign n32380 = n32358 & n32365;
  assign n32381 = n32372 & n32380;
  assign n32382 = n32379 & n32381;
  assign n32383 = ~n32351 & n32382;
  assign n32384 = n32351 & ~n32382;
  assign n32385 = ~n32383 & ~n32384;
  assign n32386 = n31509 & ~n32385;
  assign n32387 = ~n32300 & ~n32386;
  assign n32388 = P1_P3_EAX_REG_21_ & P1_P3_EAX_REG_22_;
  assign n32389 = n32246 & n32388;
  assign n32390 = P1_P3_EAX_REG_23_ & ~n32389;
  assign n32391 = ~P1_P3_EAX_REG_23_ & n32389;
  assign n32392 = ~n32390 & ~n32391;
  assign n32393 = n31515 & ~n32392;
  assign n32394 = ~n32298 & ~n32299;
  assign n32395 = n32387 & n32394;
  assign n5056 = n32393 | ~n32395;
  assign n32397 = P1_BUF2_REG_24_ & n31960;
  assign n32398 = P1_BUF2_REG_8_ & n31962;
  assign n32399 = P1_P3_EAX_REG_24_ & ~n31508;
  assign n32400 = ~n32351 & ~n32382;
  assign n32401 = P1_P3_INSTQUEUE_REG_7__1_ & n32303;
  assign n32402 = P1_P3_INSTQUEUE_REG_6__1_ & n32305;
  assign n32403 = P1_P3_INSTQUEUE_REG_5__1_ & n32307;
  assign n32404 = P1_P3_INSTQUEUE_REG_4__1_ & n32309;
  assign n32405 = ~n32401 & ~n32402;
  assign n32406 = ~n32403 & n32405;
  assign n32407 = ~n32404 & n32406;
  assign n32408 = P1_P3_INSTQUEUE_REG_3__1_ & n32315;
  assign n32409 = P1_P3_INSTQUEUE_REG_2__1_ & n32317;
  assign n32410 = P1_P3_INSTQUEUE_REG_1__1_ & n32319;
  assign n32411 = P1_P3_INSTQUEUE_REG_0__1_ & n32321;
  assign n32412 = ~n32408 & ~n32409;
  assign n32413 = ~n32410 & n32412;
  assign n32414 = ~n32411 & n32413;
  assign n32415 = P1_P3_INSTQUEUE_REG_15__1_ & n32326;
  assign n32416 = P1_P3_INSTQUEUE_REG_14__1_ & n32328;
  assign n32417 = P1_P3_INSTQUEUE_REG_13__1_ & n32330;
  assign n32418 = P1_P3_INSTQUEUE_REG_12__1_ & n32332;
  assign n32419 = ~n32415 & ~n32416;
  assign n32420 = ~n32417 & n32419;
  assign n32421 = ~n32418 & n32420;
  assign n32422 = P1_P3_INSTQUEUE_REG_11__1_ & n32338;
  assign n32423 = P1_P3_INSTQUEUE_REG_10__1_ & n32340;
  assign n32424 = P1_P3_INSTQUEUE_REG_9__1_ & n32342;
  assign n32425 = P1_P3_INSTQUEUE_REG_8__1_ & n32344;
  assign n32426 = ~n32422 & ~n32423;
  assign n32427 = ~n32424 & n32426;
  assign n32428 = ~n32425 & n32427;
  assign n32429 = n32407 & n32414;
  assign n32430 = n32421 & n32429;
  assign n32431 = n32428 & n32430;
  assign n32432 = n32400 & n32431;
  assign n32433 = ~n32400 & ~n32431;
  assign n32434 = ~n32432 & ~n32433;
  assign n32435 = n31509 & ~n32434;
  assign n32436 = ~n32399 & ~n32435;
  assign n32437 = P1_P3_EAX_REG_23_ & n32389;
  assign n32438 = ~P1_P3_EAX_REG_24_ & n32437;
  assign n32439 = P1_P3_EAX_REG_24_ & ~n32437;
  assign n32440 = ~n32438 & ~n32439;
  assign n32441 = n31515 & ~n32440;
  assign n32442 = ~n32397 & ~n32398;
  assign n32443 = n32436 & n32442;
  assign n5061 = n32441 | ~n32443;
  assign n32445 = P1_BUF2_REG_25_ & n31960;
  assign n32446 = P1_BUF2_REG_9_ & n31962;
  assign n32447 = P1_P3_EAX_REG_25_ & ~n31508;
  assign n32448 = n32400 & ~n32431;
  assign n32449 = P1_P3_INSTQUEUE_REG_7__2_ & n32303;
  assign n32450 = P1_P3_INSTQUEUE_REG_6__2_ & n32305;
  assign n32451 = P1_P3_INSTQUEUE_REG_5__2_ & n32307;
  assign n32452 = P1_P3_INSTQUEUE_REG_4__2_ & n32309;
  assign n32453 = ~n32449 & ~n32450;
  assign n32454 = ~n32451 & n32453;
  assign n32455 = ~n32452 & n32454;
  assign n32456 = P1_P3_INSTQUEUE_REG_3__2_ & n32315;
  assign n32457 = P1_P3_INSTQUEUE_REG_2__2_ & n32317;
  assign n32458 = P1_P3_INSTQUEUE_REG_1__2_ & n32319;
  assign n32459 = P1_P3_INSTQUEUE_REG_0__2_ & n32321;
  assign n32460 = ~n32456 & ~n32457;
  assign n32461 = ~n32458 & n32460;
  assign n32462 = ~n32459 & n32461;
  assign n32463 = P1_P3_INSTQUEUE_REG_15__2_ & n32326;
  assign n32464 = P1_P3_INSTQUEUE_REG_14__2_ & n32328;
  assign n32465 = P1_P3_INSTQUEUE_REG_13__2_ & n32330;
  assign n32466 = P1_P3_INSTQUEUE_REG_12__2_ & n32332;
  assign n32467 = ~n32463 & ~n32464;
  assign n32468 = ~n32465 & n32467;
  assign n32469 = ~n32466 & n32468;
  assign n32470 = P1_P3_INSTQUEUE_REG_11__2_ & n32338;
  assign n32471 = P1_P3_INSTQUEUE_REG_10__2_ & n32340;
  assign n32472 = P1_P3_INSTQUEUE_REG_9__2_ & n32342;
  assign n32473 = P1_P3_INSTQUEUE_REG_8__2_ & n32344;
  assign n32474 = ~n32470 & ~n32471;
  assign n32475 = ~n32472 & n32474;
  assign n32476 = ~n32473 & n32475;
  assign n32477 = n32455 & n32462;
  assign n32478 = n32469 & n32477;
  assign n32479 = n32476 & n32478;
  assign n32480 = n32448 & n32479;
  assign n32481 = ~n32448 & ~n32479;
  assign n32482 = ~n32480 & ~n32481;
  assign n32483 = n31509 & ~n32482;
  assign n32484 = ~n32447 & ~n32483;
  assign n32485 = P1_P3_EAX_REG_23_ & P1_P3_EAX_REG_24_;
  assign n32486 = n32389 & n32485;
  assign n32487 = P1_P3_EAX_REG_25_ & ~n32486;
  assign n32488 = ~P1_P3_EAX_REG_25_ & n32486;
  assign n32489 = ~n32487 & ~n32488;
  assign n32490 = n31515 & ~n32489;
  assign n32491 = ~n32445 & ~n32446;
  assign n32492 = n32484 & n32491;
  assign n5066 = n32490 | ~n32492;
  assign n32494 = P1_BUF2_REG_26_ & n31960;
  assign n32495 = P1_BUF2_REG_10_ & n31962;
  assign n32496 = P1_P3_EAX_REG_26_ & ~n31508;
  assign n32497 = n32448 & ~n32479;
  assign n32498 = P1_P3_INSTQUEUE_REG_7__3_ & n32303;
  assign n32499 = P1_P3_INSTQUEUE_REG_6__3_ & n32305;
  assign n32500 = P1_P3_INSTQUEUE_REG_5__3_ & n32307;
  assign n32501 = P1_P3_INSTQUEUE_REG_4__3_ & n32309;
  assign n32502 = ~n32498 & ~n32499;
  assign n32503 = ~n32500 & n32502;
  assign n32504 = ~n32501 & n32503;
  assign n32505 = P1_P3_INSTQUEUE_REG_3__3_ & n32315;
  assign n32506 = P1_P3_INSTQUEUE_REG_2__3_ & n32317;
  assign n32507 = P1_P3_INSTQUEUE_REG_1__3_ & n32319;
  assign n32508 = P1_P3_INSTQUEUE_REG_0__3_ & n32321;
  assign n32509 = ~n32505 & ~n32506;
  assign n32510 = ~n32507 & n32509;
  assign n32511 = ~n32508 & n32510;
  assign n32512 = P1_P3_INSTQUEUE_REG_15__3_ & n32326;
  assign n32513 = P1_P3_INSTQUEUE_REG_14__3_ & n32328;
  assign n32514 = P1_P3_INSTQUEUE_REG_13__3_ & n32330;
  assign n32515 = P1_P3_INSTQUEUE_REG_12__3_ & n32332;
  assign n32516 = ~n32512 & ~n32513;
  assign n32517 = ~n32514 & n32516;
  assign n32518 = ~n32515 & n32517;
  assign n32519 = P1_P3_INSTQUEUE_REG_11__3_ & n32338;
  assign n32520 = P1_P3_INSTQUEUE_REG_10__3_ & n32340;
  assign n32521 = P1_P3_INSTQUEUE_REG_9__3_ & n32342;
  assign n32522 = P1_P3_INSTQUEUE_REG_8__3_ & n32344;
  assign n32523 = ~n32519 & ~n32520;
  assign n32524 = ~n32521 & n32523;
  assign n32525 = ~n32522 & n32524;
  assign n32526 = n32504 & n32511;
  assign n32527 = n32518 & n32526;
  assign n32528 = n32525 & n32527;
  assign n32529 = n32497 & n32528;
  assign n32530 = ~n32497 & ~n32528;
  assign n32531 = ~n32529 & ~n32530;
  assign n32532 = n31509 & ~n32531;
  assign n32533 = ~n32496 & ~n32532;
  assign n32534 = P1_P3_EAX_REG_25_ & n32486;
  assign n32535 = ~P1_P3_EAX_REG_26_ & n32534;
  assign n32536 = P1_P3_EAX_REG_26_ & ~n32534;
  assign n32537 = ~n32535 & ~n32536;
  assign n32538 = n31515 & ~n32537;
  assign n32539 = ~n32494 & ~n32495;
  assign n32540 = n32533 & n32539;
  assign n5071 = n32538 | ~n32540;
  assign n32542 = P1_BUF2_REG_27_ & n31960;
  assign n32543 = P1_BUF2_REG_11_ & n31962;
  assign n32544 = P1_P3_EAX_REG_27_ & ~n31508;
  assign n32545 = n32497 & ~n32528;
  assign n32546 = P1_P3_INSTQUEUE_REG_7__4_ & n32303;
  assign n32547 = P1_P3_INSTQUEUE_REG_6__4_ & n32305;
  assign n32548 = P1_P3_INSTQUEUE_REG_5__4_ & n32307;
  assign n32549 = P1_P3_INSTQUEUE_REG_4__4_ & n32309;
  assign n32550 = ~n32546 & ~n32547;
  assign n32551 = ~n32548 & n32550;
  assign n32552 = ~n32549 & n32551;
  assign n32553 = P1_P3_INSTQUEUE_REG_3__4_ & n32315;
  assign n32554 = P1_P3_INSTQUEUE_REG_2__4_ & n32317;
  assign n32555 = P1_P3_INSTQUEUE_REG_1__4_ & n32319;
  assign n32556 = P1_P3_INSTQUEUE_REG_0__4_ & n32321;
  assign n32557 = ~n32553 & ~n32554;
  assign n32558 = ~n32555 & n32557;
  assign n32559 = ~n32556 & n32558;
  assign n32560 = P1_P3_INSTQUEUE_REG_15__4_ & n32326;
  assign n32561 = P1_P3_INSTQUEUE_REG_14__4_ & n32328;
  assign n32562 = P1_P3_INSTQUEUE_REG_13__4_ & n32330;
  assign n32563 = P1_P3_INSTQUEUE_REG_12__4_ & n32332;
  assign n32564 = ~n32560 & ~n32561;
  assign n32565 = ~n32562 & n32564;
  assign n32566 = ~n32563 & n32565;
  assign n32567 = P1_P3_INSTQUEUE_REG_11__4_ & n32338;
  assign n32568 = P1_P3_INSTQUEUE_REG_10__4_ & n32340;
  assign n32569 = P1_P3_INSTQUEUE_REG_9__4_ & n32342;
  assign n32570 = P1_P3_INSTQUEUE_REG_8__4_ & n32344;
  assign n32571 = ~n32567 & ~n32568;
  assign n32572 = ~n32569 & n32571;
  assign n32573 = ~n32570 & n32572;
  assign n32574 = n32552 & n32559;
  assign n32575 = n32566 & n32574;
  assign n32576 = n32573 & n32575;
  assign n32577 = n32545 & n32576;
  assign n32578 = ~n32545 & ~n32576;
  assign n32579 = ~n32577 & ~n32578;
  assign n32580 = n31509 & ~n32579;
  assign n32581 = ~n32544 & ~n32580;
  assign n32582 = P1_P3_EAX_REG_25_ & P1_P3_EAX_REG_26_;
  assign n32583 = n32486 & n32582;
  assign n32584 = P1_P3_EAX_REG_27_ & ~n32583;
  assign n32585 = ~P1_P3_EAX_REG_27_ & n32583;
  assign n32586 = ~n32584 & ~n32585;
  assign n32587 = n31515 & ~n32586;
  assign n32588 = ~n32542 & ~n32543;
  assign n32589 = n32581 & n32588;
  assign n5076 = n32587 | ~n32589;
  assign n32591 = P1_BUF2_REG_28_ & n31960;
  assign n32592 = P1_BUF2_REG_12_ & n31962;
  assign n32593 = P1_P3_EAX_REG_28_ & ~n31508;
  assign n32594 = n32545 & ~n32576;
  assign n32595 = P1_P3_INSTQUEUE_REG_7__5_ & n32303;
  assign n32596 = P1_P3_INSTQUEUE_REG_6__5_ & n32305;
  assign n32597 = P1_P3_INSTQUEUE_REG_5__5_ & n32307;
  assign n32598 = P1_P3_INSTQUEUE_REG_4__5_ & n32309;
  assign n32599 = ~n32595 & ~n32596;
  assign n32600 = ~n32597 & n32599;
  assign n32601 = ~n32598 & n32600;
  assign n32602 = P1_P3_INSTQUEUE_REG_3__5_ & n32315;
  assign n32603 = P1_P3_INSTQUEUE_REG_2__5_ & n32317;
  assign n32604 = P1_P3_INSTQUEUE_REG_1__5_ & n32319;
  assign n32605 = P1_P3_INSTQUEUE_REG_0__5_ & n32321;
  assign n32606 = ~n32602 & ~n32603;
  assign n32607 = ~n32604 & n32606;
  assign n32608 = ~n32605 & n32607;
  assign n32609 = P1_P3_INSTQUEUE_REG_15__5_ & n32326;
  assign n32610 = P1_P3_INSTQUEUE_REG_14__5_ & n32328;
  assign n32611 = P1_P3_INSTQUEUE_REG_13__5_ & n32330;
  assign n32612 = P1_P3_INSTQUEUE_REG_12__5_ & n32332;
  assign n32613 = ~n32609 & ~n32610;
  assign n32614 = ~n32611 & n32613;
  assign n32615 = ~n32612 & n32614;
  assign n32616 = P1_P3_INSTQUEUE_REG_11__5_ & n32338;
  assign n32617 = P1_P3_INSTQUEUE_REG_10__5_ & n32340;
  assign n32618 = P1_P3_INSTQUEUE_REG_9__5_ & n32342;
  assign n32619 = P1_P3_INSTQUEUE_REG_8__5_ & n32344;
  assign n32620 = ~n32616 & ~n32617;
  assign n32621 = ~n32618 & n32620;
  assign n32622 = ~n32619 & n32621;
  assign n32623 = n32601 & n32608;
  assign n32624 = n32615 & n32623;
  assign n32625 = n32622 & n32624;
  assign n32626 = n32594 & n32625;
  assign n32627 = ~n32594 & ~n32625;
  assign n32628 = ~n32626 & ~n32627;
  assign n32629 = n31509 & ~n32628;
  assign n32630 = P1_P3_EAX_REG_27_ & n32583;
  assign n32631 = ~P1_P3_EAX_REG_28_ & n32630;
  assign n32632 = P1_P3_EAX_REG_28_ & ~n32630;
  assign n32633 = ~n32631 & ~n32632;
  assign n32634 = n31515 & ~n32633;
  assign n32635 = ~n32591 & ~n32592;
  assign n32636 = ~n32593 & n32635;
  assign n32637 = ~n32629 & n32636;
  assign n5081 = n32634 | ~n32637;
  assign n32639 = P1_BUF2_REG_29_ & n31960;
  assign n32640 = P1_BUF2_REG_13_ & n31962;
  assign n32641 = P1_P3_EAX_REG_29_ & ~n31508;
  assign n32642 = n32594 & ~n32625;
  assign n32643 = P1_P3_INSTQUEUE_REG_7__6_ & n32303;
  assign n32644 = P1_P3_INSTQUEUE_REG_6__6_ & n32305;
  assign n32645 = P1_P3_INSTQUEUE_REG_5__6_ & n32307;
  assign n32646 = P1_P3_INSTQUEUE_REG_4__6_ & n32309;
  assign n32647 = ~n32643 & ~n32644;
  assign n32648 = ~n32645 & n32647;
  assign n32649 = ~n32646 & n32648;
  assign n32650 = P1_P3_INSTQUEUE_REG_3__6_ & n32315;
  assign n32651 = P1_P3_INSTQUEUE_REG_2__6_ & n32317;
  assign n32652 = P1_P3_INSTQUEUE_REG_1__6_ & n32319;
  assign n32653 = P1_P3_INSTQUEUE_REG_0__6_ & n32321;
  assign n32654 = ~n32650 & ~n32651;
  assign n32655 = ~n32652 & n32654;
  assign n32656 = ~n32653 & n32655;
  assign n32657 = P1_P3_INSTQUEUE_REG_15__6_ & n32326;
  assign n32658 = P1_P3_INSTQUEUE_REG_14__6_ & n32328;
  assign n32659 = P1_P3_INSTQUEUE_REG_13__6_ & n32330;
  assign n32660 = P1_P3_INSTQUEUE_REG_12__6_ & n32332;
  assign n32661 = ~n32657 & ~n32658;
  assign n32662 = ~n32659 & n32661;
  assign n32663 = ~n32660 & n32662;
  assign n32664 = P1_P3_INSTQUEUE_REG_11__6_ & n32338;
  assign n32665 = P1_P3_INSTQUEUE_REG_10__6_ & n32340;
  assign n32666 = P1_P3_INSTQUEUE_REG_9__6_ & n32342;
  assign n32667 = P1_P3_INSTQUEUE_REG_8__6_ & n32344;
  assign n32668 = ~n32664 & ~n32665;
  assign n32669 = ~n32666 & n32668;
  assign n32670 = ~n32667 & n32669;
  assign n32671 = n32649 & n32656;
  assign n32672 = n32663 & n32671;
  assign n32673 = n32670 & n32672;
  assign n32674 = n32642 & n32673;
  assign n32675 = ~n32642 & ~n32673;
  assign n32676 = ~n32674 & ~n32675;
  assign n32677 = n31509 & ~n32676;
  assign n32678 = P1_P3_EAX_REG_27_ & P1_P3_EAX_REG_28_;
  assign n32679 = n32583 & n32678;
  assign n32680 = P1_P3_EAX_REG_29_ & ~n32679;
  assign n32681 = ~P1_P3_EAX_REG_29_ & n32679;
  assign n32682 = ~n32680 & ~n32681;
  assign n32683 = n31515 & ~n32682;
  assign n32684 = ~n32639 & ~n32640;
  assign n32685 = ~n32641 & n32684;
  assign n32686 = ~n32677 & n32685;
  assign n5086 = n32683 | ~n32686;
  assign n32688 = P1_BUF2_REG_30_ & n31960;
  assign n32689 = P1_BUF2_REG_14_ & n31962;
  assign n32690 = P1_P3_EAX_REG_30_ & ~n31508;
  assign n32691 = n32642 & ~n32673;
  assign n32692 = P1_P3_INSTQUEUE_REG_7__7_ & n32303;
  assign n32693 = P1_P3_INSTQUEUE_REG_6__7_ & n32305;
  assign n32694 = P1_P3_INSTQUEUE_REG_5__7_ & n32307;
  assign n32695 = P1_P3_INSTQUEUE_REG_4__7_ & n32309;
  assign n32696 = ~n32692 & ~n32693;
  assign n32697 = ~n32694 & n32696;
  assign n32698 = ~n32695 & n32697;
  assign n32699 = P1_P3_INSTQUEUE_REG_3__7_ & n32315;
  assign n32700 = P1_P3_INSTQUEUE_REG_2__7_ & n32317;
  assign n32701 = P1_P3_INSTQUEUE_REG_1__7_ & n32319;
  assign n32702 = P1_P3_INSTQUEUE_REG_0__7_ & n32321;
  assign n32703 = ~n32699 & ~n32700;
  assign n32704 = ~n32701 & n32703;
  assign n32705 = ~n32702 & n32704;
  assign n32706 = P1_P3_INSTQUEUE_REG_15__7_ & n32326;
  assign n32707 = P1_P3_INSTQUEUE_REG_14__7_ & n32328;
  assign n32708 = P1_P3_INSTQUEUE_REG_13__7_ & n32330;
  assign n32709 = P1_P3_INSTQUEUE_REG_12__7_ & n32332;
  assign n32710 = ~n32706 & ~n32707;
  assign n32711 = ~n32708 & n32710;
  assign n32712 = ~n32709 & n32711;
  assign n32713 = P1_P3_INSTQUEUE_REG_11__7_ & n32338;
  assign n32714 = P1_P3_INSTQUEUE_REG_10__7_ & n32340;
  assign n32715 = P1_P3_INSTQUEUE_REG_9__7_ & n32342;
  assign n32716 = P1_P3_INSTQUEUE_REG_8__7_ & n32344;
  assign n32717 = ~n32713 & ~n32714;
  assign n32718 = ~n32715 & n32717;
  assign n32719 = ~n32716 & n32718;
  assign n32720 = n32698 & n32705;
  assign n32721 = n32712 & n32720;
  assign n32722 = n32719 & n32721;
  assign n32723 = n32691 & n32722;
  assign n32724 = ~n32691 & ~n32722;
  assign n32725 = ~n32723 & ~n32724;
  assign n32726 = n31509 & ~n32725;
  assign n32727 = P1_P3_EAX_REG_29_ & n32679;
  assign n32728 = ~P1_P3_EAX_REG_30_ & n32727;
  assign n32729 = P1_P3_EAX_REG_30_ & ~n32727;
  assign n32730 = ~n32728 & ~n32729;
  assign n32731 = n31515 & ~n32730;
  assign n32732 = ~n32688 & ~n32689;
  assign n32733 = ~n32690 & n32732;
  assign n32734 = ~n32726 & n32733;
  assign n5091 = n32731 | ~n32734;
  assign n32736 = P1_P3_EAX_REG_31_ & ~n31508;
  assign n32737 = P1_BUF2_REG_31_ & n31960;
  assign n32738 = P1_P3_EAX_REG_30_ & n32727;
  assign n32739 = ~P1_P3_EAX_REG_31_ & n32738;
  assign n32740 = P1_P3_EAX_REG_31_ & ~n32738;
  assign n32741 = ~n32739 & ~n32740;
  assign n32742 = n31515 & ~n32741;
  assign n32743 = ~n32736 & ~n32737;
  assign n5096 = n32742 | ~n32743;
  assign n32745 = ~n25781 & ~n25875;
  assign n32746 = n25994 & ~n32745;
  assign n32747 = n25511 & n32746;
  assign n32748 = ~P1_P3_EBX_REG_0_ & n32747;
  assign n32749 = ~n25511 & n32746;
  assign n32750 = P1_P3_INSTQUEUE_REG_0__0_ & n32749;
  assign n32751 = P1_P3_EBX_REG_0_ & ~n32746;
  assign n32752 = ~n32748 & ~n32750;
  assign n5101 = n32751 | ~n32752;
  assign n32754 = ~P1_P3_EBX_REG_0_ & P1_P3_EBX_REG_1_;
  assign n32755 = P1_P3_EBX_REG_0_ & ~P1_P3_EBX_REG_1_;
  assign n32756 = ~n32754 & ~n32755;
  assign n32757 = n32747 & ~n32756;
  assign n32758 = P1_P3_INSTQUEUE_REG_0__1_ & n32749;
  assign n32759 = P1_P3_EBX_REG_1_ & ~n32746;
  assign n32760 = ~n32757 & ~n32758;
  assign n5106 = n32759 | ~n32760;
  assign n32762 = P1_P3_EBX_REG_0_ & P1_P3_EBX_REG_1_;
  assign n32763 = ~P1_P3_EBX_REG_2_ & n32762;
  assign n32764 = P1_P3_EBX_REG_2_ & ~n32762;
  assign n32765 = ~n32763 & ~n32764;
  assign n32766 = n32747 & ~n32765;
  assign n32767 = P1_P3_INSTQUEUE_REG_0__2_ & n32749;
  assign n32768 = P1_P3_EBX_REG_2_ & ~n32746;
  assign n32769 = ~n32766 & ~n32767;
  assign n5111 = n32768 | ~n32769;
  assign n32771 = P1_P3_EBX_REG_0_ & P1_P3_EBX_REG_2_;
  assign n32772 = P1_P3_EBX_REG_1_ & n32771;
  assign n32773 = P1_P3_EBX_REG_3_ & ~n32772;
  assign n32774 = ~P1_P3_EBX_REG_3_ & n32772;
  assign n32775 = ~n32773 & ~n32774;
  assign n32776 = n32747 & ~n32775;
  assign n32777 = P1_P3_INSTQUEUE_REG_0__3_ & n32749;
  assign n32778 = P1_P3_EBX_REG_3_ & ~n32746;
  assign n32779 = ~n32776 & ~n32777;
  assign n5116 = n32778 | ~n32779;
  assign n32781 = P1_P3_EBX_REG_3_ & n32772;
  assign n32782 = ~P1_P3_EBX_REG_4_ & n32781;
  assign n32783 = P1_P3_EBX_REG_4_ & ~n32781;
  assign n32784 = ~n32782 & ~n32783;
  assign n32785 = n32747 & ~n32784;
  assign n32786 = P1_P3_INSTQUEUE_REG_0__4_ & n32749;
  assign n32787 = P1_P3_EBX_REG_4_ & ~n32746;
  assign n32788 = ~n32785 & ~n32786;
  assign n5121 = n32787 | ~n32788;
  assign n32790 = P1_P3_EBX_REG_3_ & P1_P3_EBX_REG_4_;
  assign n32791 = n32772 & n32790;
  assign n32792 = P1_P3_EBX_REG_5_ & ~n32791;
  assign n32793 = ~P1_P3_EBX_REG_5_ & n32791;
  assign n32794 = ~n32792 & ~n32793;
  assign n32795 = n32747 & ~n32794;
  assign n32796 = P1_P3_INSTQUEUE_REG_0__5_ & n32749;
  assign n32797 = P1_P3_EBX_REG_5_ & ~n32746;
  assign n32798 = ~n32795 & ~n32796;
  assign n5126 = n32797 | ~n32798;
  assign n32800 = P1_P3_EBX_REG_5_ & n32791;
  assign n32801 = ~P1_P3_EBX_REG_6_ & n32800;
  assign n32802 = P1_P3_EBX_REG_6_ & ~n32800;
  assign n32803 = ~n32801 & ~n32802;
  assign n32804 = n32747 & ~n32803;
  assign n32805 = P1_P3_INSTQUEUE_REG_0__6_ & n32749;
  assign n32806 = P1_P3_EBX_REG_6_ & ~n32746;
  assign n32807 = ~n32804 & ~n32805;
  assign n5131 = n32806 | ~n32807;
  assign n32809 = P1_P3_EBX_REG_5_ & P1_P3_EBX_REG_6_;
  assign n32810 = n32791 & n32809;
  assign n32811 = P1_P3_EBX_REG_7_ & ~n32810;
  assign n32812 = ~P1_P3_EBX_REG_7_ & n32810;
  assign n32813 = ~n32811 & ~n32812;
  assign n32814 = n32747 & ~n32813;
  assign n32815 = P1_P3_INSTQUEUE_REG_0__7_ & n32749;
  assign n32816 = P1_P3_EBX_REG_7_ & ~n32746;
  assign n32817 = ~n32814 & ~n32815;
  assign n5136 = n32816 | ~n32817;
  assign n32819 = P1_P3_EBX_REG_7_ & n32810;
  assign n32820 = ~P1_P3_EBX_REG_8_ & n32819;
  assign n32821 = P1_P3_EBX_REG_8_ & ~n32819;
  assign n32822 = ~n32820 & ~n32821;
  assign n32823 = n32747 & ~n32822;
  assign n32824 = ~n31650 & n32749;
  assign n32825 = P1_P3_EBX_REG_8_ & ~n32746;
  assign n32826 = ~n32823 & ~n32824;
  assign n5141 = n32825 | ~n32826;
  assign n32828 = P1_P3_EBX_REG_7_ & P1_P3_EBX_REG_8_;
  assign n32829 = n32810 & n32828;
  assign n32830 = P1_P3_EBX_REG_9_ & ~n32829;
  assign n32831 = ~P1_P3_EBX_REG_9_ & n32829;
  assign n32832 = ~n32830 & ~n32831;
  assign n32833 = n32747 & ~n32832;
  assign n32834 = ~n31692 & n32749;
  assign n32835 = P1_P3_EBX_REG_9_ & ~n32746;
  assign n32836 = ~n32833 & ~n32834;
  assign n5146 = n32835 | ~n32836;
  assign n32838 = P1_P3_EBX_REG_10_ & ~n32746;
  assign n32839 = ~n31735 & n32749;
  assign n32840 = P1_P3_EBX_REG_9_ & n32829;
  assign n32841 = ~P1_P3_EBX_REG_10_ & n32840;
  assign n32842 = P1_P3_EBX_REG_10_ & ~n32840;
  assign n32843 = ~n32841 & ~n32842;
  assign n32844 = n32747 & ~n32843;
  assign n32845 = ~n32838 & ~n32839;
  assign n5151 = n32844 | ~n32845;
  assign n32847 = P1_P3_EBX_REG_11_ & ~n32746;
  assign n32848 = ~n31777 & n32749;
  assign n32849 = P1_P3_EBX_REG_9_ & P1_P3_EBX_REG_10_;
  assign n32850 = n32829 & n32849;
  assign n32851 = P1_P3_EBX_REG_11_ & ~n32850;
  assign n32852 = ~P1_P3_EBX_REG_11_ & n32850;
  assign n32853 = ~n32851 & ~n32852;
  assign n32854 = n32747 & ~n32853;
  assign n32855 = ~n32847 & ~n32848;
  assign n5156 = n32854 | ~n32855;
  assign n32857 = P1_P3_EBX_REG_12_ & ~n32746;
  assign n32858 = ~n31820 & n32749;
  assign n32859 = P1_P3_EBX_REG_11_ & n32850;
  assign n32860 = ~P1_P3_EBX_REG_12_ & n32859;
  assign n32861 = P1_P3_EBX_REG_12_ & ~n32859;
  assign n32862 = ~n32860 & ~n32861;
  assign n32863 = n32747 & ~n32862;
  assign n32864 = ~n32857 & ~n32858;
  assign n5161 = n32863 | ~n32864;
  assign n32866 = P1_P3_EBX_REG_13_ & ~n32746;
  assign n32867 = ~n31863 & n32749;
  assign n32868 = P1_P3_EBX_REG_11_ & P1_P3_EBX_REG_12_;
  assign n32869 = n32850 & n32868;
  assign n32870 = P1_P3_EBX_REG_13_ & ~n32869;
  assign n32871 = ~P1_P3_EBX_REG_13_ & n32869;
  assign n32872 = ~n32870 & ~n32871;
  assign n32873 = n32747 & ~n32872;
  assign n32874 = ~n32866 & ~n32867;
  assign n5166 = n32873 | ~n32874;
  assign n32876 = P1_P3_EBX_REG_14_ & ~n32746;
  assign n32877 = ~n31906 & n32749;
  assign n32878 = P1_P3_EBX_REG_13_ & n32869;
  assign n32879 = ~P1_P3_EBX_REG_14_ & n32878;
  assign n32880 = P1_P3_EBX_REG_14_ & ~n32878;
  assign n32881 = ~n32879 & ~n32880;
  assign n32882 = n32747 & ~n32881;
  assign n32883 = ~n32876 & ~n32877;
  assign n5171 = n32882 | ~n32883;
  assign n32885 = P1_P3_EBX_REG_15_ & ~n32746;
  assign n32886 = ~n31948 & n32749;
  assign n32887 = P1_P3_EBX_REG_13_ & P1_P3_EBX_REG_14_;
  assign n32888 = n32869 & n32887;
  assign n32889 = P1_P3_EBX_REG_15_ & ~n32888;
  assign n32890 = ~P1_P3_EBX_REG_15_ & n32888;
  assign n32891 = ~n32889 & ~n32890;
  assign n32892 = n32747 & ~n32891;
  assign n32893 = ~n32885 & ~n32886;
  assign n5176 = n32892 | ~n32893;
  assign n32895 = P1_P3_EBX_REG_16_ & ~n32746;
  assign n32896 = ~n32020 & n32749;
  assign n32897 = P1_P3_EBX_REG_15_ & n32888;
  assign n32898 = ~P1_P3_EBX_REG_16_ & n32897;
  assign n32899 = P1_P3_EBX_REG_16_ & ~n32897;
  assign n32900 = ~n32898 & ~n32899;
  assign n32901 = n32747 & ~n32900;
  assign n32902 = ~n32895 & ~n32896;
  assign n5181 = n32901 | ~n32902;
  assign n32904 = P1_P3_EBX_REG_17_ & ~n32746;
  assign n32905 = ~n32064 & n32749;
  assign n32906 = P1_P3_EBX_REG_15_ & P1_P3_EBX_REG_16_;
  assign n32907 = n32888 & n32906;
  assign n32908 = P1_P3_EBX_REG_17_ & ~n32907;
  assign n32909 = ~P1_P3_EBX_REG_17_ & n32907;
  assign n32910 = ~n32908 & ~n32909;
  assign n32911 = n32747 & ~n32910;
  assign n32912 = ~n32904 & ~n32905;
  assign n5186 = n32911 | ~n32912;
  assign n32914 = P1_P3_EBX_REG_18_ & ~n32746;
  assign n32915 = ~n32109 & n32749;
  assign n32916 = P1_P3_EBX_REG_17_ & n32907;
  assign n32917 = ~P1_P3_EBX_REG_18_ & n32916;
  assign n32918 = P1_P3_EBX_REG_18_ & ~n32916;
  assign n32919 = ~n32917 & ~n32918;
  assign n32920 = n32747 & ~n32919;
  assign n32921 = ~n32914 & ~n32915;
  assign n5191 = n32920 | ~n32921;
  assign n32923 = P1_P3_EBX_REG_19_ & ~n32746;
  assign n32924 = ~n32153 & n32749;
  assign n32925 = P1_P3_EBX_REG_17_ & P1_P3_EBX_REG_18_;
  assign n32926 = n32907 & n32925;
  assign n32927 = P1_P3_EBX_REG_19_ & ~n32926;
  assign n32928 = ~P1_P3_EBX_REG_19_ & n32926;
  assign n32929 = ~n32927 & ~n32928;
  assign n32930 = n32747 & ~n32929;
  assign n32931 = ~n32923 & ~n32924;
  assign n5196 = n32930 | ~n32931;
  assign n32933 = P1_P3_EBX_REG_20_ & ~n32746;
  assign n32934 = ~n32198 & n32749;
  assign n32935 = P1_P3_EBX_REG_19_ & n32926;
  assign n32936 = ~P1_P3_EBX_REG_20_ & n32935;
  assign n32937 = P1_P3_EBX_REG_20_ & ~n32935;
  assign n32938 = ~n32936 & ~n32937;
  assign n32939 = n32747 & ~n32938;
  assign n32940 = ~n32933 & ~n32934;
  assign n5201 = n32939 | ~n32940;
  assign n32942 = P1_P3_EBX_REG_21_ & ~n32746;
  assign n32943 = ~n32242 & n32749;
  assign n32944 = P1_P3_EBX_REG_19_ & P1_P3_EBX_REG_20_;
  assign n32945 = n32926 & n32944;
  assign n32946 = P1_P3_EBX_REG_21_ & ~n32945;
  assign n32947 = ~P1_P3_EBX_REG_21_ & n32945;
  assign n32948 = ~n32946 & ~n32947;
  assign n32949 = n32747 & ~n32948;
  assign n32950 = ~n32942 & ~n32943;
  assign n5206 = n32949 | ~n32950;
  assign n32952 = P1_P3_EBX_REG_22_ & ~n32746;
  assign n32953 = ~n32287 & n32749;
  assign n32954 = P1_P3_EBX_REG_21_ & n32945;
  assign n32955 = ~P1_P3_EBX_REG_22_ & n32954;
  assign n32956 = P1_P3_EBX_REG_22_ & ~n32954;
  assign n32957 = ~n32955 & ~n32956;
  assign n32958 = n32747 & ~n32957;
  assign n32959 = ~n32952 & ~n32953;
  assign n5211 = n32958 | ~n32959;
  assign n32961 = P1_P3_EBX_REG_23_ & ~n32746;
  assign n32962 = ~n32385 & n32749;
  assign n32963 = P1_P3_EBX_REG_21_ & P1_P3_EBX_REG_22_;
  assign n32964 = n32945 & n32963;
  assign n32965 = P1_P3_EBX_REG_23_ & ~n32964;
  assign n32966 = ~P1_P3_EBX_REG_23_ & n32964;
  assign n32967 = ~n32965 & ~n32966;
  assign n32968 = n32747 & ~n32967;
  assign n32969 = ~n32961 & ~n32962;
  assign n5216 = n32968 | ~n32969;
  assign n32971 = P1_P3_EBX_REG_24_ & ~n32746;
  assign n32972 = ~n32434 & n32749;
  assign n32973 = P1_P3_EBX_REG_23_ & n32964;
  assign n32974 = ~P1_P3_EBX_REG_24_ & n32973;
  assign n32975 = P1_P3_EBX_REG_24_ & ~n32973;
  assign n32976 = ~n32974 & ~n32975;
  assign n32977 = n32747 & ~n32976;
  assign n32978 = ~n32971 & ~n32972;
  assign n5221 = n32977 | ~n32978;
  assign n32980 = P1_P3_EBX_REG_25_ & ~n32746;
  assign n32981 = ~n32482 & n32749;
  assign n32982 = P1_P3_EBX_REG_23_ & P1_P3_EBX_REG_24_;
  assign n32983 = n32964 & n32982;
  assign n32984 = P1_P3_EBX_REG_25_ & ~n32983;
  assign n32985 = ~P1_P3_EBX_REG_25_ & n32983;
  assign n32986 = ~n32984 & ~n32985;
  assign n32987 = n32747 & ~n32986;
  assign n32988 = ~n32980 & ~n32981;
  assign n5226 = n32987 | ~n32988;
  assign n32990 = P1_P3_EBX_REG_26_ & ~n32746;
  assign n32991 = ~n32531 & n32749;
  assign n32992 = P1_P3_EBX_REG_25_ & n32983;
  assign n32993 = ~P1_P3_EBX_REG_26_ & n32992;
  assign n32994 = P1_P3_EBX_REG_26_ & ~n32992;
  assign n32995 = ~n32993 & ~n32994;
  assign n32996 = n32747 & ~n32995;
  assign n32997 = ~n32990 & ~n32991;
  assign n5231 = n32996 | ~n32997;
  assign n32999 = P1_P3_EBX_REG_27_ & ~n32746;
  assign n33000 = ~n32579 & n32749;
  assign n33001 = P1_P3_EBX_REG_25_ & P1_P3_EBX_REG_26_;
  assign n33002 = n32983 & n33001;
  assign n33003 = P1_P3_EBX_REG_27_ & ~n33002;
  assign n33004 = ~P1_P3_EBX_REG_27_ & n33002;
  assign n33005 = ~n33003 & ~n33004;
  assign n33006 = n32747 & ~n33005;
  assign n33007 = ~n32999 & ~n33000;
  assign n5236 = n33006 | ~n33007;
  assign n33009 = P1_P3_EBX_REG_28_ & ~n32746;
  assign n33010 = ~n32628 & n32749;
  assign n33011 = P1_P3_EBX_REG_27_ & n33002;
  assign n33012 = ~P1_P3_EBX_REG_28_ & n33011;
  assign n33013 = P1_P3_EBX_REG_28_ & ~n33011;
  assign n33014 = ~n33012 & ~n33013;
  assign n33015 = n32747 & ~n33014;
  assign n33016 = ~n33009 & ~n33010;
  assign n5241 = n33015 | ~n33016;
  assign n33018 = P1_P3_EBX_REG_29_ & ~n32746;
  assign n33019 = ~n32676 & n32749;
  assign n33020 = P1_P3_EBX_REG_27_ & P1_P3_EBX_REG_28_;
  assign n33021 = n33002 & n33020;
  assign n33022 = P1_P3_EBX_REG_29_ & ~n33021;
  assign n33023 = ~P1_P3_EBX_REG_29_ & n33021;
  assign n33024 = ~n33022 & ~n33023;
  assign n33025 = n32747 & ~n33024;
  assign n33026 = ~n33018 & ~n33019;
  assign n5246 = n33025 | ~n33026;
  assign n33028 = P1_P3_EBX_REG_30_ & ~n32746;
  assign n33029 = ~n32725 & n32749;
  assign n33030 = P1_P3_EBX_REG_29_ & n33021;
  assign n33031 = ~P1_P3_EBX_REG_30_ & n33030;
  assign n33032 = P1_P3_EBX_REG_30_ & ~n33030;
  assign n33033 = ~n33031 & ~n33032;
  assign n33034 = n32747 & ~n33033;
  assign n33035 = ~n33028 & ~n33029;
  assign n5251 = n33034 | ~n33035;
  assign n33037 = P1_P3_EBX_REG_31_ & ~n32746;
  assign n33038 = P1_P3_EBX_REG_30_ & n33030;
  assign n33039 = ~P1_P3_EBX_REG_31_ & n33038;
  assign n33040 = P1_P3_EBX_REG_31_ & ~n33038;
  assign n33041 = ~n33039 & ~n33040;
  assign n33042 = n32747 & ~n33041;
  assign n5256 = n33037 | n33042;
  assign n33044 = ~n26005 & ~n26044;
  assign n33045 = ~n27608 & n33044;
  assign n33046 = n25872 & n25880;
  assign n33047 = n25994 & ~n33046;
  assign n33048 = n33045 & ~n33047;
  assign n33049 = P1_P3_STATE2_REG_2_ & ~n33048;
  assign n33050 = n25722 & n33049;
  assign n33051 = ~n25355 & n33050;
  assign n33052 = ~P1_P3_EBX_REG_31_ & n33051;
  assign n33053 = n25640 & n33049;
  assign n33054 = ~n25358 & n33053;
  assign n33055 = n25358 & n33053;
  assign n33056 = ~n25355 & n33055;
  assign n33057 = ~n33052 & ~n33054;
  assign n33058 = ~n33056 & n33057;
  assign n33059 = P1_P3_EBX_REG_0_ & ~n33058;
  assign n33060 = n25355 & n33055;
  assign n33061 = P1_P3_REIP_REG_0_ & n33060;
  assign n33062 = P1_P3_EBX_REG_31_ & n33051;
  assign n33063 = P1_P3_EBX_REG_0_ & n33062;
  assign n33064 = n25717 & n33049;
  assign n33065 = ~P1_P3_INSTQUEUERD_ADDR_REG_0_ & n33064;
  assign n33066 = n25713 & n33049;
  assign n33067 = ~P1_P3_INSTQUEUERD_ADDR_REG_0_ & n33066;
  assign n33068 = ~n33065 & ~n33067;
  assign n33069 = ~n33061 & ~n33063;
  assign n33070 = n33068 & n33069;
  assign n33071 = n25355 & n33050;
  assign n33072 = P1_P3_REIP_REG_0_ & n33071;
  assign n33073 = P1_P3_STATE2_REG_1_ & ~n33048;
  assign n33074 = n31185 & n33073;
  assign n33075 = P1_P3_PHYADDRPOINTER_REG_0_ & n33074;
  assign n33076 = P1_P3_REIP_REG_0_ & n33048;
  assign n33077 = P1_P3_STATE2_REG_3_ & ~n33048;
  assign n33078 = P1_P3_PHYADDRPOINTER_REG_0_ & n33077;
  assign n33079 = ~n33076 & ~n33078;
  assign n33080 = ~n31185 & n33073;
  assign n33081 = P1_P3_PHYADDRPOINTER_REG_0_ & n33080;
  assign n33082 = n33079 & ~n33081;
  assign n33083 = ~n33059 & n33070;
  assign n33084 = ~n33072 & n33083;
  assign n33085 = ~n33075 & n33084;
  assign n5261 = ~n33082 | ~n33085;
  assign n33087 = P1_P3_EBX_REG_1_ & ~n33058;
  assign n33088 = ~P1_P3_REIP_REG_1_ & n33060;
  assign n33089 = ~n32756 & n33062;
  assign n33090 = ~n25364 & ~n25369;
  assign n33091 = n33064 & ~n33090;
  assign n33092 = n33066 & ~n33090;
  assign n33093 = ~n33091 & ~n33092;
  assign n33094 = ~n33088 & ~n33089;
  assign n33095 = n33093 & n33094;
  assign n33096 = ~P1_P3_REIP_REG_1_ & n33071;
  assign n33097 = ~P1_P3_PHYADDRPOINTER_REG_1_ & n33074;
  assign n33098 = P1_P3_REIP_REG_1_ & n33048;
  assign n33099 = P1_P3_PHYADDRPOINTER_REG_1_ & n33077;
  assign n33100 = ~n33098 & ~n33099;
  assign n33101 = P1_P3_PHYADDRPOINTER_REG_0_ & P1_P3_PHYADDRPOINTER_REG_1_;
  assign n33102 = ~P1_P3_PHYADDRPOINTER_REG_0_ & ~P1_P3_PHYADDRPOINTER_REG_1_;
  assign n33103 = ~n33101 & ~n33102;
  assign n33104 = n33080 & ~n33103;
  assign n33105 = n33100 & ~n33104;
  assign n33106 = ~n33087 & n33095;
  assign n33107 = ~n33096 & n33106;
  assign n33108 = ~n33097 & n33107;
  assign n5266 = ~n33105 | ~n33108;
  assign n33110 = P1_P3_EBX_REG_2_ & ~n33058;
  assign n33111 = P1_P3_REIP_REG_1_ & ~P1_P3_REIP_REG_2_;
  assign n33112 = ~P1_P3_REIP_REG_1_ & P1_P3_REIP_REG_2_;
  assign n33113 = ~n33111 & ~n33112;
  assign n33114 = n33060 & ~n33113;
  assign n33115 = ~P1_P3_EBX_REG_0_ & ~P1_P3_EBX_REG_1_;
  assign n33116 = P1_P3_EBX_REG_2_ & ~n33115;
  assign n33117 = ~P1_P3_EBX_REG_2_ & n33115;
  assign n33118 = ~n33116 & ~n33117;
  assign n33119 = n33062 & n33118;
  assign n33120 = ~n25842 & n33064;
  assign n33121 = ~n25842 & n33066;
  assign n33122 = ~n33120 & ~n33121;
  assign n33123 = ~n33114 & ~n33119;
  assign n33124 = n33122 & n33123;
  assign n33125 = n33071 & ~n33113;
  assign n33126 = ~n30519 & n33074;
  assign n33127 = P1_P3_REIP_REG_2_ & n33048;
  assign n33128 = P1_P3_PHYADDRPOINTER_REG_2_ & n33077;
  assign n33129 = ~n33127 & ~n33128;
  assign n33130 = ~P1_P3_PHYADDRPOINTER_REG_0_ & P1_P3_PHYADDRPOINTER_REG_1_;
  assign n33131 = ~n30519 & ~n33130;
  assign n33132 = n30519 & n33130;
  assign n33133 = ~n33131 & ~n33132;
  assign n33134 = n33080 & n33133;
  assign n33135 = n33129 & ~n33134;
  assign n33136 = ~n33110 & n33124;
  assign n33137 = ~n33125 & n33136;
  assign n33138 = ~n33126 & n33137;
  assign n5271 = ~n33135 | ~n33138;
  assign n33140 = P1_P3_EBX_REG_3_ & ~n33058;
  assign n33141 = P1_P3_REIP_REG_1_ & P1_P3_REIP_REG_2_;
  assign n33142 = ~P1_P3_REIP_REG_3_ & n33141;
  assign n33143 = P1_P3_REIP_REG_3_ & ~n33141;
  assign n33144 = ~n33142 & ~n33143;
  assign n33145 = n33060 & ~n33144;
  assign n33146 = ~P1_P3_EBX_REG_3_ & n33117;
  assign n33147 = P1_P3_EBX_REG_3_ & ~n33117;
  assign n33148 = ~n33146 & ~n33147;
  assign n33149 = n33062 & n33148;
  assign n33150 = ~P1_P3_INSTQUEUERD_ADDR_REG_3_ & n25890;
  assign n33151 = ~n25891 & ~n33150;
  assign n33152 = n33064 & ~n33151;
  assign n33153 = n33066 & ~n33151;
  assign n33154 = ~n33152 & ~n33153;
  assign n33155 = ~n33145 & ~n33149;
  assign n33156 = n33154 & n33155;
  assign n33157 = n33071 & ~n33144;
  assign n33158 = ~n30541 & n33074;
  assign n33159 = P1_P3_REIP_REG_3_ & n33048;
  assign n33160 = P1_P3_PHYADDRPOINTER_REG_3_ & n33077;
  assign n33161 = ~n33159 & ~n33160;
  assign n33162 = n30541 & n33132;
  assign n33163 = ~n30541 & ~n33132;
  assign n33164 = ~n33162 & ~n33163;
  assign n33165 = n33080 & n33164;
  assign n33166 = n33161 & ~n33165;
  assign n33167 = ~n33140 & n33156;
  assign n33168 = ~n33157 & n33167;
  assign n33169 = ~n33158 & n33168;
  assign n5276 = ~n33166 | ~n33169;
  assign n33171 = P1_P3_INSTQUEUERD_ADDR_REG_3_ & n25890;
  assign n33172 = ~P1_P3_INSTQUEUERD_ADDR_REG_4_ & n33171;
  assign n33173 = P1_P3_INSTQUEUERD_ADDR_REG_4_ & ~n33171;
  assign n33174 = ~n33172 & ~n33173;
  assign n33175 = n33066 & ~n33174;
  assign n33176 = n33064 & ~n33174;
  assign n33177 = ~n33175 & ~n33176;
  assign n33178 = P1_P3_EBX_REG_4_ & ~n33058;
  assign n33179 = P1_P3_EBX_REG_4_ & ~n33146;
  assign n33180 = ~P1_P3_EBX_REG_3_ & ~P1_P3_EBX_REG_4_;
  assign n33181 = n33117 & n33180;
  assign n33182 = ~n33179 & ~n33181;
  assign n33183 = n33062 & n33182;
  assign n33184 = n27607 & ~n33048;
  assign n33185 = P1_P3_REIP_REG_3_ & n33141;
  assign n33186 = ~P1_P3_REIP_REG_4_ & n33185;
  assign n33187 = P1_P3_REIP_REG_4_ & ~n33185;
  assign n33188 = ~n33186 & ~n33187;
  assign n33189 = n33060 & ~n33188;
  assign n33190 = ~n33183 & ~n33184;
  assign n33191 = ~n33189 & n33190;
  assign n33192 = n33071 & ~n33188;
  assign n33193 = ~n30562 & n33074;
  assign n33194 = n33177 & ~n33178;
  assign n33195 = n33191 & n33194;
  assign n33196 = ~n33192 & n33195;
  assign n33197 = ~n33193 & n33196;
  assign n33198 = P1_P3_REIP_REG_4_ & n33048;
  assign n33199 = P1_P3_PHYADDRPOINTER_REG_4_ & n33077;
  assign n33200 = ~n33198 & ~n33199;
  assign n33201 = ~n30562 & ~n33162;
  assign n33202 = n30541 & n30562;
  assign n33203 = n33132 & n33202;
  assign n33204 = ~n33201 & ~n33203;
  assign n33205 = n33080 & n33204;
  assign n33206 = n33200 & ~n33205;
  assign n5281 = ~n33197 | ~n33206;
  assign n33208 = P1_P3_INSTQUEUERD_ADDR_REG_4_ & n33171;
  assign n33209 = n33066 & n33208;
  assign n33210 = n33064 & n33208;
  assign n33211 = ~n33209 & ~n33210;
  assign n33212 = P1_P3_EBX_REG_5_ & ~n33058;
  assign n33213 = ~P1_P3_EBX_REG_5_ & n33181;
  assign n33214 = P1_P3_EBX_REG_5_ & ~n33181;
  assign n33215 = ~n33213 & ~n33214;
  assign n33216 = n33062 & n33215;
  assign n33217 = P1_P3_REIP_REG_4_ & n33185;
  assign n33218 = ~P1_P3_REIP_REG_5_ & n33217;
  assign n33219 = P1_P3_REIP_REG_5_ & ~n33217;
  assign n33220 = ~n33218 & ~n33219;
  assign n33221 = n33060 & ~n33220;
  assign n33222 = ~n33184 & ~n33216;
  assign n33223 = ~n33221 & n33222;
  assign n33224 = n33071 & ~n33220;
  assign n33225 = ~n30585 & n33074;
  assign n33226 = n33211 & ~n33212;
  assign n33227 = n33223 & n33226;
  assign n33228 = ~n33224 & n33227;
  assign n33229 = ~n33225 & n33228;
  assign n33230 = P1_P3_REIP_REG_5_ & n33048;
  assign n33231 = P1_P3_PHYADDRPOINTER_REG_5_ & n33077;
  assign n33232 = ~n33230 & ~n33231;
  assign n33233 = n30585 & n33203;
  assign n33234 = ~n30585 & ~n33203;
  assign n33235 = ~n33233 & ~n33234;
  assign n33236 = n33080 & n33235;
  assign n33237 = n33232 & ~n33236;
  assign n5286 = ~n33229 | ~n33237;
  assign n33239 = P1_P3_REIP_REG_5_ & n33217;
  assign n33240 = ~P1_P3_REIP_REG_6_ & n33239;
  assign n33241 = P1_P3_REIP_REG_6_ & ~n33239;
  assign n33242 = ~n33240 & ~n33241;
  assign n33243 = n33071 & ~n33242;
  assign n33244 = P1_P3_EBX_REG_6_ & ~n33058;
  assign n33245 = P1_P3_EBX_REG_6_ & ~n33213;
  assign n33246 = ~P1_P3_EBX_REG_5_ & ~P1_P3_EBX_REG_6_;
  assign n33247 = n33181 & n33246;
  assign n33248 = ~n33245 & ~n33247;
  assign n33249 = n33062 & n33248;
  assign n33250 = n33060 & ~n33242;
  assign n33251 = ~n33184 & ~n33249;
  assign n33252 = ~n33250 & n33251;
  assign n33253 = ~n30608 & ~n33233;
  assign n33254 = n30585 & n30608;
  assign n33255 = n33203 & n33254;
  assign n33256 = ~n33253 & ~n33255;
  assign n33257 = n33080 & n33256;
  assign n33258 = P1_P3_REIP_REG_6_ & n33048;
  assign n33259 = P1_P3_PHYADDRPOINTER_REG_6_ & n33077;
  assign n33260 = ~n33258 & ~n33259;
  assign n33261 = ~n30608 & n33074;
  assign n33262 = n33260 & ~n33261;
  assign n33263 = ~n33243 & ~n33244;
  assign n33264 = n33252 & n33263;
  assign n33265 = ~n33257 & n33264;
  assign n5291 = ~n33262 | ~n33265;
  assign n33267 = P1_P3_REIP_REG_6_ & n33239;
  assign n33268 = ~P1_P3_REIP_REG_7_ & n33267;
  assign n33269 = P1_P3_REIP_REG_7_ & ~n33267;
  assign n33270 = ~n33268 & ~n33269;
  assign n33271 = n33071 & ~n33270;
  assign n33272 = P1_P3_EBX_REG_7_ & ~n33058;
  assign n33273 = ~P1_P3_EBX_REG_7_ & n33247;
  assign n33274 = P1_P3_EBX_REG_7_ & ~n33247;
  assign n33275 = ~n33273 & ~n33274;
  assign n33276 = n33062 & n33275;
  assign n33277 = n33060 & ~n33270;
  assign n33278 = ~n33184 & ~n33276;
  assign n33279 = ~n33277 & n33278;
  assign n33280 = n30631 & n33255;
  assign n33281 = ~n30631 & ~n33255;
  assign n33282 = ~n33280 & ~n33281;
  assign n33283 = n33080 & n33282;
  assign n33284 = P1_P3_REIP_REG_7_ & n33048;
  assign n33285 = P1_P3_PHYADDRPOINTER_REG_7_ & n33077;
  assign n33286 = ~n33284 & ~n33285;
  assign n33287 = ~n30631 & n33074;
  assign n33288 = n33286 & ~n33287;
  assign n33289 = ~n33271 & ~n33272;
  assign n33290 = n33279 & n33289;
  assign n33291 = ~n33283 & n33290;
  assign n5296 = ~n33288 | ~n33291;
  assign n33293 = P1_P3_REIP_REG_7_ & n33267;
  assign n33294 = ~P1_P3_REIP_REG_8_ & n33293;
  assign n33295 = P1_P3_REIP_REG_8_ & ~n33293;
  assign n33296 = ~n33294 & ~n33295;
  assign n33297 = n33071 & ~n33296;
  assign n33298 = P1_P3_EBX_REG_8_ & ~n33058;
  assign n33299 = P1_P3_EBX_REG_8_ & ~n33273;
  assign n33300 = ~P1_P3_EBX_REG_7_ & ~P1_P3_EBX_REG_8_;
  assign n33301 = n33247 & n33300;
  assign n33302 = ~n33299 & ~n33301;
  assign n33303 = n33062 & n33302;
  assign n33304 = n33060 & ~n33296;
  assign n33305 = ~n33184 & ~n33303;
  assign n33306 = ~n33304 & n33305;
  assign n33307 = ~n30654 & ~n33280;
  assign n33308 = n30631 & n30654;
  assign n33309 = n33255 & n33308;
  assign n33310 = ~n33307 & ~n33309;
  assign n33311 = n33080 & n33310;
  assign n33312 = P1_P3_REIP_REG_8_ & n33048;
  assign n33313 = P1_P3_PHYADDRPOINTER_REG_8_ & n33077;
  assign n33314 = ~n33312 & ~n33313;
  assign n33315 = ~n30654 & n33074;
  assign n33316 = n33314 & ~n33315;
  assign n33317 = ~n33297 & ~n33298;
  assign n33318 = n33306 & n33317;
  assign n33319 = ~n33311 & n33318;
  assign n5301 = ~n33316 | ~n33319;
  assign n33321 = P1_P3_REIP_REG_8_ & n33293;
  assign n33322 = ~P1_P3_REIP_REG_9_ & n33321;
  assign n33323 = P1_P3_REIP_REG_9_ & ~n33321;
  assign n33324 = ~n33322 & ~n33323;
  assign n33325 = n33071 & ~n33324;
  assign n33326 = P1_P3_EBX_REG_9_ & ~n33058;
  assign n33327 = ~P1_P3_EBX_REG_9_ & n33301;
  assign n33328 = P1_P3_EBX_REG_9_ & ~n33301;
  assign n33329 = ~n33327 & ~n33328;
  assign n33330 = n33062 & n33329;
  assign n33331 = n33060 & ~n33324;
  assign n33332 = ~n33184 & ~n33330;
  assign n33333 = ~n33331 & n33332;
  assign n33334 = n30677 & n33309;
  assign n33335 = ~n30677 & ~n33309;
  assign n33336 = ~n33334 & ~n33335;
  assign n33337 = n33080 & n33336;
  assign n33338 = P1_P3_REIP_REG_9_ & n33048;
  assign n33339 = P1_P3_PHYADDRPOINTER_REG_9_ & n33077;
  assign n33340 = ~n33338 & ~n33339;
  assign n33341 = ~n30677 & n33074;
  assign n33342 = n33340 & ~n33341;
  assign n33343 = ~n33325 & ~n33326;
  assign n33344 = n33333 & n33343;
  assign n33345 = ~n33337 & n33344;
  assign n5306 = ~n33342 | ~n33345;
  assign n33347 = P1_P3_REIP_REG_9_ & n33321;
  assign n33348 = ~P1_P3_REIP_REG_10_ & n33347;
  assign n33349 = P1_P3_REIP_REG_10_ & ~n33347;
  assign n33350 = ~n33348 & ~n33349;
  assign n33351 = n33071 & ~n33350;
  assign n33352 = P1_P3_EBX_REG_10_ & ~n33058;
  assign n33353 = P1_P3_EBX_REG_10_ & ~n33327;
  assign n33354 = ~P1_P3_EBX_REG_9_ & ~P1_P3_EBX_REG_10_;
  assign n33355 = n33301 & n33354;
  assign n33356 = ~n33353 & ~n33355;
  assign n33357 = n33062 & n33356;
  assign n33358 = n33060 & ~n33350;
  assign n33359 = ~n33184 & ~n33357;
  assign n33360 = ~n33358 & n33359;
  assign n33361 = ~n30700 & ~n33334;
  assign n33362 = n30677 & n30700;
  assign n33363 = n33309 & n33362;
  assign n33364 = ~n33361 & ~n33363;
  assign n33365 = n33080 & n33364;
  assign n33366 = P1_P3_REIP_REG_10_ & n33048;
  assign n33367 = P1_P3_PHYADDRPOINTER_REG_10_ & n33077;
  assign n33368 = ~n33366 & ~n33367;
  assign n33369 = ~n30700 & n33074;
  assign n33370 = n33368 & ~n33369;
  assign n33371 = ~n33351 & ~n33352;
  assign n33372 = n33360 & n33371;
  assign n33373 = ~n33365 & n33372;
  assign n5311 = ~n33370 | ~n33373;
  assign n33375 = P1_P3_REIP_REG_10_ & n33347;
  assign n33376 = ~P1_P3_REIP_REG_11_ & n33375;
  assign n33377 = P1_P3_REIP_REG_11_ & ~n33375;
  assign n33378 = ~n33376 & ~n33377;
  assign n33379 = n33071 & ~n33378;
  assign n33380 = P1_P3_EBX_REG_11_ & ~n33058;
  assign n33381 = ~P1_P3_EBX_REG_11_ & n33355;
  assign n33382 = P1_P3_EBX_REG_11_ & ~n33355;
  assign n33383 = ~n33381 & ~n33382;
  assign n33384 = n33062 & n33383;
  assign n33385 = n33060 & ~n33378;
  assign n33386 = ~n33184 & ~n33384;
  assign n33387 = ~n33385 & n33386;
  assign n33388 = n30723 & n33363;
  assign n33389 = ~n30723 & ~n33363;
  assign n33390 = ~n33388 & ~n33389;
  assign n33391 = n33080 & n33390;
  assign n33392 = P1_P3_REIP_REG_11_ & n33048;
  assign n33393 = P1_P3_PHYADDRPOINTER_REG_11_ & n33077;
  assign n33394 = ~n33392 & ~n33393;
  assign n33395 = ~n30723 & n33074;
  assign n33396 = n33394 & ~n33395;
  assign n33397 = ~n33379 & ~n33380;
  assign n33398 = n33387 & n33397;
  assign n33399 = ~n33391 & n33398;
  assign n5316 = ~n33396 | ~n33399;
  assign n33401 = P1_P3_REIP_REG_11_ & n33375;
  assign n33402 = ~P1_P3_REIP_REG_12_ & n33401;
  assign n33403 = P1_P3_REIP_REG_12_ & ~n33401;
  assign n33404 = ~n33402 & ~n33403;
  assign n33405 = n33071 & ~n33404;
  assign n33406 = P1_P3_EBX_REG_12_ & ~n33058;
  assign n33407 = P1_P3_EBX_REG_12_ & ~n33381;
  assign n33408 = ~P1_P3_EBX_REG_11_ & ~P1_P3_EBX_REG_12_;
  assign n33409 = n33355 & n33408;
  assign n33410 = ~n33407 & ~n33409;
  assign n33411 = n33062 & n33410;
  assign n33412 = n33060 & ~n33404;
  assign n33413 = ~n33184 & ~n33411;
  assign n33414 = ~n33412 & n33413;
  assign n33415 = ~n30746 & ~n33388;
  assign n33416 = n30723 & n30746;
  assign n33417 = n33363 & n33416;
  assign n33418 = ~n33415 & ~n33417;
  assign n33419 = n33080 & n33418;
  assign n33420 = P1_P3_REIP_REG_12_ & n33048;
  assign n33421 = P1_P3_PHYADDRPOINTER_REG_12_ & n33077;
  assign n33422 = ~n33420 & ~n33421;
  assign n33423 = ~n30746 & n33074;
  assign n33424 = n33422 & ~n33423;
  assign n33425 = ~n33405 & ~n33406;
  assign n33426 = n33414 & n33425;
  assign n33427 = ~n33419 & n33426;
  assign n5321 = ~n33424 | ~n33427;
  assign n33429 = P1_P3_REIP_REG_12_ & n33401;
  assign n33430 = ~P1_P3_REIP_REG_13_ & n33429;
  assign n33431 = P1_P3_REIP_REG_13_ & ~n33429;
  assign n33432 = ~n33430 & ~n33431;
  assign n33433 = n33071 & ~n33432;
  assign n33434 = P1_P3_EBX_REG_13_ & ~n33058;
  assign n33435 = ~P1_P3_EBX_REG_13_ & n33409;
  assign n33436 = P1_P3_EBX_REG_13_ & ~n33409;
  assign n33437 = ~n33435 & ~n33436;
  assign n33438 = n33062 & n33437;
  assign n33439 = n33060 & ~n33432;
  assign n33440 = ~n33184 & ~n33438;
  assign n33441 = ~n33439 & n33440;
  assign n33442 = n30769 & n33417;
  assign n33443 = ~n30769 & ~n33417;
  assign n33444 = ~n33442 & ~n33443;
  assign n33445 = n33080 & n33444;
  assign n33446 = P1_P3_REIP_REG_13_ & n33048;
  assign n33447 = P1_P3_PHYADDRPOINTER_REG_13_ & n33077;
  assign n33448 = ~n33446 & ~n33447;
  assign n33449 = ~n30769 & n33074;
  assign n33450 = n33448 & ~n33449;
  assign n33451 = ~n33433 & ~n33434;
  assign n33452 = n33441 & n33451;
  assign n33453 = ~n33445 & n33452;
  assign n5326 = ~n33450 | ~n33453;
  assign n33455 = P1_P3_REIP_REG_13_ & n33429;
  assign n33456 = ~P1_P3_REIP_REG_14_ & n33455;
  assign n33457 = P1_P3_REIP_REG_14_ & ~n33455;
  assign n33458 = ~n33456 & ~n33457;
  assign n33459 = n33071 & ~n33458;
  assign n33460 = P1_P3_EBX_REG_14_ & ~n33058;
  assign n33461 = P1_P3_EBX_REG_14_ & ~n33435;
  assign n33462 = ~P1_P3_EBX_REG_13_ & ~P1_P3_EBX_REG_14_;
  assign n33463 = n33409 & n33462;
  assign n33464 = ~n33461 & ~n33463;
  assign n33465 = n33062 & n33464;
  assign n33466 = n33060 & ~n33458;
  assign n33467 = ~n33184 & ~n33465;
  assign n33468 = ~n33466 & n33467;
  assign n33469 = ~n30792 & ~n33442;
  assign n33470 = n30769 & n30792;
  assign n33471 = n33417 & n33470;
  assign n33472 = ~n33469 & ~n33471;
  assign n33473 = n33080 & n33472;
  assign n33474 = P1_P3_REIP_REG_14_ & n33048;
  assign n33475 = P1_P3_PHYADDRPOINTER_REG_14_ & n33077;
  assign n33476 = ~n33474 & ~n33475;
  assign n33477 = ~n30792 & n33074;
  assign n33478 = n33476 & ~n33477;
  assign n33479 = ~n33459 & ~n33460;
  assign n33480 = n33468 & n33479;
  assign n33481 = ~n33473 & n33480;
  assign n5331 = ~n33478 | ~n33481;
  assign n33483 = P1_P3_REIP_REG_14_ & n33455;
  assign n33484 = ~P1_P3_REIP_REG_15_ & n33483;
  assign n33485 = P1_P3_REIP_REG_15_ & ~n33483;
  assign n33486 = ~n33484 & ~n33485;
  assign n33487 = n33071 & ~n33486;
  assign n33488 = P1_P3_EBX_REG_15_ & ~n33058;
  assign n33489 = ~P1_P3_EBX_REG_15_ & n33463;
  assign n33490 = P1_P3_EBX_REG_15_ & ~n33463;
  assign n33491 = ~n33489 & ~n33490;
  assign n33492 = n33062 & n33491;
  assign n33493 = n33060 & ~n33486;
  assign n33494 = ~n33184 & ~n33492;
  assign n33495 = ~n33493 & n33494;
  assign n33496 = n30815 & n33471;
  assign n33497 = ~n30815 & ~n33471;
  assign n33498 = ~n33496 & ~n33497;
  assign n33499 = n33080 & n33498;
  assign n33500 = P1_P3_REIP_REG_15_ & n33048;
  assign n33501 = P1_P3_PHYADDRPOINTER_REG_15_ & n33077;
  assign n33502 = ~n33500 & ~n33501;
  assign n33503 = ~n30815 & n33074;
  assign n33504 = n33502 & ~n33503;
  assign n33505 = ~n33487 & ~n33488;
  assign n33506 = n33495 & n33505;
  assign n33507 = ~n33499 & n33506;
  assign n5336 = ~n33504 | ~n33507;
  assign n33509 = P1_P3_REIP_REG_15_ & n33483;
  assign n33510 = ~P1_P3_REIP_REG_16_ & n33509;
  assign n33511 = P1_P3_REIP_REG_16_ & ~n33509;
  assign n33512 = ~n33510 & ~n33511;
  assign n33513 = n33071 & ~n33512;
  assign n33514 = P1_P3_EBX_REG_16_ & ~n33058;
  assign n33515 = P1_P3_EBX_REG_16_ & ~n33489;
  assign n33516 = ~P1_P3_EBX_REG_15_ & ~P1_P3_EBX_REG_16_;
  assign n33517 = n33463 & n33516;
  assign n33518 = ~n33515 & ~n33517;
  assign n33519 = n33062 & n33518;
  assign n33520 = n33060 & ~n33512;
  assign n33521 = ~n33184 & ~n33519;
  assign n33522 = ~n33520 & n33521;
  assign n33523 = ~n30838 & ~n33496;
  assign n33524 = n30815 & n30838;
  assign n33525 = n33471 & n33524;
  assign n33526 = ~n33523 & ~n33525;
  assign n33527 = n33080 & n33526;
  assign n33528 = P1_P3_REIP_REG_16_ & n33048;
  assign n33529 = P1_P3_PHYADDRPOINTER_REG_16_ & n33077;
  assign n33530 = ~n33528 & ~n33529;
  assign n33531 = ~n30838 & n33074;
  assign n33532 = n33530 & ~n33531;
  assign n33533 = ~n33513 & ~n33514;
  assign n33534 = n33522 & n33533;
  assign n33535 = ~n33527 & n33534;
  assign n5341 = ~n33532 | ~n33535;
  assign n33537 = P1_P3_REIP_REG_16_ & n33509;
  assign n33538 = ~P1_P3_REIP_REG_17_ & n33537;
  assign n33539 = P1_P3_REIP_REG_17_ & ~n33537;
  assign n33540 = ~n33538 & ~n33539;
  assign n33541 = n33071 & ~n33540;
  assign n33542 = P1_P3_EBX_REG_17_ & ~n33058;
  assign n33543 = ~P1_P3_EBX_REG_17_ & n33517;
  assign n33544 = P1_P3_EBX_REG_17_ & ~n33517;
  assign n33545 = ~n33543 & ~n33544;
  assign n33546 = n33062 & n33545;
  assign n33547 = n33060 & ~n33540;
  assign n33548 = ~n33184 & ~n33546;
  assign n33549 = ~n33547 & n33548;
  assign n33550 = n30861 & n33525;
  assign n33551 = ~n30861 & ~n33525;
  assign n33552 = ~n33550 & ~n33551;
  assign n33553 = n33080 & n33552;
  assign n33554 = P1_P3_REIP_REG_17_ & n33048;
  assign n33555 = P1_P3_PHYADDRPOINTER_REG_17_ & n33077;
  assign n33556 = ~n33554 & ~n33555;
  assign n33557 = ~n30861 & n33074;
  assign n33558 = n33556 & ~n33557;
  assign n33559 = ~n33541 & ~n33542;
  assign n33560 = n33549 & n33559;
  assign n33561 = ~n33553 & n33560;
  assign n5346 = ~n33558 | ~n33561;
  assign n33563 = P1_P3_REIP_REG_17_ & n33537;
  assign n33564 = ~P1_P3_REIP_REG_18_ & n33563;
  assign n33565 = P1_P3_REIP_REG_18_ & ~n33563;
  assign n33566 = ~n33564 & ~n33565;
  assign n33567 = n33071 & ~n33566;
  assign n33568 = P1_P3_EBX_REG_18_ & ~n33058;
  assign n33569 = P1_P3_EBX_REG_18_ & ~n33543;
  assign n33570 = ~P1_P3_EBX_REG_17_ & ~P1_P3_EBX_REG_18_;
  assign n33571 = n33517 & n33570;
  assign n33572 = ~n33569 & ~n33571;
  assign n33573 = n33062 & n33572;
  assign n33574 = n33060 & ~n33566;
  assign n33575 = ~n33184 & ~n33573;
  assign n33576 = ~n33574 & n33575;
  assign n33577 = ~n30884 & ~n33550;
  assign n33578 = n30861 & n30884;
  assign n33579 = n33525 & n33578;
  assign n33580 = ~n33577 & ~n33579;
  assign n33581 = n33080 & n33580;
  assign n33582 = P1_P3_REIP_REG_18_ & n33048;
  assign n33583 = P1_P3_PHYADDRPOINTER_REG_18_ & n33077;
  assign n33584 = ~n33582 & ~n33583;
  assign n33585 = ~n30884 & n33074;
  assign n33586 = n33584 & ~n33585;
  assign n33587 = ~n33567 & ~n33568;
  assign n33588 = n33576 & n33587;
  assign n33589 = ~n33581 & n33588;
  assign n5351 = ~n33586 | ~n33589;
  assign n33591 = P1_P3_REIP_REG_18_ & n33563;
  assign n33592 = ~P1_P3_REIP_REG_19_ & n33591;
  assign n33593 = P1_P3_REIP_REG_19_ & ~n33591;
  assign n33594 = ~n33592 & ~n33593;
  assign n33595 = n33071 & ~n33594;
  assign n33596 = P1_P3_EBX_REG_19_ & ~n33058;
  assign n33597 = ~P1_P3_EBX_REG_19_ & n33571;
  assign n33598 = P1_P3_EBX_REG_19_ & ~n33571;
  assign n33599 = ~n33597 & ~n33598;
  assign n33600 = n33062 & n33599;
  assign n33601 = n33060 & ~n33594;
  assign n33602 = ~n33184 & ~n33600;
  assign n33603 = ~n33601 & n33602;
  assign n33604 = n30907 & n33579;
  assign n33605 = ~n30907 & ~n33579;
  assign n33606 = ~n33604 & ~n33605;
  assign n33607 = n33080 & n33606;
  assign n33608 = P1_P3_REIP_REG_19_ & n33048;
  assign n33609 = P1_P3_PHYADDRPOINTER_REG_19_ & n33077;
  assign n33610 = ~n33608 & ~n33609;
  assign n33611 = ~n30907 & n33074;
  assign n33612 = n33610 & ~n33611;
  assign n33613 = ~n33595 & ~n33596;
  assign n33614 = n33603 & n33613;
  assign n33615 = ~n33607 & n33614;
  assign n5356 = ~n33612 | ~n33615;
  assign n33617 = P1_P3_REIP_REG_19_ & n33591;
  assign n33618 = ~P1_P3_REIP_REG_20_ & n33617;
  assign n33619 = P1_P3_REIP_REG_20_ & ~n33617;
  assign n33620 = ~n33618 & ~n33619;
  assign n33621 = n33071 & ~n33620;
  assign n33622 = P1_P3_EBX_REG_20_ & ~n33058;
  assign n33623 = n33060 & ~n33620;
  assign n33624 = P1_P3_EBX_REG_20_ & ~n33597;
  assign n33625 = ~P1_P3_EBX_REG_19_ & ~P1_P3_EBX_REG_20_;
  assign n33626 = n33571 & n33625;
  assign n33627 = ~n33624 & ~n33626;
  assign n33628 = n33062 & n33627;
  assign n33629 = ~n33623 & ~n33628;
  assign n33630 = ~n30930 & ~n33604;
  assign n33631 = n30907 & n30930;
  assign n33632 = n33579 & n33631;
  assign n33633 = ~n33630 & ~n33632;
  assign n33634 = n33080 & n33633;
  assign n33635 = P1_P3_REIP_REG_20_ & n33048;
  assign n33636 = P1_P3_PHYADDRPOINTER_REG_20_ & n33077;
  assign n33637 = ~n33635 & ~n33636;
  assign n33638 = ~n30930 & n33074;
  assign n33639 = n33637 & ~n33638;
  assign n33640 = ~n33621 & ~n33622;
  assign n33641 = n33629 & n33640;
  assign n33642 = ~n33634 & n33641;
  assign n5361 = ~n33639 | ~n33642;
  assign n33644 = P1_P3_REIP_REG_20_ & n33617;
  assign n33645 = ~P1_P3_REIP_REG_21_ & n33644;
  assign n33646 = P1_P3_REIP_REG_21_ & ~n33644;
  assign n33647 = ~n33645 & ~n33646;
  assign n33648 = n33071 & ~n33647;
  assign n33649 = P1_P3_EBX_REG_21_ & ~n33058;
  assign n33650 = n33060 & ~n33647;
  assign n33651 = ~P1_P3_EBX_REG_21_ & n33626;
  assign n33652 = P1_P3_EBX_REG_21_ & ~n33626;
  assign n33653 = ~n33651 & ~n33652;
  assign n33654 = n33062 & n33653;
  assign n33655 = ~n33650 & ~n33654;
  assign n33656 = n30953 & n33632;
  assign n33657 = ~n30953 & ~n33632;
  assign n33658 = ~n33656 & ~n33657;
  assign n33659 = n33080 & n33658;
  assign n33660 = P1_P3_REIP_REG_21_ & n33048;
  assign n33661 = P1_P3_PHYADDRPOINTER_REG_21_ & n33077;
  assign n33662 = ~n33660 & ~n33661;
  assign n33663 = ~n30953 & n33074;
  assign n33664 = n33662 & ~n33663;
  assign n33665 = ~n33648 & ~n33649;
  assign n33666 = n33655 & n33665;
  assign n33667 = ~n33659 & n33666;
  assign n5366 = ~n33664 | ~n33667;
  assign n33669 = P1_P3_REIP_REG_21_ & n33644;
  assign n33670 = ~P1_P3_REIP_REG_22_ & n33669;
  assign n33671 = P1_P3_REIP_REG_22_ & ~n33669;
  assign n33672 = ~n33670 & ~n33671;
  assign n33673 = n33071 & ~n33672;
  assign n33674 = P1_P3_EBX_REG_22_ & ~n33058;
  assign n33675 = n33060 & ~n33672;
  assign n33676 = P1_P3_EBX_REG_22_ & ~n33651;
  assign n33677 = ~P1_P3_EBX_REG_21_ & ~P1_P3_EBX_REG_22_;
  assign n33678 = n33626 & n33677;
  assign n33679 = ~n33676 & ~n33678;
  assign n33680 = n33062 & n33679;
  assign n33681 = ~n33675 & ~n33680;
  assign n33682 = ~n30976 & ~n33656;
  assign n33683 = n30953 & n30976;
  assign n33684 = n33632 & n33683;
  assign n33685 = ~n33682 & ~n33684;
  assign n33686 = n33080 & n33685;
  assign n33687 = P1_P3_REIP_REG_22_ & n33048;
  assign n33688 = P1_P3_PHYADDRPOINTER_REG_22_ & n33077;
  assign n33689 = ~n33687 & ~n33688;
  assign n33690 = ~n30976 & n33074;
  assign n33691 = n33689 & ~n33690;
  assign n33692 = ~n33673 & ~n33674;
  assign n33693 = n33681 & n33692;
  assign n33694 = ~n33686 & n33693;
  assign n5371 = ~n33691 | ~n33694;
  assign n33696 = P1_P3_REIP_REG_22_ & n33669;
  assign n33697 = ~P1_P3_REIP_REG_23_ & n33696;
  assign n33698 = P1_P3_REIP_REG_23_ & ~n33696;
  assign n33699 = ~n33697 & ~n33698;
  assign n33700 = n33071 & ~n33699;
  assign n33701 = P1_P3_EBX_REG_23_ & ~n33058;
  assign n33702 = n33060 & ~n33699;
  assign n33703 = ~P1_P3_EBX_REG_23_ & n33678;
  assign n33704 = P1_P3_EBX_REG_23_ & ~n33678;
  assign n33705 = ~n33703 & ~n33704;
  assign n33706 = n33062 & n33705;
  assign n33707 = ~n33702 & ~n33706;
  assign n33708 = n30999 & n33684;
  assign n33709 = ~n30999 & ~n33684;
  assign n33710 = ~n33708 & ~n33709;
  assign n33711 = n33080 & n33710;
  assign n33712 = P1_P3_REIP_REG_23_ & n33048;
  assign n33713 = P1_P3_PHYADDRPOINTER_REG_23_ & n33077;
  assign n33714 = ~n33712 & ~n33713;
  assign n33715 = ~n30999 & n33074;
  assign n33716 = n33714 & ~n33715;
  assign n33717 = ~n33700 & ~n33701;
  assign n33718 = n33707 & n33717;
  assign n33719 = ~n33711 & n33718;
  assign n5376 = ~n33716 | ~n33719;
  assign n33721 = P1_P3_REIP_REG_23_ & n33696;
  assign n33722 = ~P1_P3_REIP_REG_24_ & n33721;
  assign n33723 = P1_P3_REIP_REG_24_ & ~n33721;
  assign n33724 = ~n33722 & ~n33723;
  assign n33725 = n33071 & ~n33724;
  assign n33726 = P1_P3_EBX_REG_24_ & ~n33058;
  assign n33727 = n33060 & ~n33724;
  assign n33728 = P1_P3_EBX_REG_24_ & ~n33703;
  assign n33729 = ~P1_P3_EBX_REG_23_ & ~P1_P3_EBX_REG_24_;
  assign n33730 = n33678 & n33729;
  assign n33731 = ~n33728 & ~n33730;
  assign n33732 = n33062 & n33731;
  assign n33733 = ~n33727 & ~n33732;
  assign n33734 = ~n31023 & ~n33708;
  assign n33735 = n30999 & n31023;
  assign n33736 = n33684 & n33735;
  assign n33737 = ~n33734 & ~n33736;
  assign n33738 = n33080 & n33737;
  assign n33739 = P1_P3_REIP_REG_24_ & n33048;
  assign n33740 = P1_P3_PHYADDRPOINTER_REG_24_ & n33077;
  assign n33741 = ~n33739 & ~n33740;
  assign n33742 = ~n31023 & n33074;
  assign n33743 = n33741 & ~n33742;
  assign n33744 = ~n33725 & ~n33726;
  assign n33745 = n33733 & n33744;
  assign n33746 = ~n33738 & n33745;
  assign n5381 = ~n33743 | ~n33746;
  assign n33748 = P1_P3_REIP_REG_24_ & n33721;
  assign n33749 = ~P1_P3_REIP_REG_25_ & n33748;
  assign n33750 = P1_P3_REIP_REG_25_ & ~n33748;
  assign n33751 = ~n33749 & ~n33750;
  assign n33752 = n33071 & ~n33751;
  assign n33753 = P1_P3_EBX_REG_25_ & ~n33058;
  assign n33754 = n33060 & ~n33751;
  assign n33755 = ~P1_P3_EBX_REG_25_ & n33730;
  assign n33756 = P1_P3_EBX_REG_25_ & ~n33730;
  assign n33757 = ~n33755 & ~n33756;
  assign n33758 = n33062 & n33757;
  assign n33759 = ~n33754 & ~n33758;
  assign n33760 = n31046 & n33736;
  assign n33761 = ~n31046 & ~n33736;
  assign n33762 = ~n33760 & ~n33761;
  assign n33763 = n33080 & n33762;
  assign n33764 = P1_P3_REIP_REG_25_ & n33048;
  assign n33765 = P1_P3_PHYADDRPOINTER_REG_25_ & n33077;
  assign n33766 = ~n33764 & ~n33765;
  assign n33767 = ~n31046 & n33074;
  assign n33768 = n33766 & ~n33767;
  assign n33769 = ~n33752 & ~n33753;
  assign n33770 = n33759 & n33769;
  assign n33771 = ~n33763 & n33770;
  assign n5386 = ~n33768 | ~n33771;
  assign n33773 = P1_P3_REIP_REG_25_ & n33748;
  assign n33774 = ~P1_P3_REIP_REG_26_ & n33773;
  assign n33775 = P1_P3_REIP_REG_26_ & ~n33773;
  assign n33776 = ~n33774 & ~n33775;
  assign n33777 = n33071 & ~n33776;
  assign n33778 = P1_P3_EBX_REG_26_ & ~n33058;
  assign n33779 = n33060 & ~n33776;
  assign n33780 = P1_P3_EBX_REG_26_ & ~n33755;
  assign n33781 = ~P1_P3_EBX_REG_25_ & ~P1_P3_EBX_REG_26_;
  assign n33782 = n33730 & n33781;
  assign n33783 = ~n33780 & ~n33782;
  assign n33784 = n33062 & n33783;
  assign n33785 = ~n33779 & ~n33784;
  assign n33786 = ~n31069 & ~n33760;
  assign n33787 = n31046 & n31069;
  assign n33788 = n33736 & n33787;
  assign n33789 = ~n33786 & ~n33788;
  assign n33790 = n33080 & n33789;
  assign n33791 = P1_P3_REIP_REG_26_ & n33048;
  assign n33792 = P1_P3_PHYADDRPOINTER_REG_26_ & n33077;
  assign n33793 = ~n33791 & ~n33792;
  assign n33794 = ~n31069 & n33074;
  assign n33795 = n33793 & ~n33794;
  assign n33796 = ~n33777 & ~n33778;
  assign n33797 = n33785 & n33796;
  assign n33798 = ~n33790 & n33797;
  assign n5391 = ~n33795 | ~n33798;
  assign n33800 = P1_P3_REIP_REG_26_ & n33773;
  assign n33801 = ~P1_P3_REIP_REG_27_ & n33800;
  assign n33802 = P1_P3_REIP_REG_27_ & ~n33800;
  assign n33803 = ~n33801 & ~n33802;
  assign n33804 = n33071 & ~n33803;
  assign n33805 = P1_P3_EBX_REG_27_ & ~n33058;
  assign n33806 = n33060 & ~n33803;
  assign n33807 = ~P1_P3_EBX_REG_27_ & n33782;
  assign n33808 = P1_P3_EBX_REG_27_ & ~n33782;
  assign n33809 = ~n33807 & ~n33808;
  assign n33810 = n33062 & n33809;
  assign n33811 = ~n33806 & ~n33810;
  assign n33812 = n31092 & n33788;
  assign n33813 = ~n31092 & ~n33788;
  assign n33814 = ~n33812 & ~n33813;
  assign n33815 = n33080 & n33814;
  assign n33816 = P1_P3_REIP_REG_27_ & n33048;
  assign n33817 = P1_P3_PHYADDRPOINTER_REG_27_ & n33077;
  assign n33818 = ~n33816 & ~n33817;
  assign n33819 = ~n31092 & n33074;
  assign n33820 = n33818 & ~n33819;
  assign n33821 = ~n33804 & ~n33805;
  assign n33822 = n33811 & n33821;
  assign n33823 = ~n33815 & n33822;
  assign n5396 = ~n33820 | ~n33823;
  assign n33825 = P1_P3_REIP_REG_27_ & n33800;
  assign n33826 = ~P1_P3_REIP_REG_28_ & n33825;
  assign n33827 = P1_P3_REIP_REG_28_ & ~n33825;
  assign n33828 = ~n33826 & ~n33827;
  assign n33829 = n33071 & ~n33828;
  assign n33830 = P1_P3_EBX_REG_28_ & ~n33058;
  assign n33831 = n33060 & ~n33828;
  assign n33832 = P1_P3_EBX_REG_28_ & ~n33807;
  assign n33833 = ~P1_P3_EBX_REG_27_ & ~P1_P3_EBX_REG_28_;
  assign n33834 = n33782 & n33833;
  assign n33835 = ~n33832 & ~n33834;
  assign n33836 = n33062 & n33835;
  assign n33837 = ~n33831 & ~n33836;
  assign n33838 = ~n31116 & ~n33812;
  assign n33839 = n31092 & n31116;
  assign n33840 = n33788 & n33839;
  assign n33841 = ~n33838 & ~n33840;
  assign n33842 = n33080 & n33841;
  assign n33843 = P1_P3_REIP_REG_28_ & n33048;
  assign n33844 = P1_P3_PHYADDRPOINTER_REG_28_ & n33077;
  assign n33845 = ~n33843 & ~n33844;
  assign n33846 = ~n31116 & n33074;
  assign n33847 = n33845 & ~n33846;
  assign n33848 = ~n33829 & ~n33830;
  assign n33849 = n33837 & n33848;
  assign n33850 = ~n33842 & n33849;
  assign n5401 = ~n33847 | ~n33850;
  assign n33852 = P1_P3_REIP_REG_28_ & n33825;
  assign n33853 = ~P1_P3_REIP_REG_29_ & n33852;
  assign n33854 = P1_P3_REIP_REG_29_ & ~n33852;
  assign n33855 = ~n33853 & ~n33854;
  assign n33856 = n33071 & ~n33855;
  assign n33857 = P1_P3_EBX_REG_29_ & ~n33058;
  assign n33858 = n33060 & ~n33855;
  assign n33859 = P1_P3_EBX_REG_29_ & ~n33834;
  assign n33860 = ~P1_P3_EBX_REG_29_ & n33834;
  assign n33861 = ~n33859 & ~n33860;
  assign n33862 = n33062 & n33861;
  assign n33863 = ~n33858 & ~n33862;
  assign n33864 = ~n31139 & ~n33840;
  assign n33865 = n31139 & n33840;
  assign n33866 = ~n33864 & ~n33865;
  assign n33867 = n33080 & n33866;
  assign n33868 = P1_P3_REIP_REG_29_ & n33048;
  assign n33869 = P1_P3_PHYADDRPOINTER_REG_29_ & n33077;
  assign n33870 = ~n33868 & ~n33869;
  assign n33871 = ~n31139 & n33074;
  assign n33872 = n33870 & ~n33871;
  assign n33873 = ~n33856 & ~n33857;
  assign n33874 = n33863 & n33873;
  assign n33875 = ~n33867 & n33874;
  assign n5406 = ~n33872 | ~n33875;
  assign n33877 = P1_P3_REIP_REG_29_ & n33852;
  assign n33878 = ~P1_P3_REIP_REG_30_ & n33877;
  assign n33879 = P1_P3_REIP_REG_30_ & ~n33877;
  assign n33880 = ~n33878 & ~n33879;
  assign n33881 = n33071 & ~n33880;
  assign n33882 = P1_P3_EBX_REG_30_ & ~n33058;
  assign n33883 = n33060 & ~n33880;
  assign n33884 = ~P1_P3_EBX_REG_30_ & n33860;
  assign n33885 = P1_P3_EBX_REG_30_ & ~n33860;
  assign n33886 = ~n33884 & ~n33885;
  assign n33887 = n33062 & n33886;
  assign n33888 = ~n33883 & ~n33887;
  assign n33889 = n31162 & n33865;
  assign n33890 = ~n31162 & ~n33865;
  assign n33891 = ~n33889 & ~n33890;
  assign n33892 = n33080 & n33891;
  assign n33893 = P1_P3_REIP_REG_30_ & n33048;
  assign n33894 = P1_P3_PHYADDRPOINTER_REG_30_ & n33077;
  assign n33895 = ~n33893 & ~n33894;
  assign n33896 = ~n31162 & n33074;
  assign n33897 = n33895 & ~n33896;
  assign n33898 = ~n33881 & ~n33882;
  assign n33899 = n33888 & n33898;
  assign n33900 = ~n33892 & n33899;
  assign n5411 = ~n33897 | ~n33900;
  assign n33902 = ~n31185 & n33889;
  assign n33903 = n31185 & ~n33889;
  assign n33904 = ~n33902 & ~n33903;
  assign n33905 = ~n31185 & n33074;
  assign n33906 = n33904 & ~n33905;
  assign n33907 = P1_P3_EBX_REG_31_ & ~n33058;
  assign n33908 = P1_P3_EBX_REG_31_ & n33884;
  assign n33909 = ~P1_P3_EBX_REG_31_ & ~n33884;
  assign n33910 = ~n33908 & ~n33909;
  assign n33911 = n33062 & ~n33910;
  assign n33912 = P1_P3_REIP_REG_30_ & n33877;
  assign n33913 = ~P1_P3_REIP_REG_31_ & n33912;
  assign n33914 = P1_P3_REIP_REG_31_ & ~n33912;
  assign n33915 = ~n33913 & ~n33914;
  assign n33916 = n33060 & ~n33915;
  assign n33917 = P1_P3_PHYADDRPOINTER_REG_31_ & n33077;
  assign n33918 = P1_P3_REIP_REG_31_ & n33048;
  assign n33919 = ~n33917 & ~n33918;
  assign n33920 = n33071 & ~n33915;
  assign n33921 = n33919 & ~n33920;
  assign n33922 = ~n33907 & ~n33911;
  assign n33923 = ~n33916 & n33922;
  assign n33924 = n33921 & n33923;
  assign n33925 = n33906 & n33924;
  assign n33926 = ~n33080 & ~n33905;
  assign n33927 = n33924 & n33926;
  assign n5416 = ~n33925 & ~n33927;
  assign n33929 = ~P1_P3_DATAWIDTH_REG_1_ & ~P1_P3_REIP_REG_1_;
  assign n33930 = ~P1_P3_DATAWIDTH_REG_30_ & ~P1_P3_DATAWIDTH_REG_31_;
  assign n33931 = P1_P3_DATAWIDTH_REG_0_ & P1_P3_DATAWIDTH_REG_1_;
  assign n33932 = ~P1_P3_DATAWIDTH_REG_28_ & ~P1_P3_DATAWIDTH_REG_29_;
  assign n33933 = ~P1_P3_DATAWIDTH_REG_26_ & ~P1_P3_DATAWIDTH_REG_27_;
  assign n33934 = n33930 & ~n33931;
  assign n33935 = n33932 & n33934;
  assign n33936 = n33933 & n33935;
  assign n33937 = ~P1_P3_DATAWIDTH_REG_22_ & ~P1_P3_DATAWIDTH_REG_23_;
  assign n33938 = ~P1_P3_DATAWIDTH_REG_24_ & n33937;
  assign n33939 = ~P1_P3_DATAWIDTH_REG_25_ & n33938;
  assign n33940 = ~P1_P3_DATAWIDTH_REG_18_ & ~P1_P3_DATAWIDTH_REG_19_;
  assign n33941 = ~P1_P3_DATAWIDTH_REG_20_ & n33940;
  assign n33942 = ~P1_P3_DATAWIDTH_REG_21_ & n33941;
  assign n33943 = n33939 & n33942;
  assign n33944 = ~P1_P3_DATAWIDTH_REG_14_ & ~P1_P3_DATAWIDTH_REG_15_;
  assign n33945 = ~P1_P3_DATAWIDTH_REG_16_ & n33944;
  assign n33946 = ~P1_P3_DATAWIDTH_REG_17_ & n33945;
  assign n33947 = ~P1_P3_DATAWIDTH_REG_10_ & ~P1_P3_DATAWIDTH_REG_11_;
  assign n33948 = ~P1_P3_DATAWIDTH_REG_12_ & n33947;
  assign n33949 = ~P1_P3_DATAWIDTH_REG_13_ & n33948;
  assign n33950 = n33946 & n33949;
  assign n33951 = ~P1_P3_DATAWIDTH_REG_6_ & ~P1_P3_DATAWIDTH_REG_7_;
  assign n33952 = ~P1_P3_DATAWIDTH_REG_8_ & n33951;
  assign n33953 = ~P1_P3_DATAWIDTH_REG_9_ & n33952;
  assign n33954 = ~P1_P3_DATAWIDTH_REG_2_ & ~P1_P3_DATAWIDTH_REG_3_;
  assign n33955 = ~P1_P3_DATAWIDTH_REG_4_ & n33954;
  assign n33956 = ~P1_P3_DATAWIDTH_REG_5_ & n33955;
  assign n33957 = n33953 & n33956;
  assign n33958 = n33936 & n33943;
  assign n33959 = n33950 & n33958;
  assign n33960 = n33957 & n33959;
  assign n33961 = n33929 & n33960;
  assign n33962 = P1_P3_BYTEENABLE_REG_3_ & ~n33960;
  assign n33963 = ~P1_P3_DATAWIDTH_REG_0_ & ~P1_P3_REIP_REG_0_;
  assign n33964 = ~P1_P3_DATAWIDTH_REG_1_ & n33963;
  assign n33965 = n33960 & n33964;
  assign n33966 = ~n33961 & ~n33962;
  assign n5421 = n33965 | ~n33966;
  assign n33968 = P1_P3_REIP_REG_0_ & P1_P3_REIP_REG_1_;
  assign n33969 = P1_P3_DATAWIDTH_REG_0_ & ~P1_P3_REIP_REG_0_;
  assign n33970 = ~P1_P3_DATAWIDTH_REG_0_ & ~P1_P3_DATAWIDTH_REG_1_;
  assign n33971 = ~n33969 & ~n33970;
  assign n33972 = ~P1_P3_REIP_REG_1_ & ~n33971;
  assign n33973 = ~n33968 & ~n33972;
  assign n33974 = n33960 & ~n33973;
  assign n33975 = P1_P3_BYTEENABLE_REG_2_ & ~n33960;
  assign n5426 = n33974 | n33975;
  assign n33977 = P1_P3_REIP_REG_1_ & n33960;
  assign n33978 = P1_P3_BYTEENABLE_REG_1_ & ~n33960;
  assign n33979 = ~n33977 & ~n33978;
  assign n5431 = n33965 | ~n33979;
  assign n33981 = ~P1_P3_REIP_REG_0_ & ~P1_P3_REIP_REG_1_;
  assign n33982 = n33960 & ~n33981;
  assign n33983 = P1_P3_BYTEENABLE_REG_0_ & ~n33960;
  assign n5436 = n33982 | n33983;
  assign n33985 = P1_P3_W_R_N_REG & ~n25094;
  assign n33986 = ~P1_P3_READREQUEST_REG & n25094;
  assign n5441 = n33985 | n33986;
  assign n33988 = n25762 & n25994;
  assign n33989 = ~n25710 & n25994;
  assign n33990 = P1_P3_FLUSH_REG & ~n33989;
  assign n5446 = n33988 | n33990;
  assign n33992 = P1_P3_MORE_REG & ~n33989;
  assign n33993 = ~n25756 & n33989;
  assign n5451 = n33992 | n33993;
  assign n33995 = BS & ~n25315;
  assign n33996 = P1_P3_STATEBS16_REG & n25315;
  assign n33997 = ~P1_P3_STATE_REG_0_ & n25270;
  assign n33998 = ~n33995 & ~n33996;
  assign n5456 = n33997 | ~n33998;
  assign n34000 = ~n25640 & ~n25713;
  assign n34001 = ~n25358 & ~n34000;
  assign n34002 = ~P1_P3_STATEBS16_REG & n25640;
  assign n34003 = ~n25267 & ~n34002;
  assign n34004 = P1_P3_STATE2_REG_2_ & ~n34001;
  assign n34005 = n34003 & n34004;
  assign n34006 = P1_P3_STATE2_REG_0_ & ~n34005;
  assign n34007 = ~n26010 & ~n34006;
  assign n34008 = ~n25267 & n25352;
  assign n34009 = ~n26000 & ~n34008;
  assign n34010 = ~P1_P3_STATE2_REG_0_ & ~n34009;
  assign n34011 = ~n26072 & ~n34010;
  assign n34012 = ~n33047 & n34011;
  assign n34013 = ~n34007 & ~n34012;
  assign n34014 = P1_P3_REQUESTPENDING_REG & n34012;
  assign n5461 = n34013 | n34014;
  assign n34016 = P1_P3_D_C_N_REG & ~n25094;
  assign n34017 = ~P1_P3_CODEFETCH_REG & n25094;
  assign n34018 = ~n34016 & ~n34017;
  assign n5466 = n33997 | ~n34018;
  assign n34020 = P1_P3_MEMORYFETCH_REG & n25094;
  assign n34021 = P1_P3_M_IO_N_REG & ~n25094;
  assign n5471 = n34020 | n34021;
  assign n34023 = P1_P3_STATE2_REG_0_ & n27607;
  assign n34024 = n25709 & n25994;
  assign n34025 = P1_P3_CODEFETCH_REG & ~n34024;
  assign n5476 = n34023 | n34025;
  assign n34027 = P1_P3_STATE_REG_0_ & P1_P3_ADS_N_REG;
  assign n5481 = ~n25315 | n34027;
  assign n34029 = P1_P3_STATE2_REG_2_ & ~n25722;
  assign n34030 = ~n25717 & n34029;
  assign n34031 = ~n27607 & ~n33047;
  assign n34032 = ~n34030 & ~n34031;
  assign n34033 = P1_P3_READREQUEST_REG & n34031;
  assign n5486 = n34032 | n34033;
  assign n34035 = P1_P3_STATE2_REG_2_ & n25639;
  assign n34036 = ~n34031 & ~n34035;
  assign n34037 = P1_P3_MEMORYFETCH_REG & n34031;
  assign n5491 = n34036 | n34037;
  assign n34039 = P1_P2_STATE_REG_1_ & ~P1_P2_STATE_REG_0_;
  assign n34040 = P1_P2_BYTEENABLE_REG_3_ & n34039;
  assign n34041 = P1_P2_BE_N_REG_3_ & ~n34039;
  assign n5496 = n34040 | n34041;
  assign n34043 = P1_P2_BYTEENABLE_REG_2_ & n34039;
  assign n34044 = P1_P2_BE_N_REG_2_ & ~n34039;
  assign n5501 = n34043 | n34044;
  assign n34046 = P1_P2_BYTEENABLE_REG_1_ & n34039;
  assign n34047 = P1_P2_BE_N_REG_1_ & ~n34039;
  assign n5506 = n34046 | n34047;
  assign n34049 = P1_P2_BYTEENABLE_REG_0_ & n34039;
  assign n34050 = P1_P2_BE_N_REG_0_ & ~n34039;
  assign n5511 = n34049 | n34050;
  assign n34052 = P1_P2_STATE_REG_2_ & n34039;
  assign n34053 = P1_P2_REIP_REG_30_ & n34052;
  assign n34054 = ~P1_P2_STATE_REG_2_ & n34039;
  assign n34055 = P1_P2_REIP_REG_31_ & n34054;
  assign n34056 = P1_P2_ADDRESS_REG_29_ & ~n34039;
  assign n34057 = ~n34053 & ~n34055;
  assign n5516 = n34056 | ~n34057;
  assign n34059 = P1_P2_REIP_REG_29_ & n34052;
  assign n34060 = P1_P2_REIP_REG_30_ & n34054;
  assign n34061 = P1_P2_ADDRESS_REG_28_ & ~n34039;
  assign n34062 = ~n34059 & ~n34060;
  assign n5521 = n34061 | ~n34062;
  assign n34064 = P1_P2_REIP_REG_28_ & n34052;
  assign n34065 = P1_P2_REIP_REG_29_ & n34054;
  assign n34066 = P1_P2_ADDRESS_REG_27_ & ~n34039;
  assign n34067 = ~n34064 & ~n34065;
  assign n5526 = n34066 | ~n34067;
  assign n34069 = P1_P2_REIP_REG_27_ & n34052;
  assign n34070 = P1_P2_REIP_REG_28_ & n34054;
  assign n34071 = P1_P2_ADDRESS_REG_26_ & ~n34039;
  assign n34072 = ~n34069 & ~n34070;
  assign n5531 = n34071 | ~n34072;
  assign n34074 = P1_P2_REIP_REG_26_ & n34052;
  assign n34075 = P1_P2_REIP_REG_27_ & n34054;
  assign n34076 = P1_P2_ADDRESS_REG_25_ & ~n34039;
  assign n34077 = ~n34074 & ~n34075;
  assign n5536 = n34076 | ~n34077;
  assign n34079 = P1_P2_REIP_REG_25_ & n34052;
  assign n34080 = P1_P2_REIP_REG_26_ & n34054;
  assign n34081 = P1_P2_ADDRESS_REG_24_ & ~n34039;
  assign n34082 = ~n34079 & ~n34080;
  assign n5541 = n34081 | ~n34082;
  assign n34084 = P1_P2_REIP_REG_24_ & n34052;
  assign n34085 = P1_P2_REIP_REG_25_ & n34054;
  assign n34086 = P1_P2_ADDRESS_REG_23_ & ~n34039;
  assign n34087 = ~n34084 & ~n34085;
  assign n5546 = n34086 | ~n34087;
  assign n34089 = P1_P2_REIP_REG_23_ & n34052;
  assign n34090 = P1_P2_REIP_REG_24_ & n34054;
  assign n34091 = P1_P2_ADDRESS_REG_22_ & ~n34039;
  assign n34092 = ~n34089 & ~n34090;
  assign n5551 = n34091 | ~n34092;
  assign n34094 = P1_P2_REIP_REG_22_ & n34052;
  assign n34095 = P1_P2_REIP_REG_23_ & n34054;
  assign n34096 = P1_P2_ADDRESS_REG_21_ & ~n34039;
  assign n34097 = ~n34094 & ~n34095;
  assign n5556 = n34096 | ~n34097;
  assign n34099 = P1_P2_REIP_REG_21_ & n34052;
  assign n34100 = P1_P2_REIP_REG_22_ & n34054;
  assign n34101 = P1_P2_ADDRESS_REG_20_ & ~n34039;
  assign n34102 = ~n34099 & ~n34100;
  assign n5561 = n34101 | ~n34102;
  assign n34104 = P1_P2_REIP_REG_20_ & n34052;
  assign n34105 = P1_P2_REIP_REG_21_ & n34054;
  assign n34106 = P1_P2_ADDRESS_REG_19_ & ~n34039;
  assign n34107 = ~n34104 & ~n34105;
  assign n5566 = n34106 | ~n34107;
  assign n34109 = P1_P2_REIP_REG_19_ & n34052;
  assign n34110 = P1_P2_REIP_REG_20_ & n34054;
  assign n34111 = P1_P2_ADDRESS_REG_18_ & ~n34039;
  assign n34112 = ~n34109 & ~n34110;
  assign n5571 = n34111 | ~n34112;
  assign n34114 = P1_P2_REIP_REG_18_ & n34052;
  assign n34115 = P1_P2_REIP_REG_19_ & n34054;
  assign n34116 = P1_P2_ADDRESS_REG_17_ & ~n34039;
  assign n34117 = ~n34114 & ~n34115;
  assign n5576 = n34116 | ~n34117;
  assign n34119 = P1_P2_REIP_REG_17_ & n34052;
  assign n34120 = P1_P2_REIP_REG_18_ & n34054;
  assign n34121 = P1_P2_ADDRESS_REG_16_ & ~n34039;
  assign n34122 = ~n34119 & ~n34120;
  assign n5581 = n34121 | ~n34122;
  assign n34124 = P1_P2_REIP_REG_16_ & n34052;
  assign n34125 = P1_P2_REIP_REG_17_ & n34054;
  assign n34126 = P1_P2_ADDRESS_REG_15_ & ~n34039;
  assign n34127 = ~n34124 & ~n34125;
  assign n5586 = n34126 | ~n34127;
  assign n34129 = P1_P2_REIP_REG_15_ & n34052;
  assign n34130 = P1_P2_REIP_REG_16_ & n34054;
  assign n34131 = P1_P2_ADDRESS_REG_14_ & ~n34039;
  assign n34132 = ~n34129 & ~n34130;
  assign n5591 = n34131 | ~n34132;
  assign n34134 = P1_P2_REIP_REG_14_ & n34052;
  assign n34135 = P1_P2_REIP_REG_15_ & n34054;
  assign n34136 = P1_P2_ADDRESS_REG_13_ & ~n34039;
  assign n34137 = ~n34134 & ~n34135;
  assign n5596 = n34136 | ~n34137;
  assign n34139 = P1_P2_REIP_REG_13_ & n34052;
  assign n34140 = P1_P2_REIP_REG_14_ & n34054;
  assign n34141 = P1_P2_ADDRESS_REG_12_ & ~n34039;
  assign n34142 = ~n34139 & ~n34140;
  assign n5601 = n34141 | ~n34142;
  assign n34144 = P1_P2_REIP_REG_12_ & n34052;
  assign n34145 = P1_P2_REIP_REG_13_ & n34054;
  assign n34146 = P1_P2_ADDRESS_REG_11_ & ~n34039;
  assign n34147 = ~n34144 & ~n34145;
  assign n5606 = n34146 | ~n34147;
  assign n34149 = P1_P2_REIP_REG_11_ & n34052;
  assign n34150 = P1_P2_REIP_REG_12_ & n34054;
  assign n34151 = P1_P2_ADDRESS_REG_10_ & ~n34039;
  assign n34152 = ~n34149 & ~n34150;
  assign n5611 = n34151 | ~n34152;
  assign n34154 = P1_P2_REIP_REG_10_ & n34052;
  assign n34155 = P1_P2_REIP_REG_11_ & n34054;
  assign n34156 = P1_P2_ADDRESS_REG_9_ & ~n34039;
  assign n34157 = ~n34154 & ~n34155;
  assign n5616 = n34156 | ~n34157;
  assign n34159 = P1_P2_REIP_REG_9_ & n34052;
  assign n34160 = P1_P2_REIP_REG_10_ & n34054;
  assign n34161 = P1_P2_ADDRESS_REG_8_ & ~n34039;
  assign n34162 = ~n34159 & ~n34160;
  assign n5621 = n34161 | ~n34162;
  assign n34164 = P1_P2_REIP_REG_8_ & n34052;
  assign n34165 = P1_P2_REIP_REG_9_ & n34054;
  assign n34166 = P1_P2_ADDRESS_REG_7_ & ~n34039;
  assign n34167 = ~n34164 & ~n34165;
  assign n5626 = n34166 | ~n34167;
  assign n34169 = P1_P2_REIP_REG_7_ & n34052;
  assign n34170 = P1_P2_REIP_REG_8_ & n34054;
  assign n34171 = P1_P2_ADDRESS_REG_6_ & ~n34039;
  assign n34172 = ~n34169 & ~n34170;
  assign n5631 = n34171 | ~n34172;
  assign n34174 = P1_P2_REIP_REG_6_ & n34052;
  assign n34175 = P1_P2_REIP_REG_7_ & n34054;
  assign n34176 = P1_P2_ADDRESS_REG_5_ & ~n34039;
  assign n34177 = ~n34174 & ~n34175;
  assign n5636 = n34176 | ~n34177;
  assign n34179 = P1_P2_REIP_REG_5_ & n34052;
  assign n34180 = P1_P2_REIP_REG_6_ & n34054;
  assign n34181 = P1_P2_ADDRESS_REG_4_ & ~n34039;
  assign n34182 = ~n34179 & ~n34180;
  assign n5641 = n34181 | ~n34182;
  assign n34184 = P1_P2_REIP_REG_4_ & n34052;
  assign n34185 = P1_P2_REIP_REG_5_ & n34054;
  assign n34186 = P1_P2_ADDRESS_REG_3_ & ~n34039;
  assign n34187 = ~n34184 & ~n34185;
  assign n5646 = n34186 | ~n34187;
  assign n34189 = P1_P2_REIP_REG_3_ & n34052;
  assign n34190 = P1_P2_REIP_REG_4_ & n34054;
  assign n34191 = P1_P2_ADDRESS_REG_2_ & ~n34039;
  assign n34192 = ~n34189 & ~n34190;
  assign n5651 = n34191 | ~n34192;
  assign n34194 = P1_P2_REIP_REG_2_ & n34052;
  assign n34195 = P1_P2_REIP_REG_3_ & n34054;
  assign n34196 = P1_P2_ADDRESS_REG_1_ & ~n34039;
  assign n34197 = ~n34194 & ~n34195;
  assign n5656 = n34196 | ~n34197;
  assign n34199 = P1_P2_REIP_REG_1_ & n34052;
  assign n34200 = P1_P2_REIP_REG_2_ & n34054;
  assign n34201 = P1_P2_ADDRESS_REG_0_ & ~n34039;
  assign n34202 = ~n34199 & ~n34200;
  assign n5661 = n34201 | ~n34202;
  assign n34204 = ~P1_P2_STATE_REG_2_ & P1_P2_STATE_REG_1_;
  assign n34205 = NA & n34204;
  assign n34206 = P1_P2_STATE_REG_0_ & ~n34205;
  assign n34207 = ~HOLD & ~P1_P2_REQUESTPENDING_REG;
  assign n34208 = P1_READY12_REG & P1_READY21_REG;
  assign n34209 = ~n34207 & n34208;
  assign n34210 = n34204 & n34209;
  assign n34211 = ~P1_P2_STATE_REG_2_ & ~P1_P2_STATE_REG_1_;
  assign n34212 = HOLD & ~P1_P2_REQUESTPENDING_REG;
  assign n34213 = n34211 & n34212;
  assign n34214 = ~n34210 & ~n34213;
  assign n34215 = n34206 & ~n34214;
  assign n34216 = ~n34052 & ~n34215;
  assign n34217 = ~HOLD & P1_P2_REQUESTPENDING_REG;
  assign n34218 = P1_P2_STATE_REG_0_ & ~n34217;
  assign n34219 = ~n34207 & n34218;
  assign n34220 = ~NA & ~P1_P2_STATE_REG_0_;
  assign n34221 = n34207 & ~n34208;
  assign n34222 = ~n34208 & n34217;
  assign n34223 = P1_P2_STATE_REG_1_ & ~n34221;
  assign n34224 = ~n34222 & n34223;
  assign n34225 = ~n34219 & ~n34220;
  assign n34226 = ~n34224 & n34225;
  assign n34227 = P1_P2_STATE_REG_2_ & ~n34226;
  assign n5666 = ~n34216 | n34227;
  assign n34229 = P1_P2_STATE_REG_2_ & ~n34218;
  assign n34230 = P1_P2_STATE_REG_0_ & P1_P2_REQUESTPENDING_REG;
  assign n34231 = ~P1_P2_STATE_REG_2_ & n34230;
  assign n34232 = ~n34229 & ~n34231;
  assign n34233 = ~P1_P2_STATE_REG_1_ & ~n34232;
  assign n34234 = HOLD & ~n34208;
  assign n34235 = P1_P2_STATE_REG_0_ & ~n34234;
  assign n34236 = P1_P2_STATE_REG_2_ & ~n34235;
  assign n34237 = ~n34221 & ~n34236;
  assign n34238 = P1_P2_STATE_REG_1_ & n34237;
  assign n34239 = n34039 & n34208;
  assign n34240 = ~n34054 & ~n34239;
  assign n34241 = ~n34233 & ~n34238;
  assign n5671 = ~n34240 | ~n34241;
  assign n34243 = P1_P2_STATE_REG_1_ & ~n34222;
  assign n34244 = n34230 & ~n34243;
  assign n34245 = ~P1_P2_STATE_REG_2_ & ~n34244;
  assign n34246 = P1_P2_STATE_REG_2_ & n34218;
  assign n34247 = NA & ~P1_P2_STATE_REG_0_;
  assign n34248 = P1_P2_STATE_REG_2_ & ~n34217;
  assign n34249 = ~n34247 & ~n34248;
  assign n34250 = ~P1_P2_STATE_REG_1_ & ~n34249;
  assign n34251 = ~n34245 & ~n34246;
  assign n5676 = n34250 | ~n34251;
  assign n34253 = ~BS & ~n34211;
  assign n34254 = P1_P2_STATE_REG_0_ & n34204;
  assign n34255 = ~P1_P2_STATE_REG_1_ & ~P1_P2_STATE_REG_0_;
  assign n34256 = ~n34254 & ~n34255;
  assign n34257 = n34253 & ~n34256;
  assign n34258 = P1_P2_DATAWIDTH_REG_0_ & n34256;
  assign n5681 = n34257 | n34258;
  assign n34260 = P1_P2_DATAWIDTH_REG_1_ & n34256;
  assign n34261 = ~n34253 & ~n34256;
  assign n5686 = n34260 | n34261;
  assign n5691 = P1_P2_DATAWIDTH_REG_2_ & n34256;
  assign n5696 = P1_P2_DATAWIDTH_REG_3_ & n34256;
  assign n5701 = P1_P2_DATAWIDTH_REG_4_ & n34256;
  assign n5706 = P1_P2_DATAWIDTH_REG_5_ & n34256;
  assign n5711 = P1_P2_DATAWIDTH_REG_6_ & n34256;
  assign n5716 = P1_P2_DATAWIDTH_REG_7_ & n34256;
  assign n5721 = P1_P2_DATAWIDTH_REG_8_ & n34256;
  assign n5726 = P1_P2_DATAWIDTH_REG_9_ & n34256;
  assign n5731 = P1_P2_DATAWIDTH_REG_10_ & n34256;
  assign n5736 = P1_P2_DATAWIDTH_REG_11_ & n34256;
  assign n5741 = P1_P2_DATAWIDTH_REG_12_ & n34256;
  assign n5746 = P1_P2_DATAWIDTH_REG_13_ & n34256;
  assign n5751 = P1_P2_DATAWIDTH_REG_14_ & n34256;
  assign n5756 = P1_P2_DATAWIDTH_REG_15_ & n34256;
  assign n5761 = P1_P2_DATAWIDTH_REG_16_ & n34256;
  assign n5766 = P1_P2_DATAWIDTH_REG_17_ & n34256;
  assign n5771 = P1_P2_DATAWIDTH_REG_18_ & n34256;
  assign n5776 = P1_P2_DATAWIDTH_REG_19_ & n34256;
  assign n5781 = P1_P2_DATAWIDTH_REG_20_ & n34256;
  assign n5786 = P1_P2_DATAWIDTH_REG_21_ & n34256;
  assign n5791 = P1_P2_DATAWIDTH_REG_22_ & n34256;
  assign n5796 = P1_P2_DATAWIDTH_REG_23_ & n34256;
  assign n5801 = P1_P2_DATAWIDTH_REG_24_ & n34256;
  assign n5806 = P1_P2_DATAWIDTH_REG_25_ & n34256;
  assign n5811 = P1_P2_DATAWIDTH_REG_26_ & n34256;
  assign n5816 = P1_P2_DATAWIDTH_REG_27_ & n34256;
  assign n5821 = P1_P2_DATAWIDTH_REG_28_ & n34256;
  assign n5826 = P1_P2_DATAWIDTH_REG_29_ & n34256;
  assign n5831 = P1_P2_DATAWIDTH_REG_30_ & n34256;
  assign n5836 = P1_P2_DATAWIDTH_REG_31_ & n34256;
  assign n34293 = P1_P2_STATE2_REG_2_ & P1_P2_STATE2_REG_1_;
  assign n34294 = P1_P2_STATE2_REG_1_ & n34208;
  assign n34295 = ~P1_P2_STATE2_REG_0_ & ~n34294;
  assign n34296 = ~P1_P2_STATEBS16_REG & ~n34208;
  assign n34297 = P1_P2_STATE_REG_2_ & ~P1_P2_STATE_REG_1_;
  assign n34298 = ~n34204 & ~n34297;
  assign n34299 = ~P1_P2_STATE_REG_0_ & ~n34298;
  assign n34300 = n34296 & n34299;
  assign n34301 = P1_P2_INSTQUEUERD_ADDR_REG_1_ & P1_P2_INSTQUEUERD_ADDR_REG_0_;
  assign n34302 = ~P1_P2_INSTQUEUERD_ADDR_REG_2_ & n34301;
  assign n34303 = P1_P2_INSTQUEUERD_ADDR_REG_3_ & n34302;
  assign n34304 = P1_P2_INSTQUEUE_REG_11__5_ & n34303;
  assign n34305 = P1_P2_INSTQUEUERD_ADDR_REG_1_ & ~P1_P2_INSTQUEUERD_ADDR_REG_0_;
  assign n34306 = ~P1_P2_INSTQUEUERD_ADDR_REG_2_ & n34305;
  assign n34307 = P1_P2_INSTQUEUERD_ADDR_REG_3_ & n34306;
  assign n34308 = P1_P2_INSTQUEUE_REG_10__5_ & n34307;
  assign n34309 = ~n34304 & ~n34308;
  assign n34310 = ~P1_P2_INSTQUEUERD_ADDR_REG_1_ & P1_P2_INSTQUEUERD_ADDR_REG_0_;
  assign n34311 = ~P1_P2_INSTQUEUERD_ADDR_REG_2_ & n34310;
  assign n34312 = P1_P2_INSTQUEUERD_ADDR_REG_3_ & n34311;
  assign n34313 = P1_P2_INSTQUEUE_REG_9__5_ & n34312;
  assign n34314 = ~P1_P2_INSTQUEUERD_ADDR_REG_1_ & ~P1_P2_INSTQUEUERD_ADDR_REG_0_;
  assign n34315 = ~P1_P2_INSTQUEUERD_ADDR_REG_2_ & n34314;
  assign n34316 = P1_P2_INSTQUEUERD_ADDR_REG_3_ & n34315;
  assign n34317 = P1_P2_INSTQUEUE_REG_8__5_ & n34316;
  assign n34318 = ~n34313 & ~n34317;
  assign n34319 = P1_P2_INSTQUEUERD_ADDR_REG_3_ & P1_P2_INSTQUEUERD_ADDR_REG_2_;
  assign n34320 = n34301 & n34319;
  assign n34321 = P1_P2_INSTQUEUE_REG_15__5_ & n34320;
  assign n34322 = n34305 & n34319;
  assign n34323 = P1_P2_INSTQUEUE_REG_14__5_ & n34322;
  assign n34324 = n34310 & n34319;
  assign n34325 = P1_P2_INSTQUEUE_REG_13__5_ & n34324;
  assign n34326 = n34314 & n34319;
  assign n34327 = P1_P2_INSTQUEUE_REG_12__5_ & n34326;
  assign n34328 = ~n34321 & ~n34323;
  assign n34329 = ~n34325 & n34328;
  assign n34330 = ~n34327 & n34329;
  assign n34331 = ~P1_P2_INSTQUEUERD_ADDR_REG_3_ & P1_P2_INSTQUEUERD_ADDR_REG_2_;
  assign n34332 = n34301 & n34331;
  assign n34333 = P1_P2_INSTQUEUE_REG_7__5_ & n34332;
  assign n34334 = n34305 & n34331;
  assign n34335 = P1_P2_INSTQUEUE_REG_6__5_ & n34334;
  assign n34336 = n34310 & n34331;
  assign n34337 = P1_P2_INSTQUEUE_REG_5__5_ & n34336;
  assign n34338 = n34314 & n34331;
  assign n34339 = P1_P2_INSTQUEUE_REG_4__5_ & n34338;
  assign n34340 = ~n34333 & ~n34335;
  assign n34341 = ~n34337 & n34340;
  assign n34342 = ~n34339 & n34341;
  assign n34343 = ~P1_P2_INSTQUEUERD_ADDR_REG_3_ & n34302;
  assign n34344 = P1_P2_INSTQUEUE_REG_3__5_ & n34343;
  assign n34345 = ~P1_P2_INSTQUEUERD_ADDR_REG_3_ & ~P1_P2_INSTQUEUERD_ADDR_REG_2_;
  assign n34346 = n34305 & n34345;
  assign n34347 = P1_P2_INSTQUEUE_REG_2__5_ & n34346;
  assign n34348 = n34310 & n34345;
  assign n34349 = P1_P2_INSTQUEUE_REG_1__5_ & n34348;
  assign n34350 = ~P1_P2_INSTQUEUERD_ADDR_REG_3_ & n34315;
  assign n34351 = P1_P2_INSTQUEUE_REG_0__5_ & n34350;
  assign n34352 = ~n34344 & ~n34347;
  assign n34353 = ~n34349 & n34352;
  assign n34354 = ~n34351 & n34353;
  assign n34355 = n34309 & n34318;
  assign n34356 = n34330 & n34355;
  assign n34357 = n34342 & n34356;
  assign n34358 = n34354 & n34357;
  assign n34359 = P1_P2_INSTQUEUE_REG_11__6_ & n34303;
  assign n34360 = P1_P2_INSTQUEUE_REG_10__6_ & n34307;
  assign n34361 = ~n34359 & ~n34360;
  assign n34362 = P1_P2_INSTQUEUE_REG_9__6_ & n34312;
  assign n34363 = P1_P2_INSTQUEUE_REG_8__6_ & n34316;
  assign n34364 = ~n34362 & ~n34363;
  assign n34365 = P1_P2_INSTQUEUE_REG_15__6_ & n34320;
  assign n34366 = P1_P2_INSTQUEUE_REG_14__6_ & n34322;
  assign n34367 = P1_P2_INSTQUEUE_REG_13__6_ & n34324;
  assign n34368 = P1_P2_INSTQUEUE_REG_12__6_ & n34326;
  assign n34369 = ~n34365 & ~n34366;
  assign n34370 = ~n34367 & n34369;
  assign n34371 = ~n34368 & n34370;
  assign n34372 = P1_P2_INSTQUEUE_REG_7__6_ & n34332;
  assign n34373 = P1_P2_INSTQUEUE_REG_6__6_ & n34334;
  assign n34374 = P1_P2_INSTQUEUE_REG_5__6_ & n34336;
  assign n34375 = P1_P2_INSTQUEUE_REG_4__6_ & n34338;
  assign n34376 = ~n34372 & ~n34373;
  assign n34377 = ~n34374 & n34376;
  assign n34378 = ~n34375 & n34377;
  assign n34379 = P1_P2_INSTQUEUE_REG_3__6_ & n34343;
  assign n34380 = P1_P2_INSTQUEUE_REG_2__6_ & n34346;
  assign n34381 = P1_P2_INSTQUEUE_REG_1__6_ & n34348;
  assign n34382 = P1_P2_INSTQUEUE_REG_0__6_ & n34350;
  assign n34383 = ~n34379 & ~n34380;
  assign n34384 = ~n34381 & n34383;
  assign n34385 = ~n34382 & n34384;
  assign n34386 = n34361 & n34364;
  assign n34387 = n34371 & n34386;
  assign n34388 = n34378 & n34387;
  assign n34389 = n34385 & n34388;
  assign n34390 = n34358 & n34389;
  assign n34391 = P1_P2_INSTQUEUE_REG_11__4_ & n34303;
  assign n34392 = P1_P2_INSTQUEUE_REG_10__4_ & n34307;
  assign n34393 = ~n34391 & ~n34392;
  assign n34394 = P1_P2_INSTQUEUE_REG_9__4_ & n34312;
  assign n34395 = P1_P2_INSTQUEUE_REG_8__4_ & n34316;
  assign n34396 = ~n34394 & ~n34395;
  assign n34397 = P1_P2_INSTQUEUE_REG_15__4_ & n34320;
  assign n34398 = P1_P2_INSTQUEUE_REG_14__4_ & n34322;
  assign n34399 = P1_P2_INSTQUEUE_REG_13__4_ & n34324;
  assign n34400 = P1_P2_INSTQUEUE_REG_12__4_ & n34326;
  assign n34401 = ~n34397 & ~n34398;
  assign n34402 = ~n34399 & n34401;
  assign n34403 = ~n34400 & n34402;
  assign n34404 = P1_P2_INSTQUEUE_REG_7__4_ & n34332;
  assign n34405 = P1_P2_INSTQUEUE_REG_6__4_ & n34334;
  assign n34406 = P1_P2_INSTQUEUE_REG_5__4_ & n34336;
  assign n34407 = P1_P2_INSTQUEUE_REG_4__4_ & n34338;
  assign n34408 = ~n34404 & ~n34405;
  assign n34409 = ~n34406 & n34408;
  assign n34410 = ~n34407 & n34409;
  assign n34411 = P1_P2_INSTQUEUE_REG_3__4_ & n34343;
  assign n34412 = P1_P2_INSTQUEUE_REG_2__4_ & n34346;
  assign n34413 = P1_P2_INSTQUEUE_REG_1__4_ & n34348;
  assign n34414 = P1_P2_INSTQUEUE_REG_0__4_ & n34350;
  assign n34415 = ~n34411 & ~n34412;
  assign n34416 = ~n34413 & n34415;
  assign n34417 = ~n34414 & n34416;
  assign n34418 = n34393 & n34396;
  assign n34419 = n34403 & n34418;
  assign n34420 = n34410 & n34419;
  assign n34421 = n34417 & n34420;
  assign n34422 = P1_P2_INSTQUEUE_REG_11__7_ & n34303;
  assign n34423 = P1_P2_INSTQUEUE_REG_10__7_ & n34307;
  assign n34424 = ~n34422 & ~n34423;
  assign n34425 = P1_P2_INSTQUEUE_REG_9__7_ & n34312;
  assign n34426 = P1_P2_INSTQUEUE_REG_8__7_ & n34316;
  assign n34427 = ~n34425 & ~n34426;
  assign n34428 = P1_P2_INSTQUEUE_REG_15__7_ & n34320;
  assign n34429 = P1_P2_INSTQUEUE_REG_14__7_ & n34322;
  assign n34430 = P1_P2_INSTQUEUE_REG_13__7_ & n34324;
  assign n34431 = P1_P2_INSTQUEUE_REG_12__7_ & n34326;
  assign n34432 = ~n34428 & ~n34429;
  assign n34433 = ~n34430 & n34432;
  assign n34434 = ~n34431 & n34433;
  assign n34435 = P1_P2_INSTQUEUE_REG_7__7_ & n34332;
  assign n34436 = P1_P2_INSTQUEUE_REG_6__7_ & n34334;
  assign n34437 = P1_P2_INSTQUEUE_REG_5__7_ & n34336;
  assign n34438 = P1_P2_INSTQUEUE_REG_4__7_ & n34338;
  assign n34439 = ~n34435 & ~n34436;
  assign n34440 = ~n34437 & n34439;
  assign n34441 = ~n34438 & n34440;
  assign n34442 = P1_P2_INSTQUEUE_REG_3__7_ & n34343;
  assign n34443 = P1_P2_INSTQUEUE_REG_2__7_ & n34346;
  assign n34444 = P1_P2_INSTQUEUE_REG_1__7_ & n34348;
  assign n34445 = P1_P2_INSTQUEUE_REG_0__7_ & n34350;
  assign n34446 = ~n34442 & ~n34443;
  assign n34447 = ~n34444 & n34446;
  assign n34448 = ~n34445 & n34447;
  assign n34449 = n34424 & n34427;
  assign n34450 = n34434 & n34449;
  assign n34451 = n34441 & n34450;
  assign n34452 = n34448 & n34451;
  assign n34453 = P1_P2_INSTQUEUE_REG_11__3_ & n34303;
  assign n34454 = P1_P2_INSTQUEUE_REG_10__3_ & n34307;
  assign n34455 = ~n34453 & ~n34454;
  assign n34456 = P1_P2_INSTQUEUE_REG_9__3_ & n34312;
  assign n34457 = P1_P2_INSTQUEUE_REG_8__3_ & n34316;
  assign n34458 = ~n34456 & ~n34457;
  assign n34459 = P1_P2_INSTQUEUE_REG_15__3_ & n34320;
  assign n34460 = P1_P2_INSTQUEUE_REG_14__3_ & n34322;
  assign n34461 = P1_P2_INSTQUEUE_REG_13__3_ & n34324;
  assign n34462 = P1_P2_INSTQUEUE_REG_12__3_ & n34326;
  assign n34463 = ~n34459 & ~n34460;
  assign n34464 = ~n34461 & n34463;
  assign n34465 = ~n34462 & n34464;
  assign n34466 = P1_P2_INSTQUEUE_REG_7__3_ & n34332;
  assign n34467 = P1_P2_INSTQUEUE_REG_6__3_ & n34334;
  assign n34468 = P1_P2_INSTQUEUE_REG_5__3_ & n34336;
  assign n34469 = P1_P2_INSTQUEUE_REG_4__3_ & n34338;
  assign n34470 = ~n34466 & ~n34467;
  assign n34471 = ~n34468 & n34470;
  assign n34472 = ~n34469 & n34471;
  assign n34473 = P1_P2_INSTQUEUE_REG_3__3_ & n34343;
  assign n34474 = P1_P2_INSTQUEUE_REG_2__3_ & n34346;
  assign n34475 = P1_P2_INSTQUEUE_REG_1__3_ & n34348;
  assign n34476 = P1_P2_INSTQUEUE_REG_0__3_ & n34350;
  assign n34477 = ~n34473 & ~n34474;
  assign n34478 = ~n34475 & n34477;
  assign n34479 = ~n34476 & n34478;
  assign n34480 = n34455 & n34458;
  assign n34481 = n34465 & n34480;
  assign n34482 = n34472 & n34481;
  assign n34483 = n34479 & n34482;
  assign n34484 = P1_P2_INSTQUEUE_REG_11__2_ & n34303;
  assign n34485 = P1_P2_INSTQUEUE_REG_10__2_ & n34307;
  assign n34486 = ~n34484 & ~n34485;
  assign n34487 = P1_P2_INSTQUEUE_REG_9__2_ & n34312;
  assign n34488 = P1_P2_INSTQUEUE_REG_8__2_ & n34316;
  assign n34489 = ~n34487 & ~n34488;
  assign n34490 = P1_P2_INSTQUEUE_REG_15__2_ & n34320;
  assign n34491 = P1_P2_INSTQUEUE_REG_14__2_ & n34322;
  assign n34492 = P1_P2_INSTQUEUE_REG_13__2_ & n34324;
  assign n34493 = P1_P2_INSTQUEUE_REG_12__2_ & n34326;
  assign n34494 = ~n34490 & ~n34491;
  assign n34495 = ~n34492 & n34494;
  assign n34496 = ~n34493 & n34495;
  assign n34497 = P1_P2_INSTQUEUE_REG_7__2_ & n34332;
  assign n34498 = P1_P2_INSTQUEUE_REG_6__2_ & n34334;
  assign n34499 = P1_P2_INSTQUEUE_REG_5__2_ & n34336;
  assign n34500 = P1_P2_INSTQUEUE_REG_4__2_ & n34338;
  assign n34501 = ~n34497 & ~n34498;
  assign n34502 = ~n34499 & n34501;
  assign n34503 = ~n34500 & n34502;
  assign n34504 = P1_P2_INSTQUEUE_REG_3__2_ & n34343;
  assign n34505 = P1_P2_INSTQUEUE_REG_2__2_ & n34346;
  assign n34506 = P1_P2_INSTQUEUE_REG_1__2_ & n34348;
  assign n34507 = P1_P2_INSTQUEUE_REG_0__2_ & n34350;
  assign n34508 = ~n34504 & ~n34505;
  assign n34509 = ~n34506 & n34508;
  assign n34510 = ~n34507 & n34509;
  assign n34511 = n34486 & n34489;
  assign n34512 = n34496 & n34511;
  assign n34513 = n34503 & n34512;
  assign n34514 = n34510 & n34513;
  assign n34515 = ~n34452 & ~n34483;
  assign n34516 = n34514 & n34515;
  assign n34517 = n34390 & n34421;
  assign n34518 = n34516 & n34517;
  assign n34519 = P1_P2_INSTQUEUE_REG_11__1_ & n34303;
  assign n34520 = P1_P2_INSTQUEUE_REG_10__1_ & n34307;
  assign n34521 = ~n34519 & ~n34520;
  assign n34522 = P1_P2_INSTQUEUE_REG_9__1_ & n34312;
  assign n34523 = P1_P2_INSTQUEUE_REG_8__1_ & n34316;
  assign n34524 = ~n34522 & ~n34523;
  assign n34525 = P1_P2_INSTQUEUE_REG_15__1_ & n34320;
  assign n34526 = P1_P2_INSTQUEUE_REG_14__1_ & n34322;
  assign n34527 = P1_P2_INSTQUEUE_REG_13__1_ & n34324;
  assign n34528 = P1_P2_INSTQUEUE_REG_12__1_ & n34326;
  assign n34529 = ~n34525 & ~n34526;
  assign n34530 = ~n34527 & n34529;
  assign n34531 = ~n34528 & n34530;
  assign n34532 = P1_P2_INSTQUEUE_REG_7__1_ & n34332;
  assign n34533 = P1_P2_INSTQUEUE_REG_6__1_ & n34334;
  assign n34534 = P1_P2_INSTQUEUE_REG_5__1_ & n34336;
  assign n34535 = P1_P2_INSTQUEUE_REG_4__1_ & n34338;
  assign n34536 = ~n34532 & ~n34533;
  assign n34537 = ~n34534 & n34536;
  assign n34538 = ~n34535 & n34537;
  assign n34539 = P1_P2_INSTQUEUE_REG_3__1_ & n34343;
  assign n34540 = P1_P2_INSTQUEUE_REG_2__1_ & n34346;
  assign n34541 = P1_P2_INSTQUEUE_REG_1__1_ & n34348;
  assign n34542 = P1_P2_INSTQUEUE_REG_0__1_ & n34350;
  assign n34543 = ~n34539 & ~n34540;
  assign n34544 = ~n34541 & n34543;
  assign n34545 = ~n34542 & n34544;
  assign n34546 = n34521 & n34524;
  assign n34547 = n34531 & n34546;
  assign n34548 = n34538 & n34547;
  assign n34549 = n34545 & n34548;
  assign n34550 = P1_P2_INSTQUEUE_REG_11__0_ & n34303;
  assign n34551 = P1_P2_INSTQUEUE_REG_10__0_ & n34307;
  assign n34552 = ~n34550 & ~n34551;
  assign n34553 = P1_P2_INSTQUEUE_REG_9__0_ & n34312;
  assign n34554 = P1_P2_INSTQUEUE_REG_8__0_ & n34316;
  assign n34555 = ~n34553 & ~n34554;
  assign n34556 = P1_P2_INSTQUEUE_REG_15__0_ & n34320;
  assign n34557 = P1_P2_INSTQUEUE_REG_14__0_ & n34322;
  assign n34558 = P1_P2_INSTQUEUE_REG_13__0_ & n34324;
  assign n34559 = P1_P2_INSTQUEUE_REG_12__0_ & n34326;
  assign n34560 = ~n34556 & ~n34557;
  assign n34561 = ~n34558 & n34560;
  assign n34562 = ~n34559 & n34561;
  assign n34563 = P1_P2_INSTQUEUE_REG_7__0_ & n34332;
  assign n34564 = P1_P2_INSTQUEUE_REG_6__0_ & n34334;
  assign n34565 = P1_P2_INSTQUEUE_REG_5__0_ & n34336;
  assign n34566 = P1_P2_INSTQUEUE_REG_4__0_ & n34338;
  assign n34567 = ~n34563 & ~n34564;
  assign n34568 = ~n34565 & n34567;
  assign n34569 = ~n34566 & n34568;
  assign n34570 = P1_P2_INSTQUEUE_REG_3__0_ & n34343;
  assign n34571 = P1_P2_INSTQUEUE_REG_2__0_ & n34346;
  assign n34572 = P1_P2_INSTQUEUE_REG_1__0_ & n34348;
  assign n34573 = P1_P2_INSTQUEUE_REG_0__0_ & n34350;
  assign n34574 = ~n34570 & ~n34571;
  assign n34575 = ~n34572 & n34574;
  assign n34576 = ~n34573 & n34575;
  assign n34577 = n34552 & n34555;
  assign n34578 = n34562 & n34577;
  assign n34579 = n34569 & n34578;
  assign n34580 = n34576 & n34579;
  assign n34581 = n34549 & ~n34580;
  assign n34582 = n34518 & n34581;
  assign n34583 = n34300 & n34582;
  assign n34584 = ~P1_P2_STATE2_REG_1_ & ~n34583;
  assign n34585 = ~n34208 & n34299;
  assign n34586 = ~n34514 & ~n34549;
  assign n34587 = n34585 & n34586;
  assign n34588 = ~n34208 & ~n34514;
  assign n34589 = n34549 & n34588;
  assign n34590 = ~n34208 & n34514;
  assign n34591 = n34549 & ~n34585;
  assign n34592 = n34590 & ~n34591;
  assign n34593 = ~n34587 & ~n34589;
  assign n34594 = ~n34592 & n34593;
  assign n34595 = P1_P2_INSTQUEUERD_ADDR_REG_4_ & ~P1_P2_INSTQUEUEWR_ADDR_REG_4_;
  assign n34596 = ~P1_P2_INSTQUEUERD_ADDR_REG_3_ & P1_P2_INSTQUEUEWR_ADDR_REG_3_;
  assign n34597 = P1_P2_INSTQUEUERD_ADDR_REG_3_ & ~P1_P2_INSTQUEUEWR_ADDR_REG_3_;
  assign n34598 = ~P1_P2_INSTQUEUERD_ADDR_REG_2_ & P1_P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n34599 = P1_P2_INSTQUEUERD_ADDR_REG_2_ & ~P1_P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n34600 = P1_P2_INSTQUEUERD_ADDR_REG_0_ & ~P1_P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n34601 = P1_P2_INSTQUEUEWR_ADDR_REG_1_ & ~n34600;
  assign n34602 = ~P1_P2_INSTQUEUEWR_ADDR_REG_1_ & n34600;
  assign n34603 = ~P1_P2_INSTQUEUERD_ADDR_REG_1_ & ~n34602;
  assign n34604 = ~n34601 & ~n34603;
  assign n34605 = ~n34599 & ~n34604;
  assign n34606 = ~n34598 & ~n34605;
  assign n34607 = ~n34597 & ~n34606;
  assign n34608 = ~n34596 & ~n34607;
  assign n34609 = ~P1_P2_INSTQUEUERD_ADDR_REG_4_ & P1_P2_INSTQUEUEWR_ADDR_REG_4_;
  assign n34610 = n34608 & ~n34609;
  assign n34611 = ~n34595 & ~n34610;
  assign n34612 = ~n34595 & ~n34609;
  assign n34613 = ~n34608 & ~n34612;
  assign n34614 = n34608 & n34612;
  assign n34615 = ~n34613 & ~n34614;
  assign n34616 = ~n34596 & ~n34597;
  assign n34617 = ~n34606 & ~n34616;
  assign n34618 = n34606 & n34616;
  assign n34619 = ~n34617 & ~n34618;
  assign n34620 = ~P1_P2_INSTQUEUERD_ADDR_REG_1_ & P1_P2_INSTQUEUEWR_ADDR_REG_1_;
  assign n34621 = P1_P2_INSTQUEUERD_ADDR_REG_1_ & ~P1_P2_INSTQUEUEWR_ADDR_REG_1_;
  assign n34622 = ~n34620 & ~n34621;
  assign n34623 = ~n34600 & ~n34622;
  assign n34624 = n34600 & n34622;
  assign n34625 = ~n34623 & ~n34624;
  assign n34626 = ~n34598 & ~n34599;
  assign n34627 = ~n34604 & ~n34626;
  assign n34628 = n34604 & n34626;
  assign n34629 = ~n34627 & ~n34628;
  assign n34630 = n34615 & n34619;
  assign n34631 = n34625 & n34630;
  assign n34632 = n34629 & n34631;
  assign n34633 = n34611 & ~n34632;
  assign n34634 = ~n34549 & ~n34633;
  assign n34635 = n34549 & ~n34633;
  assign n34636 = ~n34634 & ~n34635;
  assign n34637 = ~n34452 & n34483;
  assign n34638 = ~n34358 & ~n34389;
  assign n34639 = n34421 & n34638;
  assign n34640 = n34637 & n34639;
  assign n34641 = n34580 & n34640;
  assign n34642 = n34636 & n34641;
  assign n34643 = ~n34514 & ~n34642;
  assign n34644 = ~n34483 & ~n34580;
  assign n34645 = ~n34452 & n34644;
  assign n34646 = n34517 & n34645;
  assign n34647 = ~n34634 & n34646;
  assign n34648 = ~n34635 & n34647;
  assign n34649 = n34514 & ~n34648;
  assign n34650 = ~n34643 & ~n34649;
  assign n34651 = n34594 & n34650;
  assign n34652 = ~P1_P2_FLUSH_REG & ~P1_P2_MORE_REG;
  assign n34653 = n34651 & ~n34652;
  assign n34654 = ~n34549 & n34580;
  assign n34655 = ~n34514 & n34654;
  assign n34656 = n34640 & n34655;
  assign n34657 = ~n34633 & n34656;
  assign n34658 = n34549 & n34580;
  assign n34659 = ~n34514 & n34658;
  assign n34660 = n34640 & n34659;
  assign n34661 = ~n34633 & n34660;
  assign n34662 = n34582 & ~n34633;
  assign n34663 = ~n34549 & ~n34580;
  assign n34664 = n34518 & n34663;
  assign n34665 = ~n34633 & n34664;
  assign n34666 = ~n34657 & ~n34661;
  assign n34667 = ~n34662 & n34666;
  assign n34668 = ~n34665 & n34667;
  assign n34669 = ~n34358 & n34389;
  assign n34670 = ~n34421 & n34669;
  assign n34671 = n34516 & n34670;
  assign n34672 = n34663 & n34671;
  assign n34673 = ~P1_P2_INSTQUEUERD_ADDR_REG_0_ & P1_P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n34674 = ~n34600 & ~n34673;
  assign n34675 = n34625 & n34674;
  assign n34676 = ~n34629 & ~n34675;
  assign n34677 = n34630 & ~n34676;
  assign n34678 = n34611 & ~n34677;
  assign n34679 = n34672 & ~n34678;
  assign n34680 = n34658 & n34671;
  assign n34681 = ~n34678 & n34680;
  assign n34682 = n34516 & n34639;
  assign n34683 = n34581 & n34682;
  assign n34684 = n34615 & ~n34676;
  assign n34685 = n34619 & n34684;
  assign n34686 = n34611 & ~n34685;
  assign n34687 = n34683 & ~n34686;
  assign n34688 = n34663 & n34682;
  assign n34689 = ~n34625 & ~n34674;
  assign n34690 = n34630 & ~n34689;
  assign n34691 = n34629 & n34690;
  assign n34692 = n34611 & ~n34691;
  assign n34693 = n34688 & ~n34692;
  assign n34694 = ~n34679 & ~n34681;
  assign n34695 = ~n34687 & n34694;
  assign n34696 = ~n34693 & n34695;
  assign n34697 = n34668 & n34696;
  assign n34698 = ~n34651 & ~n34697;
  assign n34699 = ~n34549 & ~n34692;
  assign n34700 = n34549 & ~n34686;
  assign n34701 = ~n34699 & ~n34700;
  assign n34702 = ~n34580 & n34682;
  assign n34703 = n34701 & n34702;
  assign n34704 = n34483 & n34514;
  assign n34705 = n34358 & ~n34389;
  assign n34706 = n34704 & n34705;
  assign n34707 = n34658 & n34706;
  assign n34708 = ~n34452 & n34707;
  assign n34709 = n34518 & ~n34580;
  assign n34710 = ~n34656 & ~n34708;
  assign n34711 = ~n34709 & n34710;
  assign n34712 = n34389 & n34483;
  assign n34713 = ~n34421 & n34514;
  assign n34714 = ~n34452 & n34658;
  assign n34715 = n34713 & n34714;
  assign n34716 = n34358 & ~n34514;
  assign n34717 = n34421 & n34452;
  assign n34718 = n34716 & n34717;
  assign n34719 = ~n34715 & ~n34718;
  assign n34720 = n34712 & ~n34719;
  assign n34721 = n34663 & n34717;
  assign n34722 = n34706 & n34721;
  assign n34723 = n34483 & ~n34514;
  assign n34724 = n34452 & n34654;
  assign n34725 = n34639 & n34723;
  assign n34726 = n34724 & n34725;
  assign n34727 = ~n34549 & n34682;
  assign n34728 = ~n34726 & ~n34727;
  assign n34729 = ~n34720 & ~n34722;
  assign n34730 = n34728 & n34729;
  assign n34731 = n34389 & ~n34452;
  assign n34732 = ~n34705 & ~n34731;
  assign n34733 = n34483 & n34732;
  assign n34734 = ~n34514 & ~n34733;
  assign n34735 = ~n34452 & ~n34705;
  assign n34736 = ~n34669 & n34735;
  assign n34737 = ~n34483 & n34736;
  assign n34738 = n34581 & ~n34737;
  assign n34739 = n34638 & n34658;
  assign n34740 = n34358 & n34452;
  assign n34741 = ~n34515 & ~n34740;
  assign n34742 = ~n34549 & n34741;
  assign n34743 = n34389 & n34421;
  assign n34744 = n34580 & n34743;
  assign n34745 = ~n34739 & ~n34742;
  assign n34746 = ~n34744 & n34745;
  assign n34747 = ~n34738 & n34746;
  assign n34748 = n34514 & ~n34747;
  assign n34749 = ~n34483 & ~n34743;
  assign n34750 = n34358 & n34749;
  assign n34751 = n34452 & n34549;
  assign n34752 = n34580 & ~n34751;
  assign n34753 = n34483 & ~n34752;
  assign n34754 = ~n34358 & n34753;
  assign n34755 = ~n34452 & ~n34638;
  assign n34756 = ~n34581 & n34755;
  assign n34757 = ~n34421 & ~n34756;
  assign n34758 = n34389 & ~n34549;
  assign n34759 = n34452 & n34758;
  assign n34760 = n34421 & ~n34549;
  assign n34761 = n34669 & n34760;
  assign n34762 = ~n34638 & n34654;
  assign n34763 = ~n34759 & ~n34761;
  assign n34764 = ~n34762 & n34763;
  assign n34765 = ~n34750 & ~n34754;
  assign n34766 = ~n34757 & n34765;
  assign n34767 = n34764 & n34766;
  assign n34768 = ~n34734 & ~n34748;
  assign n34769 = n34767 & n34768;
  assign n34770 = n34730 & n34769;
  assign n34771 = ~n34707 & n34770;
  assign n34772 = P1_P2_INSTQUEUERD_ADDR_REG_0_ & ~n34771;
  assign n34773 = n34711 & ~n34772;
  assign n34774 = ~P1_P2_INSTQUEUERD_ADDR_REG_2_ & ~n34773;
  assign n34775 = P1_P2_INSTQUEUERD_ADDR_REG_1_ & n34774;
  assign n34776 = P1_P2_INSTQUEUERD_ADDR_REG_2_ & ~n34711;
  assign n34777 = ~P1_P2_INSTQUEUERD_ADDR_REG_1_ & n34776;
  assign n34778 = ~P1_P2_INSTQUEUERD_ADDR_REG_2_ & P1_P2_INSTQUEUERD_ADDR_REG_1_;
  assign n34779 = P1_P2_INSTQUEUERD_ADDR_REG_2_ & ~P1_P2_INSTQUEUERD_ADDR_REG_1_;
  assign n34780 = ~n34778 & ~n34779;
  assign n34781 = n34660 & ~n34780;
  assign n34782 = P1_P2_INSTQUEUERD_ADDR_REG_2_ & ~n34301;
  assign n34783 = ~n34302 & ~n34782;
  assign n34784 = ~n34658 & ~n34663;
  assign n34785 = n34783 & ~n34784;
  assign n34786 = n34671 & n34785;
  assign n34787 = ~n34781 & ~n34786;
  assign n34788 = n34549 & n34712;
  assign n34789 = ~n34713 & ~n34718;
  assign n34790 = n34788 & ~n34789;
  assign n34791 = n34717 & ~n34784;
  assign n34792 = n34706 & n34791;
  assign n34793 = ~n34790 & ~n34792;
  assign n34794 = n34728 & n34793;
  assign n34795 = n34769 & n34794;
  assign n34796 = n34782 & ~n34795;
  assign n34797 = n34787 & ~n34796;
  assign n34798 = ~n34775 & ~n34777;
  assign n34799 = n34797 & n34798;
  assign n34800 = n34421 & n34580;
  assign n34801 = ~n34483 & ~n34654;
  assign n34802 = n34735 & ~n34800;
  assign n34803 = n34801 & n34802;
  assign n34804 = ~n34761 & n34803;
  assign n34805 = n34514 & ~n34804;
  assign n34806 = ~n34514 & ~n34641;
  assign n34807 = n34581 & ~n34736;
  assign n34808 = ~n34805 & ~n34806;
  assign n34809 = ~n34807 & n34808;
  assign n34810 = n34678 & n34680;
  assign n34811 = n34633 & n34660;
  assign n34812 = n34633 & n34664;
  assign n34813 = ~n34811 & ~n34812;
  assign n34814 = ~n34208 & ~n34813;
  assign n34815 = ~n34810 & ~n34814;
  assign n34816 = n34672 & n34678;
  assign n34817 = ~n34669 & n34713;
  assign n34818 = ~n34816 & ~n34817;
  assign n34819 = n34633 & n34656;
  assign n34820 = n34582 & n34633;
  assign n34821 = ~n34819 & ~n34820;
  assign n34822 = n34585 & ~n34821;
  assign n34823 = n34818 & ~n34822;
  assign n34824 = n34809 & n34815;
  assign n34825 = n34823 & n34824;
  assign n34826 = ~n34799 & ~n34825;
  assign n34827 = P1_P2_INSTQUEUERD_ADDR_REG_2_ & n34825;
  assign n34828 = ~n34826 & ~n34827;
  assign n34829 = P1_P2_INSTQUEUERD_ADDR_REG_1_ & n34331;
  assign n34830 = ~n34773 & n34829;
  assign n34831 = P1_P2_INSTQUEUERD_ADDR_REG_2_ & n34301;
  assign n34832 = P1_P2_INSTQUEUERD_ADDR_REG_3_ & ~n34831;
  assign n34833 = ~n34794 & n34832;
  assign n34834 = P1_P2_INSTQUEUERD_ADDR_REG_2_ & P1_P2_INSTQUEUERD_ADDR_REG_1_;
  assign n34835 = ~P1_P2_INSTQUEUERD_ADDR_REG_3_ & n34834;
  assign n34836 = P1_P2_INSTQUEUERD_ADDR_REG_3_ & ~n34834;
  assign n34837 = ~n34835 & ~n34836;
  assign n34838 = n34660 & ~n34837;
  assign n34839 = ~n34833 & ~n34838;
  assign n34840 = ~n34421 & n34708;
  assign n34841 = n34421 & n34708;
  assign n34842 = ~n34582 & ~n34664;
  assign n34843 = ~n34656 & n34842;
  assign n34844 = ~n34840 & ~n34841;
  assign n34845 = n34843 & n34844;
  assign n34846 = n34769 & n34845;
  assign n34847 = n34836 & ~n34846;
  assign n34848 = P1_P2_INSTQUEUERD_ADDR_REG_3_ & ~P1_P2_INSTQUEUERD_ADDR_REG_0_;
  assign n34849 = ~n34769 & n34848;
  assign n34850 = ~n34301 & n34345;
  assign n34851 = ~P1_P2_INSTQUEUERD_ADDR_REG_2_ & ~n34301;
  assign n34852 = P1_P2_INSTQUEUERD_ADDR_REG_3_ & ~n34851;
  assign n34853 = ~n34850 & ~n34852;
  assign n34854 = ~n34784 & n34853;
  assign n34855 = n34671 & n34854;
  assign n34856 = ~n34849 & ~n34855;
  assign n34857 = n34839 & ~n34847;
  assign n34858 = n34856 & n34857;
  assign n34859 = ~n34830 & n34858;
  assign n34860 = ~n34825 & ~n34859;
  assign n34861 = P1_P2_INSTQUEUERD_ADDR_REG_3_ & n34825;
  assign n34862 = ~n34860 & ~n34861;
  assign n34863 = ~n34828 & ~n34862;
  assign n34864 = P1_P2_INSTQUEUERD_ADDR_REG_4_ & n34825;
  assign n34865 = P1_P2_INSTQUEUERD_ADDR_REG_3_ & n34834;
  assign n34866 = ~P1_P2_INSTQUEUERD_ADDR_REG_4_ & n34865;
  assign n34867 = P1_P2_INSTQUEUERD_ADDR_REG_4_ & ~n34865;
  assign n34868 = ~n34866 & ~n34867;
  assign n34869 = n34660 & ~n34868;
  assign n34870 = ~n34825 & n34869;
  assign n34871 = ~n34864 & ~n34870;
  assign n34872 = ~n34863 & n34871;
  assign n34873 = ~P1_P2_INSTQUEUEWR_ADDR_REG_3_ & ~n34862;
  assign n34874 = ~P1_P2_INSTQUEUEWR_ADDR_REG_4_ & ~n34871;
  assign n34875 = P1_P2_INSTQUEUEWR_ADDR_REG_2_ & n34828;
  assign n34876 = P1_P2_INSTQUEUEWR_ADDR_REG_3_ & n34862;
  assign n34877 = n34669 & n34715;
  assign n34878 = ~n34672 & ~n34877;
  assign n34879 = n34707 & n34717;
  assign n34880 = n34770 & ~n34879;
  assign n34881 = n34878 & n34880;
  assign n34882 = ~P1_P2_INSTQUEUERD_ADDR_REG_0_ & ~n34881;
  assign n34883 = P1_P2_INSTQUEUERD_ADDR_REG_0_ & ~n34711;
  assign n34884 = P1_P2_INSTQUEUERD_ADDR_REG_0_ & n34660;
  assign n34885 = ~n34882 & ~n34883;
  assign n34886 = ~n34884 & n34885;
  assign n34887 = ~n34825 & ~n34886;
  assign n34888 = P1_P2_INSTQUEUERD_ADDR_REG_0_ & n34825;
  assign n34889 = ~n34887 & ~n34888;
  assign n34890 = P1_P2_INSTQUEUEWR_ADDR_REG_0_ & n34889;
  assign n34891 = ~P1_P2_INSTQUEUEWR_ADDR_REG_1_ & ~n34890;
  assign n34892 = ~P1_P2_INSTQUEUEWR_ADDR_REG_2_ & ~n34828;
  assign n34893 = ~P1_P2_INSTQUEUERD_ADDR_REG_1_ & ~n34773;
  assign n34894 = ~P1_P2_INSTQUEUERD_ADDR_REG_1_ & n34660;
  assign n34895 = ~n34301 & ~n34314;
  assign n34896 = ~n34878 & n34895;
  assign n34897 = ~n34894 & ~n34896;
  assign n34898 = n34305 & ~n34880;
  assign n34899 = n34897 & ~n34898;
  assign n34900 = ~n34893 & n34899;
  assign n34901 = ~n34825 & ~n34900;
  assign n34902 = P1_P2_INSTQUEUERD_ADDR_REG_1_ & n34825;
  assign n34903 = ~n34901 & ~n34902;
  assign n34904 = P1_P2_INSTQUEUEWR_ADDR_REG_1_ & n34890;
  assign n34905 = ~n34903 & ~n34904;
  assign n34906 = ~n34891 & ~n34892;
  assign n34907 = ~n34905 & n34906;
  assign n34908 = ~n34875 & ~n34876;
  assign n34909 = ~n34907 & n34908;
  assign n34910 = ~n34873 & ~n34874;
  assign n34911 = ~n34909 & n34910;
  assign n34912 = P1_P2_INSTQUEUEWR_ADDR_REG_4_ & n34871;
  assign n34913 = ~n34911 & ~n34912;
  assign n34914 = ~n34653 & ~n34698;
  assign n34915 = ~n34703 & n34914;
  assign n34916 = n34872 & n34915;
  assign n34917 = ~n34913 & n34916;
  assign n34918 = n34584 & n34917;
  assign n34919 = P1_P2_STATE2_REG_0_ & ~n34918;
  assign n34920 = ~n34295 & ~n34919;
  assign n34921 = P1_P2_STATE2_REG_2_ & n34920;
  assign n34922 = P1_P2_STATE2_REG_0_ & ~n34921;
  assign n34923 = n34293 & n34922;
  assign n34924 = P1_P2_STATE2_REG_3_ & ~n34922;
  assign n5841 = n34923 | n34924;
  assign n34926 = ~P1_P2_STATE2_REG_2_ & ~n34208;
  assign n34927 = P1_P2_STATE2_REG_0_ & ~n34926;
  assign n34928 = ~P1_P2_STATE2_REG_0_ & ~P1_P2_STATEBS16_REG;
  assign n34929 = ~n34927 & ~n34928;
  assign n34930 = P1_P2_STATE2_REG_1_ & n34929;
  assign n34931 = P1_P2_STATE2_REG_2_ & ~P1_P2_STATE2_REG_1_;
  assign n34932 = ~n34930 & ~n34931;
  assign n34933 = P1_P2_STATE2_REG_2_ & ~n34922;
  assign n5846 = ~n34932 | n34933;
  assign n34935 = P1_P2_STATE2_REG_0_ & n34931;
  assign n34936 = ~n34921 & n34935;
  assign n34937 = ~P1_P2_STATE2_REG_2_ & P1_P2_STATE2_REG_0_;
  assign n34938 = n34208 & n34937;
  assign n34939 = ~n34921 & ~n34938;
  assign n34940 = P1_P2_STATE2_REG_1_ & ~n34939;
  assign n34941 = ~P1_P2_STATE2_REG_3_ & ~P1_P2_STATE2_REG_1_;
  assign n34942 = ~n34208 & n34941;
  assign n34943 = n34922 & n34942;
  assign n34944 = P1_P2_STATE2_REG_1_ & ~P1_P2_STATE2_REG_0_;
  assign n34945 = ~P1_P2_STATE2_REG_2_ & n34944;
  assign n34946 = ~P1_P2_STATEBS16_REG & n34945;
  assign n34947 = ~n34936 & ~n34940;
  assign n34948 = ~n34943 & n34947;
  assign n5851 = n34946 | ~n34948;
  assign n34950 = P1_P2_STATE2_REG_3_ & ~P1_P2_INSTQUEUERD_ADDR_REG_4_;
  assign n34951 = ~P1_P2_STATE2_REG_2_ & ~P1_P2_STATE2_REG_1_;
  assign n34952 = n34950 & n34951;
  assign n34953 = ~n34921 & ~n34952;
  assign n34954 = ~P1_P2_STATE2_REG_0_ & n34953;
  assign n34955 = P1_P2_INSTADDRPOINTER_REG_0_ & P1_P2_INSTADDRPOINTER_REG_31_;
  assign n34956 = P1_P2_INSTADDRPOINTER_REG_0_ & ~P1_P2_INSTADDRPOINTER_REG_31_;
  assign n34957 = ~n34955 & ~n34956;
  assign n34958 = P1_P2_FLUSH_REG & n34957;
  assign n34959 = P1_P2_INSTQUEUERD_ADDR_REG_0_ & ~P1_P2_FLUSH_REG;
  assign n34960 = ~n34958 & ~n34959;
  assign n34961 = P1_P2_INSTADDRPOINTER_REG_0_ & ~P1_P2_INSTADDRPOINTER_REG_1_;
  assign n34962 = ~P1_P2_INSTADDRPOINTER_REG_0_ & P1_P2_INSTADDRPOINTER_REG_1_;
  assign n34963 = ~n34961 & ~n34962;
  assign n34964 = P1_P2_INSTADDRPOINTER_REG_31_ & ~n34963;
  assign n34965 = P1_P2_INSTADDRPOINTER_REG_1_ & ~P1_P2_INSTADDRPOINTER_REG_31_;
  assign n34966 = ~n34964 & ~n34965;
  assign n34967 = ~n34957 & n34966;
  assign n34968 = P1_P2_FLUSH_REG & n34967;
  assign n34969 = P1_P2_INSTQUEUERD_ADDR_REG_1_ & ~P1_P2_FLUSH_REG;
  assign n34970 = ~n34968 & ~n34969;
  assign n34971 = n34960 & n34970;
  assign n34972 = P1_P2_INSTQUEUERD_ADDR_REG_3_ & ~P1_P2_FLUSH_REG;
  assign n34973 = ~n34957 & ~n34966;
  assign n34974 = P1_P2_FLUSH_REG & n34973;
  assign n34975 = P1_P2_INSTQUEUERD_ADDR_REG_2_ & ~P1_P2_FLUSH_REG;
  assign n34976 = ~n34974 & ~n34975;
  assign n34977 = ~n34971 & n34972;
  assign n34978 = ~n34976 & n34977;
  assign n34979 = P1_P2_INSTQUEUERD_ADDR_REG_4_ & ~P1_P2_FLUSH_REG;
  assign n34980 = ~n34978 & ~n34979;
  assign n34981 = n34293 & n34980;
  assign n34982 = ~n34921 & ~n34981;
  assign n34983 = P1_P2_STATE2_REG_0_ & ~n34982;
  assign n34984 = P1_P2_STATE2_REG_3_ & P1_P2_STATE2_REG_0_;
  assign n34985 = n34951 & n34984;
  assign n34986 = ~n34938 & ~n34985;
  assign n34987 = ~n34917 & n34935;
  assign n34988 = n34986 & ~n34987;
  assign n34989 = ~n34954 & ~n34983;
  assign n5856 = ~n34988 | ~n34989;
  assign n34991 = P1_P2_INSTQUEUEWR_ADDR_REG_1_ & P1_P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n34992 = P1_P2_INSTQUEUEWR_ADDR_REG_2_ & n34991;
  assign n34993 = P1_P2_INSTQUEUEWR_ADDR_REG_3_ & n34992;
  assign n34994 = P1_P2_STATE2_REG_3_ & ~n34993;
  assign n34995 = ~P1_P2_STATE2_REG_2_ & P1_P2_STATE2_REG_1_;
  assign n34996 = ~n34931 & ~n34995;
  assign n34997 = ~n34950 & n34996;
  assign n34998 = ~P1_P2_STATE2_REG_0_ & ~n34997;
  assign n34999 = ~n34994 & n34998;
  assign n35000 = ~P1_P2_INSTQUEUEWR_ADDR_REG_2_ & n34991;
  assign n35001 = P1_P2_INSTQUEUEWR_ADDR_REG_2_ & ~n34991;
  assign n35002 = ~n35000 & ~n35001;
  assign n35003 = ~P1_P2_INSTQUEUEWR_ADDR_REG_3_ & n34992;
  assign n35004 = P1_P2_INSTQUEUEWR_ADDR_REG_3_ & ~n34992;
  assign n35005 = ~n35003 & ~n35004;
  assign n35006 = ~n35002 & ~n35005;
  assign n35007 = ~P1_P2_INSTQUEUEWR_ADDR_REG_1_ & P1_P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n35008 = P1_P2_INSTQUEUEWR_ADDR_REG_1_ & ~P1_P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n35009 = ~n35007 & ~n35008;
  assign n35010 = ~P1_P2_INSTQUEUEWR_ADDR_REG_0_ & ~n35009;
  assign n35011 = n35006 & n35010;
  assign n35012 = ~n34993 & ~n35011;
  assign n35013 = ~P1_P2_STATE2_REG_3_ & ~P1_P2_STATE2_REG_2_;
  assign n35014 = ~P1_P2_STATEBS16_REG & n35013;
  assign n35015 = ~P1_P2_STATE2_REG_2_ & ~n35014;
  assign n35016 = P1_P2_INSTQUEUEWR_ADDR_REG_0_ & ~n35009;
  assign n35017 = ~P1_P2_INSTQUEUEWR_ADDR_REG_0_ & n35009;
  assign n35018 = ~n35016 & ~n35017;
  assign n35019 = ~P1_P2_INSTQUEUEWR_ADDR_REG_0_ & ~n35018;
  assign n35020 = P1_P2_INSTQUEUEWR_ADDR_REG_0_ & n35018;
  assign n35021 = ~n35019 & ~n35020;
  assign n35022 = ~P1_P2_INSTQUEUEWR_ADDR_REG_0_ & ~n35021;
  assign n35023 = ~n35002 & ~n35010;
  assign n35024 = n35002 & n35010;
  assign n35025 = ~n35023 & ~n35024;
  assign n35026 = P1_P2_INSTQUEUEWR_ADDR_REG_0_ & ~n35018;
  assign n35027 = ~n35025 & ~n35026;
  assign n35028 = n35025 & n35026;
  assign n35029 = ~n35027 & ~n35028;
  assign n35030 = ~n35002 & n35005;
  assign n35031 = n35010 & n35030;
  assign n35032 = ~n35002 & n35010;
  assign n35033 = ~n35005 & ~n35032;
  assign n35034 = ~n35031 & ~n35033;
  assign n35035 = n35025 & ~n35034;
  assign n35036 = ~n35026 & ~n35034;
  assign n35037 = ~n35035 & ~n35036;
  assign n35038 = ~n35025 & n35034;
  assign n35039 = n35026 & n35038;
  assign n35040 = n35037 & ~n35039;
  assign n35041 = ~n35029 & ~n35040;
  assign n35042 = n35022 & n35041;
  assign n35043 = ~n35025 & ~n35034;
  assign n35044 = n35026 & n35043;
  assign n35045 = ~n35042 & ~n35044;
  assign n35046 = n35015 & ~n35045;
  assign n35047 = n35012 & ~n35046;
  assign n35048 = n34999 & ~n35047;
  assign n35049 = P1_P2_INSTQUEUE_REG_15__7_ & ~n35048;
  assign n35050 = P1_BUF1_REG_23_ & n12494;
  assign n35051 = P1_BUF2_REG_23_ & ~n12494;
  assign n35052 = ~n35050 & ~n35051;
  assign n35053 = P1_P2_STATEBS16_REG & n35013;
  assign n35054 = n34998 & n35053;
  assign n35055 = ~n35052 & n35054;
  assign n35056 = n35044 & n35055;
  assign n35057 = P1_P2_STATE2_REG_3_ & n34998;
  assign n35058 = ~n34452 & n35057;
  assign n35059 = n34993 & n35058;
  assign n35060 = ~n35056 & ~n35059;
  assign n35061 = P1_BUF1_REG_31_ & n12494;
  assign n35062 = P1_BUF2_REG_31_ & ~n12494;
  assign n35063 = ~n35061 & ~n35062;
  assign n35064 = n35054 & ~n35063;
  assign n35065 = n35042 & n35064;
  assign n35066 = n35060 & ~n35065;
  assign n35067 = n35045 & n35053;
  assign n35068 = n35015 & ~n35067;
  assign n35069 = ~n35012 & ~n35068;
  assign n35070 = P1_BUF1_REG_7_ & n12494;
  assign n35071 = P1_BUF2_REG_7_ & ~n12494;
  assign n35072 = ~n35070 & ~n35071;
  assign n35073 = n34998 & ~n35072;
  assign n35074 = n35069 & n35073;
  assign n35075 = ~n35049 & n35066;
  assign n5861 = n35074 | ~n35075;
  assign n35077 = P1_P2_INSTQUEUE_REG_15__6_ & ~n35048;
  assign n35078 = P1_BUF1_REG_22_ & n12494;
  assign n35079 = P1_BUF2_REG_22_ & ~n12494;
  assign n35080 = ~n35078 & ~n35079;
  assign n35081 = n35054 & ~n35080;
  assign n35082 = n35044 & n35081;
  assign n35083 = ~n34389 & n35057;
  assign n35084 = n34993 & n35083;
  assign n35085 = ~n35082 & ~n35084;
  assign n35086 = P1_BUF1_REG_30_ & n12494;
  assign n35087 = P1_BUF2_REG_30_ & ~n12494;
  assign n35088 = ~n35086 & ~n35087;
  assign n35089 = n35054 & ~n35088;
  assign n35090 = n35042 & n35089;
  assign n35091 = n35085 & ~n35090;
  assign n35092 = P1_BUF1_REG_6_ & n12494;
  assign n35093 = P1_BUF2_REG_6_ & ~n12494;
  assign n35094 = ~n35092 & ~n35093;
  assign n35095 = n34998 & ~n35094;
  assign n35096 = n35069 & n35095;
  assign n35097 = ~n35077 & n35091;
  assign n5866 = n35096 | ~n35097;
  assign n35099 = P1_P2_INSTQUEUE_REG_15__5_ & ~n35048;
  assign n35100 = P1_BUF1_REG_21_ & n12494;
  assign n35101 = P1_BUF2_REG_21_ & ~n12494;
  assign n35102 = ~n35100 & ~n35101;
  assign n35103 = n35054 & ~n35102;
  assign n35104 = n35044 & n35103;
  assign n35105 = ~n34358 & n35057;
  assign n35106 = n34993 & n35105;
  assign n35107 = ~n35104 & ~n35106;
  assign n35108 = P1_BUF1_REG_29_ & n12494;
  assign n35109 = P1_BUF2_REG_29_ & ~n12494;
  assign n35110 = ~n35108 & ~n35109;
  assign n35111 = n35054 & ~n35110;
  assign n35112 = n35042 & n35111;
  assign n35113 = n35107 & ~n35112;
  assign n35114 = P1_BUF1_REG_5_ & n12494;
  assign n35115 = P1_BUF2_REG_5_ & ~n12494;
  assign n35116 = ~n35114 & ~n35115;
  assign n35117 = n34998 & ~n35116;
  assign n35118 = n35069 & n35117;
  assign n35119 = ~n35099 & n35113;
  assign n5871 = n35118 | ~n35119;
  assign n35121 = P1_P2_INSTQUEUE_REG_15__4_ & ~n35048;
  assign n35122 = P1_BUF1_REG_20_ & n12494;
  assign n35123 = P1_BUF2_REG_20_ & ~n12494;
  assign n35124 = ~n35122 & ~n35123;
  assign n35125 = n35054 & ~n35124;
  assign n35126 = n35044 & n35125;
  assign n35127 = ~n34421 & n35057;
  assign n35128 = n34993 & n35127;
  assign n35129 = ~n35126 & ~n35128;
  assign n35130 = P1_BUF1_REG_28_ & n12494;
  assign n35131 = P1_BUF2_REG_28_ & ~n12494;
  assign n35132 = ~n35130 & ~n35131;
  assign n35133 = n35054 & ~n35132;
  assign n35134 = n35042 & n35133;
  assign n35135 = n35129 & ~n35134;
  assign n35136 = P1_BUF1_REG_4_ & n12494;
  assign n35137 = P1_BUF2_REG_4_ & ~n12494;
  assign n35138 = ~n35136 & ~n35137;
  assign n35139 = n34998 & ~n35138;
  assign n35140 = n35069 & n35139;
  assign n35141 = ~n35121 & n35135;
  assign n5876 = n35140 | ~n35141;
  assign n35143 = P1_P2_INSTQUEUE_REG_15__3_ & ~n35048;
  assign n35144 = P1_BUF1_REG_19_ & n12494;
  assign n35145 = P1_BUF2_REG_19_ & ~n12494;
  assign n35146 = ~n35144 & ~n35145;
  assign n35147 = n35054 & ~n35146;
  assign n35148 = n35044 & n35147;
  assign n35149 = ~n34483 & n35057;
  assign n35150 = n34993 & n35149;
  assign n35151 = ~n35148 & ~n35150;
  assign n35152 = P1_BUF1_REG_27_ & n12494;
  assign n35153 = P1_BUF2_REG_27_ & ~n12494;
  assign n35154 = ~n35152 & ~n35153;
  assign n35155 = n35054 & ~n35154;
  assign n35156 = n35042 & n35155;
  assign n35157 = n35151 & ~n35156;
  assign n35158 = P1_BUF1_REG_3_ & n12494;
  assign n35159 = P1_BUF2_REG_3_ & ~n12494;
  assign n35160 = ~n35158 & ~n35159;
  assign n35161 = n34998 & ~n35160;
  assign n35162 = n35069 & n35161;
  assign n35163 = ~n35143 & n35157;
  assign n5881 = n35162 | ~n35163;
  assign n35165 = P1_P2_INSTQUEUE_REG_15__2_ & ~n35048;
  assign n35166 = P1_BUF1_REG_18_ & n12494;
  assign n35167 = P1_BUF2_REG_18_ & ~n12494;
  assign n35168 = ~n35166 & ~n35167;
  assign n35169 = n35054 & ~n35168;
  assign n35170 = n35044 & n35169;
  assign n35171 = ~n34514 & n35057;
  assign n35172 = n34993 & n35171;
  assign n35173 = ~n35170 & ~n35172;
  assign n35174 = P1_BUF1_REG_26_ & n12494;
  assign n35175 = P1_BUF2_REG_26_ & ~n12494;
  assign n35176 = ~n35174 & ~n35175;
  assign n35177 = n35054 & ~n35176;
  assign n35178 = n35042 & n35177;
  assign n35179 = n35173 & ~n35178;
  assign n35180 = P1_BUF1_REG_2_ & n12494;
  assign n35181 = P1_BUF2_REG_2_ & ~n12494;
  assign n35182 = ~n35180 & ~n35181;
  assign n35183 = n34998 & ~n35182;
  assign n35184 = n35069 & n35183;
  assign n35185 = ~n35165 & n35179;
  assign n5886 = n35184 | ~n35185;
  assign n35187 = P1_P2_INSTQUEUE_REG_15__1_ & ~n35048;
  assign n35188 = P1_BUF1_REG_17_ & n12494;
  assign n35189 = P1_BUF2_REG_17_ & ~n12494;
  assign n35190 = ~n35188 & ~n35189;
  assign n35191 = n35054 & ~n35190;
  assign n35192 = n35044 & n35191;
  assign n35193 = ~n34549 & n35057;
  assign n35194 = n34993 & n35193;
  assign n35195 = ~n35192 & ~n35194;
  assign n35196 = P1_BUF1_REG_25_ & n12494;
  assign n35197 = P1_BUF2_REG_25_ & ~n12494;
  assign n35198 = ~n35196 & ~n35197;
  assign n35199 = n35054 & ~n35198;
  assign n35200 = n35042 & n35199;
  assign n35201 = n35195 & ~n35200;
  assign n35202 = P1_BUF1_REG_1_ & n12494;
  assign n35203 = P1_BUF2_REG_1_ & ~n12494;
  assign n35204 = ~n35202 & ~n35203;
  assign n35205 = n34998 & ~n35204;
  assign n35206 = n35069 & n35205;
  assign n35207 = ~n35187 & n35201;
  assign n5891 = n35206 | ~n35207;
  assign n35209 = P1_P2_INSTQUEUE_REG_15__0_ & ~n35048;
  assign n35210 = P1_BUF1_REG_16_ & n12494;
  assign n35211 = P1_BUF2_REG_16_ & ~n12494;
  assign n35212 = ~n35210 & ~n35211;
  assign n35213 = n35054 & ~n35212;
  assign n35214 = n35044 & n35213;
  assign n35215 = ~n34580 & n35057;
  assign n35216 = n34993 & n35215;
  assign n35217 = ~n35214 & ~n35216;
  assign n35218 = P1_BUF1_REG_24_ & n12494;
  assign n35219 = P1_BUF2_REG_24_ & ~n12494;
  assign n35220 = ~n35218 & ~n35219;
  assign n35221 = n35054 & ~n35220;
  assign n35222 = n35042 & n35221;
  assign n35223 = n35217 & ~n35222;
  assign n35224 = P1_BUF1_REG_0_ & n12494;
  assign n35225 = P1_BUF2_REG_0_ & ~n12494;
  assign n35226 = ~n35224 & ~n35225;
  assign n35227 = n34998 & ~n35226;
  assign n35228 = n35069 & n35227;
  assign n35229 = ~n35209 & n35223;
  assign n5896 = n35228 | ~n35229;
  assign n35231 = P1_P2_INSTQUEUEWR_ADDR_REG_3_ & P1_P2_INSTQUEUEWR_ADDR_REG_1_;
  assign n35232 = P1_P2_INSTQUEUEWR_ADDR_REG_2_ & ~P1_P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n35233 = n35231 & n35232;
  assign n35234 = P1_P2_STATE2_REG_3_ & ~n35233;
  assign n35235 = n34998 & ~n35234;
  assign n35236 = n35006 & n35016;
  assign n35237 = ~n35233 & ~n35236;
  assign n35238 = P1_P2_INSTQUEUEWR_ADDR_REG_0_ & ~n35021;
  assign n35239 = n35041 & n35238;
  assign n35240 = n35019 & n35043;
  assign n35241 = ~n35239 & ~n35240;
  assign n35242 = n35015 & ~n35241;
  assign n35243 = n35237 & ~n35242;
  assign n35244 = n35235 & ~n35243;
  assign n35245 = P1_P2_INSTQUEUE_REG_14__7_ & ~n35244;
  assign n35246 = n35055 & n35240;
  assign n35247 = n35058 & n35233;
  assign n35248 = ~n35246 & ~n35247;
  assign n35249 = n35064 & n35239;
  assign n35250 = n35248 & ~n35249;
  assign n35251 = n35053 & n35241;
  assign n35252 = n35015 & ~n35251;
  assign n35253 = ~n35237 & ~n35252;
  assign n35254 = n35073 & n35253;
  assign n35255 = ~n35245 & n35250;
  assign n5901 = n35254 | ~n35255;
  assign n35257 = P1_P2_INSTQUEUE_REG_14__6_ & ~n35244;
  assign n35258 = n35081 & n35240;
  assign n35259 = n35083 & n35233;
  assign n35260 = ~n35258 & ~n35259;
  assign n35261 = n35089 & n35239;
  assign n35262 = n35260 & ~n35261;
  assign n35263 = n35095 & n35253;
  assign n35264 = ~n35257 & n35262;
  assign n5906 = n35263 | ~n35264;
  assign n35266 = P1_P2_INSTQUEUE_REG_14__5_ & ~n35244;
  assign n35267 = n35103 & n35240;
  assign n35268 = n35105 & n35233;
  assign n35269 = ~n35267 & ~n35268;
  assign n35270 = n35111 & n35239;
  assign n35271 = n35269 & ~n35270;
  assign n35272 = n35117 & n35253;
  assign n35273 = ~n35266 & n35271;
  assign n5911 = n35272 | ~n35273;
  assign n35275 = P1_P2_INSTQUEUE_REG_14__4_ & ~n35244;
  assign n35276 = n35125 & n35240;
  assign n35277 = n35127 & n35233;
  assign n35278 = ~n35276 & ~n35277;
  assign n35279 = n35133 & n35239;
  assign n35280 = n35278 & ~n35279;
  assign n35281 = n35139 & n35253;
  assign n35282 = ~n35275 & n35280;
  assign n5916 = n35281 | ~n35282;
  assign n35284 = P1_P2_INSTQUEUE_REG_14__3_ & ~n35244;
  assign n35285 = n35147 & n35240;
  assign n35286 = n35149 & n35233;
  assign n35287 = ~n35285 & ~n35286;
  assign n35288 = n35155 & n35239;
  assign n35289 = n35287 & ~n35288;
  assign n35290 = n35161 & n35253;
  assign n35291 = ~n35284 & n35289;
  assign n5921 = n35290 | ~n35291;
  assign n35293 = P1_P2_INSTQUEUE_REG_14__2_ & ~n35244;
  assign n35294 = n35169 & n35240;
  assign n35295 = n35171 & n35233;
  assign n35296 = ~n35294 & ~n35295;
  assign n35297 = n35177 & n35239;
  assign n35298 = n35296 & ~n35297;
  assign n35299 = n35183 & n35253;
  assign n35300 = ~n35293 & n35298;
  assign n5926 = n35299 | ~n35300;
  assign n35302 = P1_P2_INSTQUEUE_REG_14__1_ & ~n35244;
  assign n35303 = n35191 & n35240;
  assign n35304 = n35193 & n35233;
  assign n35305 = ~n35303 & ~n35304;
  assign n35306 = n35199 & n35239;
  assign n35307 = n35305 & ~n35306;
  assign n35308 = n35205 & n35253;
  assign n35309 = ~n35302 & n35307;
  assign n5931 = n35308 | ~n35309;
  assign n35311 = P1_P2_INSTQUEUE_REG_14__0_ & ~n35244;
  assign n35312 = n35213 & n35240;
  assign n35313 = n35215 & n35233;
  assign n35314 = ~n35312 & ~n35313;
  assign n35315 = n35221 & n35239;
  assign n35316 = n35314 & ~n35315;
  assign n35317 = n35227 & n35253;
  assign n35318 = ~n35311 & n35316;
  assign n5936 = n35317 | ~n35318;
  assign n35320 = P1_P2_INSTQUEUEWR_ADDR_REG_3_ & P1_P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n35321 = n35007 & n35320;
  assign n35322 = P1_P2_STATE2_REG_3_ & ~n35321;
  assign n35323 = n34998 & ~n35322;
  assign n35324 = n35006 & n35017;
  assign n35325 = ~n35321 & ~n35324;
  assign n35326 = ~P1_P2_INSTQUEUEWR_ADDR_REG_0_ & n35021;
  assign n35327 = n35041 & n35326;
  assign n35328 = n35020 & n35043;
  assign n35329 = ~n35327 & ~n35328;
  assign n35330 = n35015 & ~n35329;
  assign n35331 = n35325 & ~n35330;
  assign n35332 = n35323 & ~n35331;
  assign n35333 = P1_P2_INSTQUEUE_REG_13__7_ & ~n35332;
  assign n35334 = n35055 & n35328;
  assign n35335 = n35058 & n35321;
  assign n35336 = ~n35334 & ~n35335;
  assign n35337 = n35064 & n35327;
  assign n35338 = n35336 & ~n35337;
  assign n35339 = n35053 & n35329;
  assign n35340 = n35015 & ~n35339;
  assign n35341 = ~n35325 & ~n35340;
  assign n35342 = n35073 & n35341;
  assign n35343 = ~n35333 & n35338;
  assign n5941 = n35342 | ~n35343;
  assign n35345 = P1_P2_INSTQUEUE_REG_13__6_ & ~n35332;
  assign n35346 = n35081 & n35328;
  assign n35347 = n35083 & n35321;
  assign n35348 = ~n35346 & ~n35347;
  assign n35349 = n35089 & n35327;
  assign n35350 = n35348 & ~n35349;
  assign n35351 = n35095 & n35341;
  assign n35352 = ~n35345 & n35350;
  assign n5946 = n35351 | ~n35352;
  assign n35354 = P1_P2_INSTQUEUE_REG_13__5_ & ~n35332;
  assign n35355 = n35103 & n35328;
  assign n35356 = n35105 & n35321;
  assign n35357 = ~n35355 & ~n35356;
  assign n35358 = n35111 & n35327;
  assign n35359 = n35357 & ~n35358;
  assign n35360 = n35117 & n35341;
  assign n35361 = ~n35354 & n35359;
  assign n5951 = n35360 | ~n35361;
  assign n35363 = P1_P2_INSTQUEUE_REG_13__4_ & ~n35332;
  assign n35364 = n35125 & n35328;
  assign n35365 = n35127 & n35321;
  assign n35366 = ~n35364 & ~n35365;
  assign n35367 = n35133 & n35327;
  assign n35368 = n35366 & ~n35367;
  assign n35369 = n35139 & n35341;
  assign n35370 = ~n35363 & n35368;
  assign n5956 = n35369 | ~n35370;
  assign n35372 = P1_P2_INSTQUEUE_REG_13__3_ & ~n35332;
  assign n35373 = n35147 & n35328;
  assign n35374 = n35149 & n35321;
  assign n35375 = ~n35373 & ~n35374;
  assign n35376 = n35155 & n35327;
  assign n35377 = n35375 & ~n35376;
  assign n35378 = n35161 & n35341;
  assign n35379 = ~n35372 & n35377;
  assign n5961 = n35378 | ~n35379;
  assign n35381 = P1_P2_INSTQUEUE_REG_13__2_ & ~n35332;
  assign n35382 = n35169 & n35328;
  assign n35383 = n35171 & n35321;
  assign n35384 = ~n35382 & ~n35383;
  assign n35385 = n35177 & n35327;
  assign n35386 = n35384 & ~n35385;
  assign n35387 = n35183 & n35341;
  assign n35388 = ~n35381 & n35386;
  assign n5966 = n35387 | ~n35388;
  assign n35390 = P1_P2_INSTQUEUE_REG_13__1_ & ~n35332;
  assign n35391 = n35191 & n35328;
  assign n35392 = n35193 & n35321;
  assign n35393 = ~n35391 & ~n35392;
  assign n35394 = n35199 & n35327;
  assign n35395 = n35393 & ~n35394;
  assign n35396 = n35205 & n35341;
  assign n35397 = ~n35390 & n35395;
  assign n5971 = n35396 | ~n35397;
  assign n35399 = P1_P2_INSTQUEUE_REG_13__0_ & ~n35332;
  assign n35400 = n35213 & n35328;
  assign n35401 = n35215 & n35321;
  assign n35402 = ~n35400 & ~n35401;
  assign n35403 = n35221 & n35327;
  assign n35404 = n35402 & ~n35403;
  assign n35405 = n35227 & n35341;
  assign n35406 = ~n35399 & n35404;
  assign n5976 = n35405 | ~n35406;
  assign n35408 = P1_P2_INSTQUEUEWR_ADDR_REG_3_ & ~P1_P2_INSTQUEUEWR_ADDR_REG_1_;
  assign n35409 = n35232 & n35408;
  assign n35410 = P1_P2_STATE2_REG_3_ & ~n35409;
  assign n35411 = n34998 & ~n35410;
  assign n35412 = P1_P2_INSTQUEUEWR_ADDR_REG_0_ & n35021;
  assign n35413 = n35041 & n35412;
  assign n35414 = ~P1_P2_INSTQUEUEWR_ADDR_REG_0_ & n35018;
  assign n35415 = n35043 & n35414;
  assign n35416 = ~n35413 & ~n35415;
  assign n35417 = n35015 & ~n35416;
  assign n35418 = n35006 & n35009;
  assign n35419 = ~n35417 & ~n35418;
  assign n35420 = n35411 & ~n35419;
  assign n35421 = P1_P2_INSTQUEUE_REG_12__7_ & ~n35420;
  assign n35422 = n35055 & n35415;
  assign n35423 = n35058 & n35409;
  assign n35424 = ~n35422 & ~n35423;
  assign n35425 = n35064 & n35413;
  assign n35426 = n35424 & ~n35425;
  assign n35427 = n35053 & n35416;
  assign n35428 = n35015 & ~n35427;
  assign n35429 = n35418 & ~n35428;
  assign n35430 = n35073 & n35429;
  assign n35431 = ~n35421 & n35426;
  assign n5981 = n35430 | ~n35431;
  assign n35433 = P1_P2_INSTQUEUE_REG_12__6_ & ~n35420;
  assign n35434 = n35081 & n35415;
  assign n35435 = n35083 & n35409;
  assign n35436 = ~n35434 & ~n35435;
  assign n35437 = n35089 & n35413;
  assign n35438 = n35436 & ~n35437;
  assign n35439 = n35095 & n35429;
  assign n35440 = ~n35433 & n35438;
  assign n5986 = n35439 | ~n35440;
  assign n35442 = P1_P2_INSTQUEUE_REG_12__5_ & ~n35420;
  assign n35443 = n35103 & n35415;
  assign n35444 = n35105 & n35409;
  assign n35445 = ~n35443 & ~n35444;
  assign n35446 = n35111 & n35413;
  assign n35447 = n35445 & ~n35446;
  assign n35448 = n35117 & n35429;
  assign n35449 = ~n35442 & n35447;
  assign n5991 = n35448 | ~n35449;
  assign n35451 = P1_P2_INSTQUEUE_REG_12__4_ & ~n35420;
  assign n35452 = n35125 & n35415;
  assign n35453 = n35127 & n35409;
  assign n35454 = ~n35452 & ~n35453;
  assign n35455 = n35133 & n35413;
  assign n35456 = n35454 & ~n35455;
  assign n35457 = n35139 & n35429;
  assign n35458 = ~n35451 & n35456;
  assign n5996 = n35457 | ~n35458;
  assign n35460 = P1_P2_INSTQUEUE_REG_12__3_ & ~n35420;
  assign n35461 = n35147 & n35415;
  assign n35462 = n35149 & n35409;
  assign n35463 = ~n35461 & ~n35462;
  assign n35464 = n35155 & n35413;
  assign n35465 = n35463 & ~n35464;
  assign n35466 = n35161 & n35429;
  assign n35467 = ~n35460 & n35465;
  assign n6001 = n35466 | ~n35467;
  assign n35469 = P1_P2_INSTQUEUE_REG_12__2_ & ~n35420;
  assign n35470 = n35169 & n35415;
  assign n35471 = n35171 & n35409;
  assign n35472 = ~n35470 & ~n35471;
  assign n35473 = n35177 & n35413;
  assign n35474 = n35472 & ~n35473;
  assign n35475 = n35183 & n35429;
  assign n35476 = ~n35469 & n35474;
  assign n6006 = n35475 | ~n35476;
  assign n35478 = P1_P2_INSTQUEUE_REG_12__1_ & ~n35420;
  assign n35479 = n35191 & n35415;
  assign n35480 = n35193 & n35409;
  assign n35481 = ~n35479 & ~n35480;
  assign n35482 = n35199 & n35413;
  assign n35483 = n35481 & ~n35482;
  assign n35484 = n35205 & n35429;
  assign n35485 = ~n35478 & n35483;
  assign n6011 = n35484 | ~n35485;
  assign n35487 = P1_P2_INSTQUEUE_REG_12__0_ & ~n35420;
  assign n35488 = n35213 & n35415;
  assign n35489 = n35215 & n35409;
  assign n35490 = ~n35488 & ~n35489;
  assign n35491 = n35221 & n35413;
  assign n35492 = n35490 & ~n35491;
  assign n35493 = n35227 & n35429;
  assign n35494 = ~n35487 & n35492;
  assign n6016 = n35493 | ~n35494;
  assign n35496 = P1_P2_INSTQUEUEWR_ADDR_REG_3_ & ~P1_P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n35497 = n34991 & n35496;
  assign n35498 = P1_P2_STATE2_REG_3_ & ~n35497;
  assign n35499 = n34998 & ~n35498;
  assign n35500 = n35002 & ~n35005;
  assign n35501 = n35010 & n35500;
  assign n35502 = ~n35497 & ~n35501;
  assign n35503 = n35029 & ~n35040;
  assign n35504 = n35022 & n35503;
  assign n35505 = n35026 & n35035;
  assign n35506 = ~n35504 & ~n35505;
  assign n35507 = n35015 & ~n35506;
  assign n35508 = n35502 & ~n35507;
  assign n35509 = n35499 & ~n35508;
  assign n35510 = P1_P2_INSTQUEUE_REG_11__7_ & ~n35509;
  assign n35511 = n35055 & n35505;
  assign n35512 = n35058 & n35497;
  assign n35513 = ~n35511 & ~n35512;
  assign n35514 = n35064 & n35504;
  assign n35515 = n35513 & ~n35514;
  assign n35516 = n35053 & n35506;
  assign n35517 = n35015 & ~n35516;
  assign n35518 = ~n35502 & ~n35517;
  assign n35519 = n35073 & n35518;
  assign n35520 = ~n35510 & n35515;
  assign n6021 = n35519 | ~n35520;
  assign n35522 = P1_P2_INSTQUEUE_REG_11__6_ & ~n35509;
  assign n35523 = n35081 & n35505;
  assign n35524 = n35083 & n35497;
  assign n35525 = ~n35523 & ~n35524;
  assign n35526 = n35089 & n35504;
  assign n35527 = n35525 & ~n35526;
  assign n35528 = n35095 & n35518;
  assign n35529 = ~n35522 & n35527;
  assign n6026 = n35528 | ~n35529;
  assign n35531 = P1_P2_INSTQUEUE_REG_11__5_ & ~n35509;
  assign n35532 = n35103 & n35505;
  assign n35533 = n35105 & n35497;
  assign n35534 = ~n35532 & ~n35533;
  assign n35535 = n35111 & n35504;
  assign n35536 = n35534 & ~n35535;
  assign n35537 = n35117 & n35518;
  assign n35538 = ~n35531 & n35536;
  assign n6031 = n35537 | ~n35538;
  assign n35540 = P1_P2_INSTQUEUE_REG_11__4_ & ~n35509;
  assign n35541 = n35125 & n35505;
  assign n35542 = n35127 & n35497;
  assign n35543 = ~n35541 & ~n35542;
  assign n35544 = n35133 & n35504;
  assign n35545 = n35543 & ~n35544;
  assign n35546 = n35139 & n35518;
  assign n35547 = ~n35540 & n35545;
  assign n6036 = n35546 | ~n35547;
  assign n35549 = P1_P2_INSTQUEUE_REG_11__3_ & ~n35509;
  assign n35550 = n35147 & n35505;
  assign n35551 = n35149 & n35497;
  assign n35552 = ~n35550 & ~n35551;
  assign n35553 = n35155 & n35504;
  assign n35554 = n35552 & ~n35553;
  assign n35555 = n35161 & n35518;
  assign n35556 = ~n35549 & n35554;
  assign n6041 = n35555 | ~n35556;
  assign n35558 = P1_P2_INSTQUEUE_REG_11__2_ & ~n35509;
  assign n35559 = n35169 & n35505;
  assign n35560 = n35171 & n35497;
  assign n35561 = ~n35559 & ~n35560;
  assign n35562 = n35177 & n35504;
  assign n35563 = n35561 & ~n35562;
  assign n35564 = n35183 & n35518;
  assign n35565 = ~n35558 & n35563;
  assign n6046 = n35564 | ~n35565;
  assign n35567 = P1_P2_INSTQUEUE_REG_11__1_ & ~n35509;
  assign n35568 = n35191 & n35505;
  assign n35569 = n35193 & n35497;
  assign n35570 = ~n35568 & ~n35569;
  assign n35571 = n35199 & n35504;
  assign n35572 = n35570 & ~n35571;
  assign n35573 = n35205 & n35518;
  assign n35574 = ~n35567 & n35572;
  assign n6051 = n35573 | ~n35574;
  assign n35576 = P1_P2_INSTQUEUE_REG_11__0_ & ~n35509;
  assign n35577 = n35213 & n35505;
  assign n35578 = n35215 & n35497;
  assign n35579 = ~n35577 & ~n35578;
  assign n35580 = n35221 & n35504;
  assign n35581 = n35579 & ~n35580;
  assign n35582 = n35227 & n35518;
  assign n35583 = ~n35576 & n35581;
  assign n6056 = n35582 | ~n35583;
  assign n35585 = ~P1_P2_INSTQUEUEWR_ADDR_REG_2_ & ~P1_P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n35586 = n35231 & n35585;
  assign n35587 = P1_P2_STATE2_REG_3_ & ~n35586;
  assign n35588 = n34998 & ~n35587;
  assign n35589 = n35016 & n35500;
  assign n35590 = ~n35586 & ~n35589;
  assign n35591 = n35238 & n35503;
  assign n35592 = n35019 & n35035;
  assign n35593 = ~n35591 & ~n35592;
  assign n35594 = n35015 & ~n35593;
  assign n35595 = n35590 & ~n35594;
  assign n35596 = n35588 & ~n35595;
  assign n35597 = P1_P2_INSTQUEUE_REG_10__7_ & ~n35596;
  assign n35598 = n35055 & n35592;
  assign n35599 = n35058 & n35586;
  assign n35600 = ~n35598 & ~n35599;
  assign n35601 = n35064 & n35591;
  assign n35602 = n35600 & ~n35601;
  assign n35603 = n35053 & n35593;
  assign n35604 = n35015 & ~n35603;
  assign n35605 = ~n35590 & ~n35604;
  assign n35606 = n35073 & n35605;
  assign n35607 = ~n35597 & n35602;
  assign n6061 = n35606 | ~n35607;
  assign n35609 = P1_P2_INSTQUEUE_REG_10__6_ & ~n35596;
  assign n35610 = n35081 & n35592;
  assign n35611 = n35083 & n35586;
  assign n35612 = ~n35610 & ~n35611;
  assign n35613 = n35089 & n35591;
  assign n35614 = n35612 & ~n35613;
  assign n35615 = n35095 & n35605;
  assign n35616 = ~n35609 & n35614;
  assign n6066 = n35615 | ~n35616;
  assign n35618 = P1_P2_INSTQUEUE_REG_10__5_ & ~n35596;
  assign n35619 = n35103 & n35592;
  assign n35620 = n35105 & n35586;
  assign n35621 = ~n35619 & ~n35620;
  assign n35622 = n35111 & n35591;
  assign n35623 = n35621 & ~n35622;
  assign n35624 = n35117 & n35605;
  assign n35625 = ~n35618 & n35623;
  assign n6071 = n35624 | ~n35625;
  assign n35627 = P1_P2_INSTQUEUE_REG_10__4_ & ~n35596;
  assign n35628 = n35125 & n35592;
  assign n35629 = n35127 & n35586;
  assign n35630 = ~n35628 & ~n35629;
  assign n35631 = n35133 & n35591;
  assign n35632 = n35630 & ~n35631;
  assign n35633 = n35139 & n35605;
  assign n35634 = ~n35627 & n35632;
  assign n6076 = n35633 | ~n35634;
  assign n35636 = P1_P2_INSTQUEUE_REG_10__3_ & ~n35596;
  assign n35637 = n35147 & n35592;
  assign n35638 = n35149 & n35586;
  assign n35639 = ~n35637 & ~n35638;
  assign n35640 = n35155 & n35591;
  assign n35641 = n35639 & ~n35640;
  assign n35642 = n35161 & n35605;
  assign n35643 = ~n35636 & n35641;
  assign n6081 = n35642 | ~n35643;
  assign n35645 = P1_P2_INSTQUEUE_REG_10__2_ & ~n35596;
  assign n35646 = n35169 & n35592;
  assign n35647 = n35171 & n35586;
  assign n35648 = ~n35646 & ~n35647;
  assign n35649 = n35177 & n35591;
  assign n35650 = n35648 & ~n35649;
  assign n35651 = n35183 & n35605;
  assign n35652 = ~n35645 & n35650;
  assign n6086 = n35651 | ~n35652;
  assign n35654 = P1_P2_INSTQUEUE_REG_10__1_ & ~n35596;
  assign n35655 = n35191 & n35592;
  assign n35656 = n35193 & n35586;
  assign n35657 = ~n35655 & ~n35656;
  assign n35658 = n35199 & n35591;
  assign n35659 = n35657 & ~n35658;
  assign n35660 = n35205 & n35605;
  assign n35661 = ~n35654 & n35659;
  assign n6091 = n35660 | ~n35661;
  assign n35663 = P1_P2_INSTQUEUE_REG_10__0_ & ~n35596;
  assign n35664 = n35213 & n35592;
  assign n35665 = n35215 & n35586;
  assign n35666 = ~n35664 & ~n35665;
  assign n35667 = n35221 & n35591;
  assign n35668 = n35666 & ~n35667;
  assign n35669 = n35227 & n35605;
  assign n35670 = ~n35663 & n35668;
  assign n6096 = n35669 | ~n35670;
  assign n35672 = n35007 & n35496;
  assign n35673 = P1_P2_STATE2_REG_3_ & ~n35672;
  assign n35674 = n34998 & ~n35673;
  assign n35675 = n35017 & n35500;
  assign n35676 = ~n35672 & ~n35675;
  assign n35677 = n35326 & n35503;
  assign n35678 = n35020 & n35035;
  assign n35679 = ~n35677 & ~n35678;
  assign n35680 = n35015 & ~n35679;
  assign n35681 = n35676 & ~n35680;
  assign n35682 = n35674 & ~n35681;
  assign n35683 = P1_P2_INSTQUEUE_REG_9__7_ & ~n35682;
  assign n35684 = n35055 & n35678;
  assign n35685 = n35058 & n35672;
  assign n35686 = ~n35684 & ~n35685;
  assign n35687 = n35064 & n35677;
  assign n35688 = n35686 & ~n35687;
  assign n35689 = n35053 & n35679;
  assign n35690 = n35015 & ~n35689;
  assign n35691 = ~n35676 & ~n35690;
  assign n35692 = n35073 & n35691;
  assign n35693 = ~n35683 & n35688;
  assign n6101 = n35692 | ~n35693;
  assign n35695 = P1_P2_INSTQUEUE_REG_9__6_ & ~n35682;
  assign n35696 = n35081 & n35678;
  assign n35697 = n35083 & n35672;
  assign n35698 = ~n35696 & ~n35697;
  assign n35699 = n35089 & n35677;
  assign n35700 = n35698 & ~n35699;
  assign n35701 = n35095 & n35691;
  assign n35702 = ~n35695 & n35700;
  assign n6106 = n35701 | ~n35702;
  assign n35704 = P1_P2_INSTQUEUE_REG_9__5_ & ~n35682;
  assign n35705 = n35103 & n35678;
  assign n35706 = n35105 & n35672;
  assign n35707 = ~n35705 & ~n35706;
  assign n35708 = n35111 & n35677;
  assign n35709 = n35707 & ~n35708;
  assign n35710 = n35117 & n35691;
  assign n35711 = ~n35704 & n35709;
  assign n6111 = n35710 | ~n35711;
  assign n35713 = P1_P2_INSTQUEUE_REG_9__4_ & ~n35682;
  assign n35714 = n35125 & n35678;
  assign n35715 = n35127 & n35672;
  assign n35716 = ~n35714 & ~n35715;
  assign n35717 = n35133 & n35677;
  assign n35718 = n35716 & ~n35717;
  assign n35719 = n35139 & n35691;
  assign n35720 = ~n35713 & n35718;
  assign n6116 = n35719 | ~n35720;
  assign n35722 = P1_P2_INSTQUEUE_REG_9__3_ & ~n35682;
  assign n35723 = n35147 & n35678;
  assign n35724 = n35149 & n35672;
  assign n35725 = ~n35723 & ~n35724;
  assign n35726 = n35155 & n35677;
  assign n35727 = n35725 & ~n35726;
  assign n35728 = n35161 & n35691;
  assign n35729 = ~n35722 & n35727;
  assign n6121 = n35728 | ~n35729;
  assign n35731 = P1_P2_INSTQUEUE_REG_9__2_ & ~n35682;
  assign n35732 = n35169 & n35678;
  assign n35733 = n35171 & n35672;
  assign n35734 = ~n35732 & ~n35733;
  assign n35735 = n35177 & n35677;
  assign n35736 = n35734 & ~n35735;
  assign n35737 = n35183 & n35691;
  assign n35738 = ~n35731 & n35736;
  assign n6126 = n35737 | ~n35738;
  assign n35740 = P1_P2_INSTQUEUE_REG_9__1_ & ~n35682;
  assign n35741 = n35191 & n35678;
  assign n35742 = n35193 & n35672;
  assign n35743 = ~n35741 & ~n35742;
  assign n35744 = n35199 & n35677;
  assign n35745 = n35743 & ~n35744;
  assign n35746 = n35205 & n35691;
  assign n35747 = ~n35740 & n35745;
  assign n6131 = n35746 | ~n35747;
  assign n35749 = P1_P2_INSTQUEUE_REG_9__0_ & ~n35682;
  assign n35750 = n35213 & n35678;
  assign n35751 = n35215 & n35672;
  assign n35752 = ~n35750 & ~n35751;
  assign n35753 = n35221 & n35677;
  assign n35754 = n35752 & ~n35753;
  assign n35755 = n35227 & n35691;
  assign n35756 = ~n35749 & n35754;
  assign n6136 = n35755 | ~n35756;
  assign n35758 = n35408 & n35585;
  assign n35759 = P1_P2_STATE2_REG_3_ & ~n35758;
  assign n35760 = n34998 & ~n35759;
  assign n35761 = n35412 & n35503;
  assign n35762 = n35035 & n35414;
  assign n35763 = ~n35761 & ~n35762;
  assign n35764 = n35015 & ~n35763;
  assign n35765 = n35009 & n35500;
  assign n35766 = ~n35764 & ~n35765;
  assign n35767 = n35760 & ~n35766;
  assign n35768 = P1_P2_INSTQUEUE_REG_8__7_ & ~n35767;
  assign n35769 = n35055 & n35762;
  assign n35770 = n35058 & n35758;
  assign n35771 = ~n35769 & ~n35770;
  assign n35772 = n35064 & n35761;
  assign n35773 = n35771 & ~n35772;
  assign n35774 = n35053 & n35763;
  assign n35775 = n35015 & ~n35774;
  assign n35776 = n35765 & ~n35775;
  assign n35777 = n35073 & n35776;
  assign n35778 = ~n35768 & n35773;
  assign n6141 = n35777 | ~n35778;
  assign n35780 = P1_P2_INSTQUEUE_REG_8__6_ & ~n35767;
  assign n35781 = n35081 & n35762;
  assign n35782 = n35083 & n35758;
  assign n35783 = ~n35781 & ~n35782;
  assign n35784 = n35089 & n35761;
  assign n35785 = n35783 & ~n35784;
  assign n35786 = n35095 & n35776;
  assign n35787 = ~n35780 & n35785;
  assign n6146 = n35786 | ~n35787;
  assign n35789 = P1_P2_INSTQUEUE_REG_8__5_ & ~n35767;
  assign n35790 = n35103 & n35762;
  assign n35791 = n35105 & n35758;
  assign n35792 = ~n35790 & ~n35791;
  assign n35793 = n35111 & n35761;
  assign n35794 = n35792 & ~n35793;
  assign n35795 = n35117 & n35776;
  assign n35796 = ~n35789 & n35794;
  assign n6151 = n35795 | ~n35796;
  assign n35798 = P1_P2_INSTQUEUE_REG_8__4_ & ~n35767;
  assign n35799 = n35125 & n35762;
  assign n35800 = n35127 & n35758;
  assign n35801 = ~n35799 & ~n35800;
  assign n35802 = n35133 & n35761;
  assign n35803 = n35801 & ~n35802;
  assign n35804 = n35139 & n35776;
  assign n35805 = ~n35798 & n35803;
  assign n6156 = n35804 | ~n35805;
  assign n35807 = P1_P2_INSTQUEUE_REG_8__3_ & ~n35767;
  assign n35808 = n35147 & n35762;
  assign n35809 = n35149 & n35758;
  assign n35810 = ~n35808 & ~n35809;
  assign n35811 = n35155 & n35761;
  assign n35812 = n35810 & ~n35811;
  assign n35813 = n35161 & n35776;
  assign n35814 = ~n35807 & n35812;
  assign n6161 = n35813 | ~n35814;
  assign n35816 = P1_P2_INSTQUEUE_REG_8__2_ & ~n35767;
  assign n35817 = n35169 & n35762;
  assign n35818 = n35171 & n35758;
  assign n35819 = ~n35817 & ~n35818;
  assign n35820 = n35177 & n35761;
  assign n35821 = n35819 & ~n35820;
  assign n35822 = n35183 & n35776;
  assign n35823 = ~n35816 & n35821;
  assign n6166 = n35822 | ~n35823;
  assign n35825 = P1_P2_INSTQUEUE_REG_8__1_ & ~n35767;
  assign n35826 = n35191 & n35762;
  assign n35827 = n35193 & n35758;
  assign n35828 = ~n35826 & ~n35827;
  assign n35829 = n35199 & n35761;
  assign n35830 = n35828 & ~n35829;
  assign n35831 = n35205 & n35776;
  assign n35832 = ~n35825 & n35830;
  assign n6171 = n35831 | ~n35832;
  assign n35834 = P1_P2_INSTQUEUE_REG_8__0_ & ~n35767;
  assign n35835 = n35213 & n35762;
  assign n35836 = n35215 & n35758;
  assign n35837 = ~n35835 & ~n35836;
  assign n35838 = n35221 & n35761;
  assign n35839 = n35837 & ~n35838;
  assign n35840 = n35227 & n35776;
  assign n35841 = ~n35834 & n35839;
  assign n6176 = n35840 | ~n35841;
  assign n35843 = P1_P2_STATE2_REG_3_ & ~n35003;
  assign n35844 = n34998 & ~n35843;
  assign n35845 = ~n35003 & ~n35031;
  assign n35846 = ~n35029 & n35040;
  assign n35847 = n35022 & n35846;
  assign n35848 = ~n35039 & ~n35847;
  assign n35849 = n35015 & ~n35848;
  assign n35850 = n35845 & ~n35849;
  assign n35851 = n35844 & ~n35850;
  assign n35852 = P1_P2_INSTQUEUE_REG_7__7_ & ~n35851;
  assign n35853 = n35039 & n35055;
  assign n35854 = n35003 & n35058;
  assign n35855 = ~n35853 & ~n35854;
  assign n35856 = n35064 & n35847;
  assign n35857 = n35855 & ~n35856;
  assign n35858 = n35053 & n35848;
  assign n35859 = n35015 & ~n35858;
  assign n35860 = ~n35845 & ~n35859;
  assign n35861 = n35073 & n35860;
  assign n35862 = ~n35852 & n35857;
  assign n6181 = n35861 | ~n35862;
  assign n35864 = P1_P2_INSTQUEUE_REG_7__6_ & ~n35851;
  assign n35865 = n35039 & n35081;
  assign n35866 = n35003 & n35083;
  assign n35867 = ~n35865 & ~n35866;
  assign n35868 = n35089 & n35847;
  assign n35869 = n35867 & ~n35868;
  assign n35870 = n35095 & n35860;
  assign n35871 = ~n35864 & n35869;
  assign n6186 = n35870 | ~n35871;
  assign n35873 = P1_P2_INSTQUEUE_REG_7__5_ & ~n35851;
  assign n35874 = n35039 & n35103;
  assign n35875 = n35003 & n35105;
  assign n35876 = ~n35874 & ~n35875;
  assign n35877 = n35111 & n35847;
  assign n35878 = n35876 & ~n35877;
  assign n35879 = n35117 & n35860;
  assign n35880 = ~n35873 & n35878;
  assign n6191 = n35879 | ~n35880;
  assign n35882 = P1_P2_INSTQUEUE_REG_7__4_ & ~n35851;
  assign n35883 = n35039 & n35125;
  assign n35884 = n35003 & n35127;
  assign n35885 = ~n35883 & ~n35884;
  assign n35886 = n35133 & n35847;
  assign n35887 = n35885 & ~n35886;
  assign n35888 = n35139 & n35860;
  assign n35889 = ~n35882 & n35887;
  assign n6196 = n35888 | ~n35889;
  assign n35891 = P1_P2_INSTQUEUE_REG_7__3_ & ~n35851;
  assign n35892 = n35039 & n35147;
  assign n35893 = n35003 & n35149;
  assign n35894 = ~n35892 & ~n35893;
  assign n35895 = n35155 & n35847;
  assign n35896 = n35894 & ~n35895;
  assign n35897 = n35161 & n35860;
  assign n35898 = ~n35891 & n35896;
  assign n6201 = n35897 | ~n35898;
  assign n35900 = P1_P2_INSTQUEUE_REG_7__2_ & ~n35851;
  assign n35901 = n35039 & n35169;
  assign n35902 = n35003 & n35171;
  assign n35903 = ~n35901 & ~n35902;
  assign n35904 = n35177 & n35847;
  assign n35905 = n35903 & ~n35904;
  assign n35906 = n35183 & n35860;
  assign n35907 = ~n35900 & n35905;
  assign n6206 = n35906 | ~n35907;
  assign n35909 = P1_P2_INSTQUEUE_REG_7__1_ & ~n35851;
  assign n35910 = n35039 & n35191;
  assign n35911 = n35003 & n35193;
  assign n35912 = ~n35910 & ~n35911;
  assign n35913 = n35199 & n35847;
  assign n35914 = n35912 & ~n35913;
  assign n35915 = n35205 & n35860;
  assign n35916 = ~n35909 & n35914;
  assign n6211 = n35915 | ~n35916;
  assign n35918 = P1_P2_INSTQUEUE_REG_7__0_ & ~n35851;
  assign n35919 = n35039 & n35213;
  assign n35920 = n35003 & n35215;
  assign n35921 = ~n35919 & ~n35920;
  assign n35922 = n35221 & n35847;
  assign n35923 = n35921 & ~n35922;
  assign n35924 = n35227 & n35860;
  assign n35925 = ~n35918 & n35923;
  assign n6216 = n35924 | ~n35925;
  assign n35927 = ~P1_P2_INSTQUEUEWR_ADDR_REG_3_ & P1_P2_INSTQUEUEWR_ADDR_REG_1_;
  assign n35928 = n35232 & n35927;
  assign n35929 = P1_P2_STATE2_REG_3_ & ~n35928;
  assign n35930 = n34998 & ~n35929;
  assign n35931 = n35016 & n35030;
  assign n35932 = ~n35928 & ~n35931;
  assign n35933 = n35238 & n35846;
  assign n35934 = n35019 & n35038;
  assign n35935 = ~n35933 & ~n35934;
  assign n35936 = n35015 & ~n35935;
  assign n35937 = n35932 & ~n35936;
  assign n35938 = n35930 & ~n35937;
  assign n35939 = P1_P2_INSTQUEUE_REG_6__7_ & ~n35938;
  assign n35940 = n35055 & n35934;
  assign n35941 = n35058 & n35928;
  assign n35942 = ~n35940 & ~n35941;
  assign n35943 = n35064 & n35933;
  assign n35944 = n35942 & ~n35943;
  assign n35945 = n35053 & n35935;
  assign n35946 = n35015 & ~n35945;
  assign n35947 = ~n35932 & ~n35946;
  assign n35948 = n35073 & n35947;
  assign n35949 = ~n35939 & n35944;
  assign n6221 = n35948 | ~n35949;
  assign n35951 = P1_P2_INSTQUEUE_REG_6__6_ & ~n35938;
  assign n35952 = n35081 & n35934;
  assign n35953 = n35083 & n35928;
  assign n35954 = ~n35952 & ~n35953;
  assign n35955 = n35089 & n35933;
  assign n35956 = n35954 & ~n35955;
  assign n35957 = n35095 & n35947;
  assign n35958 = ~n35951 & n35956;
  assign n6226 = n35957 | ~n35958;
  assign n35960 = P1_P2_INSTQUEUE_REG_6__5_ & ~n35938;
  assign n35961 = n35103 & n35934;
  assign n35962 = n35105 & n35928;
  assign n35963 = ~n35961 & ~n35962;
  assign n35964 = n35111 & n35933;
  assign n35965 = n35963 & ~n35964;
  assign n35966 = n35117 & n35947;
  assign n35967 = ~n35960 & n35965;
  assign n6231 = n35966 | ~n35967;
  assign n35969 = P1_P2_INSTQUEUE_REG_6__4_ & ~n35938;
  assign n35970 = n35125 & n35934;
  assign n35971 = n35127 & n35928;
  assign n35972 = ~n35970 & ~n35971;
  assign n35973 = n35133 & n35933;
  assign n35974 = n35972 & ~n35973;
  assign n35975 = n35139 & n35947;
  assign n35976 = ~n35969 & n35974;
  assign n6236 = n35975 | ~n35976;
  assign n35978 = P1_P2_INSTQUEUE_REG_6__3_ & ~n35938;
  assign n35979 = n35147 & n35934;
  assign n35980 = n35149 & n35928;
  assign n35981 = ~n35979 & ~n35980;
  assign n35982 = n35155 & n35933;
  assign n35983 = n35981 & ~n35982;
  assign n35984 = n35161 & n35947;
  assign n35985 = ~n35978 & n35983;
  assign n6241 = n35984 | ~n35985;
  assign n35987 = P1_P2_INSTQUEUE_REG_6__2_ & ~n35938;
  assign n35988 = n35169 & n35934;
  assign n35989 = n35171 & n35928;
  assign n35990 = ~n35988 & ~n35989;
  assign n35991 = n35177 & n35933;
  assign n35992 = n35990 & ~n35991;
  assign n35993 = n35183 & n35947;
  assign n35994 = ~n35987 & n35992;
  assign n6246 = n35993 | ~n35994;
  assign n35996 = P1_P2_INSTQUEUE_REG_6__1_ & ~n35938;
  assign n35997 = n35191 & n35934;
  assign n35998 = n35193 & n35928;
  assign n35999 = ~n35997 & ~n35998;
  assign n36000 = n35199 & n35933;
  assign n36001 = n35999 & ~n36000;
  assign n36002 = n35205 & n35947;
  assign n36003 = ~n35996 & n36001;
  assign n6251 = n36002 | ~n36003;
  assign n36005 = P1_P2_INSTQUEUE_REG_6__0_ & ~n35938;
  assign n36006 = n35213 & n35934;
  assign n36007 = n35215 & n35928;
  assign n36008 = ~n36006 & ~n36007;
  assign n36009 = n35221 & n35933;
  assign n36010 = n36008 & ~n36009;
  assign n36011 = n35227 & n35947;
  assign n36012 = ~n36005 & n36010;
  assign n6256 = n36011 | ~n36012;
  assign n36014 = ~P1_P2_INSTQUEUEWR_ADDR_REG_3_ & P1_P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n36015 = n35007 & n36014;
  assign n36016 = P1_P2_STATE2_REG_3_ & ~n36015;
  assign n36017 = n34998 & ~n36016;
  assign n36018 = n35017 & n35030;
  assign n36019 = ~n36015 & ~n36018;
  assign n36020 = n35326 & n35846;
  assign n36021 = n35020 & n35038;
  assign n36022 = ~n36020 & ~n36021;
  assign n36023 = n35015 & ~n36022;
  assign n36024 = n36019 & ~n36023;
  assign n36025 = n36017 & ~n36024;
  assign n36026 = P1_P2_INSTQUEUE_REG_5__7_ & ~n36025;
  assign n36027 = n35055 & n36021;
  assign n36028 = n35058 & n36015;
  assign n36029 = ~n36027 & ~n36028;
  assign n36030 = n35064 & n36020;
  assign n36031 = n36029 & ~n36030;
  assign n36032 = n35053 & n36022;
  assign n36033 = n35015 & ~n36032;
  assign n36034 = ~n36019 & ~n36033;
  assign n36035 = n35073 & n36034;
  assign n36036 = ~n36026 & n36031;
  assign n6261 = n36035 | ~n36036;
  assign n36038 = P1_P2_INSTQUEUE_REG_5__6_ & ~n36025;
  assign n36039 = n35081 & n36021;
  assign n36040 = n35083 & n36015;
  assign n36041 = ~n36039 & ~n36040;
  assign n36042 = n35089 & n36020;
  assign n36043 = n36041 & ~n36042;
  assign n36044 = n35095 & n36034;
  assign n36045 = ~n36038 & n36043;
  assign n6266 = n36044 | ~n36045;
  assign n36047 = P1_P2_INSTQUEUE_REG_5__5_ & ~n36025;
  assign n36048 = n35103 & n36021;
  assign n36049 = n35105 & n36015;
  assign n36050 = ~n36048 & ~n36049;
  assign n36051 = n35111 & n36020;
  assign n36052 = n36050 & ~n36051;
  assign n36053 = n35117 & n36034;
  assign n36054 = ~n36047 & n36052;
  assign n6271 = n36053 | ~n36054;
  assign n36056 = P1_P2_INSTQUEUE_REG_5__4_ & ~n36025;
  assign n36057 = n35125 & n36021;
  assign n36058 = n35127 & n36015;
  assign n36059 = ~n36057 & ~n36058;
  assign n36060 = n35133 & n36020;
  assign n36061 = n36059 & ~n36060;
  assign n36062 = n35139 & n36034;
  assign n36063 = ~n36056 & n36061;
  assign n6276 = n36062 | ~n36063;
  assign n36065 = P1_P2_INSTQUEUE_REG_5__3_ & ~n36025;
  assign n36066 = n35147 & n36021;
  assign n36067 = n35149 & n36015;
  assign n36068 = ~n36066 & ~n36067;
  assign n36069 = n35155 & n36020;
  assign n36070 = n36068 & ~n36069;
  assign n36071 = n35161 & n36034;
  assign n36072 = ~n36065 & n36070;
  assign n6281 = n36071 | ~n36072;
  assign n36074 = P1_P2_INSTQUEUE_REG_5__2_ & ~n36025;
  assign n36075 = n35169 & n36021;
  assign n36076 = n35171 & n36015;
  assign n36077 = ~n36075 & ~n36076;
  assign n36078 = n35177 & n36020;
  assign n36079 = n36077 & ~n36078;
  assign n36080 = n35183 & n36034;
  assign n36081 = ~n36074 & n36079;
  assign n6286 = n36080 | ~n36081;
  assign n36083 = P1_P2_INSTQUEUE_REG_5__1_ & ~n36025;
  assign n36084 = n35191 & n36021;
  assign n36085 = n35193 & n36015;
  assign n36086 = ~n36084 & ~n36085;
  assign n36087 = n35199 & n36020;
  assign n36088 = n36086 & ~n36087;
  assign n36089 = n35205 & n36034;
  assign n36090 = ~n36083 & n36088;
  assign n6291 = n36089 | ~n36090;
  assign n36092 = P1_P2_INSTQUEUE_REG_5__0_ & ~n36025;
  assign n36093 = n35213 & n36021;
  assign n36094 = n35215 & n36015;
  assign n36095 = ~n36093 & ~n36094;
  assign n36096 = n35221 & n36020;
  assign n36097 = n36095 & ~n36096;
  assign n36098 = n35227 & n36034;
  assign n36099 = ~n36092 & n36097;
  assign n6296 = n36098 | ~n36099;
  assign n36101 = n35038 & n35414;
  assign n36102 = n35055 & n36101;
  assign n36103 = ~P1_P2_INSTQUEUEWR_ADDR_REG_3_ & ~P1_P2_INSTQUEUEWR_ADDR_REG_1_;
  assign n36104 = n35232 & n36103;
  assign n36105 = n35058 & n36104;
  assign n36106 = n35015 & ~n35053;
  assign n36107 = n35009 & n35030;
  assign n36108 = ~n36106 & n36107;
  assign n36109 = n35073 & n36108;
  assign n36110 = ~n36102 & ~n36105;
  assign n36111 = ~n36109 & n36110;
  assign n36112 = n35412 & n35846;
  assign n36113 = n35064 & n36112;
  assign n36114 = n36111 & ~n36113;
  assign n36115 = P1_P2_STATE2_REG_3_ & ~n36104;
  assign n36116 = n34998 & ~n36115;
  assign n36117 = ~n36101 & ~n36112;
  assign n36118 = n35015 & ~n36117;
  assign n36119 = ~n36107 & ~n36118;
  assign n36120 = n36116 & ~n36119;
  assign n36121 = P1_P2_INSTQUEUE_REG_4__7_ & ~n36120;
  assign n6301 = ~n36114 | n36121;
  assign n36123 = n35081 & n36101;
  assign n36124 = n35083 & n36104;
  assign n36125 = n35095 & n36108;
  assign n36126 = ~n36123 & ~n36124;
  assign n36127 = ~n36125 & n36126;
  assign n36128 = n35089 & n36112;
  assign n36129 = n36127 & ~n36128;
  assign n36130 = P1_P2_INSTQUEUE_REG_4__6_ & ~n36120;
  assign n6306 = ~n36129 | n36130;
  assign n36132 = n35103 & n36101;
  assign n36133 = n35105 & n36104;
  assign n36134 = n35117 & n36108;
  assign n36135 = ~n36132 & ~n36133;
  assign n36136 = ~n36134 & n36135;
  assign n36137 = n35111 & n36112;
  assign n36138 = n36136 & ~n36137;
  assign n36139 = P1_P2_INSTQUEUE_REG_4__5_ & ~n36120;
  assign n6311 = ~n36138 | n36139;
  assign n36141 = n35125 & n36101;
  assign n36142 = n35127 & n36104;
  assign n36143 = n35139 & n36108;
  assign n36144 = ~n36141 & ~n36142;
  assign n36145 = ~n36143 & n36144;
  assign n36146 = n35133 & n36112;
  assign n36147 = n36145 & ~n36146;
  assign n36148 = P1_P2_INSTQUEUE_REG_4__4_ & ~n36120;
  assign n6316 = ~n36147 | n36148;
  assign n36150 = n35147 & n36101;
  assign n36151 = n35149 & n36104;
  assign n36152 = n35161 & n36108;
  assign n36153 = ~n36150 & ~n36151;
  assign n36154 = ~n36152 & n36153;
  assign n36155 = n35155 & n36112;
  assign n36156 = n36154 & ~n36155;
  assign n36157 = P1_P2_INSTQUEUE_REG_4__3_ & ~n36120;
  assign n6321 = ~n36156 | n36157;
  assign n36159 = n35169 & n36101;
  assign n36160 = n35171 & n36104;
  assign n36161 = n35183 & n36108;
  assign n36162 = ~n36159 & ~n36160;
  assign n36163 = ~n36161 & n36162;
  assign n36164 = n35177 & n36112;
  assign n36165 = n36163 & ~n36164;
  assign n36166 = P1_P2_INSTQUEUE_REG_4__2_ & ~n36120;
  assign n6326 = ~n36165 | n36166;
  assign n36168 = n35191 & n36101;
  assign n36169 = n35193 & n36104;
  assign n36170 = n35205 & n36108;
  assign n36171 = ~n36168 & ~n36169;
  assign n36172 = ~n36170 & n36171;
  assign n36173 = n35199 & n36112;
  assign n36174 = n36172 & ~n36173;
  assign n36175 = P1_P2_INSTQUEUE_REG_4__1_ & ~n36120;
  assign n6331 = ~n36174 | n36175;
  assign n36177 = n35213 & n36101;
  assign n36178 = n35215 & n36104;
  assign n36179 = n35227 & n36108;
  assign n36180 = ~n36177 & ~n36178;
  assign n36181 = ~n36179 & n36180;
  assign n36182 = n35221 & n36112;
  assign n36183 = n36181 & ~n36182;
  assign n36184 = P1_P2_INSTQUEUE_REG_4__0_ & ~n36120;
  assign n6336 = ~n36183 | n36184;
  assign n36186 = n35025 & n35034;
  assign n36187 = n35026 & n36186;
  assign n36188 = n35055 & n36187;
  assign n36189 = ~P1_P2_INSTQUEUEWR_ADDR_REG_3_ & ~P1_P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n36190 = n34991 & n36189;
  assign n36191 = n35058 & n36190;
  assign n36192 = n35002 & n35005;
  assign n36193 = n35010 & n36192;
  assign n36194 = ~n36190 & ~n36193;
  assign n36195 = ~n36106 & ~n36194;
  assign n36196 = n35073 & n36195;
  assign n36197 = ~n36188 & ~n36191;
  assign n36198 = ~n36196 & n36197;
  assign n36199 = n35029 & n35040;
  assign n36200 = n35022 & n36199;
  assign n36201 = n35064 & n36200;
  assign n36202 = n36198 & ~n36201;
  assign n36203 = P1_P2_STATE2_REG_3_ & ~n36190;
  assign n36204 = n34998 & ~n36203;
  assign n36205 = ~n36187 & ~n36200;
  assign n36206 = n35015 & ~n36205;
  assign n36207 = n36194 & ~n36206;
  assign n36208 = n36204 & ~n36207;
  assign n36209 = P1_P2_INSTQUEUE_REG_3__7_ & ~n36208;
  assign n6341 = ~n36202 | n36209;
  assign n36211 = n35081 & n36187;
  assign n36212 = n35083 & n36190;
  assign n36213 = n35095 & n36195;
  assign n36214 = ~n36211 & ~n36212;
  assign n36215 = ~n36213 & n36214;
  assign n36216 = n35089 & n36200;
  assign n36217 = n36215 & ~n36216;
  assign n36218 = P1_P2_INSTQUEUE_REG_3__6_ & ~n36208;
  assign n6346 = ~n36217 | n36218;
  assign n36220 = n35103 & n36187;
  assign n36221 = n35105 & n36190;
  assign n36222 = n35117 & n36195;
  assign n36223 = ~n36220 & ~n36221;
  assign n36224 = ~n36222 & n36223;
  assign n36225 = n35111 & n36200;
  assign n36226 = n36224 & ~n36225;
  assign n36227 = P1_P2_INSTQUEUE_REG_3__5_ & ~n36208;
  assign n6351 = ~n36226 | n36227;
  assign n36229 = n35125 & n36187;
  assign n36230 = n35127 & n36190;
  assign n36231 = n35139 & n36195;
  assign n36232 = ~n36229 & ~n36230;
  assign n36233 = ~n36231 & n36232;
  assign n36234 = n35133 & n36200;
  assign n36235 = n36233 & ~n36234;
  assign n36236 = P1_P2_INSTQUEUE_REG_3__4_ & ~n36208;
  assign n6356 = ~n36235 | n36236;
  assign n36238 = n35147 & n36187;
  assign n36239 = n35149 & n36190;
  assign n36240 = n35161 & n36195;
  assign n36241 = ~n36238 & ~n36239;
  assign n36242 = ~n36240 & n36241;
  assign n36243 = n35155 & n36200;
  assign n36244 = n36242 & ~n36243;
  assign n36245 = P1_P2_INSTQUEUE_REG_3__3_ & ~n36208;
  assign n6361 = ~n36244 | n36245;
  assign n36247 = n35169 & n36187;
  assign n36248 = n35171 & n36190;
  assign n36249 = n35183 & n36195;
  assign n36250 = ~n36247 & ~n36248;
  assign n36251 = ~n36249 & n36250;
  assign n36252 = n35177 & n36200;
  assign n36253 = n36251 & ~n36252;
  assign n36254 = P1_P2_INSTQUEUE_REG_3__2_ & ~n36208;
  assign n6366 = ~n36253 | n36254;
  assign n36256 = n35191 & n36187;
  assign n36257 = n35193 & n36190;
  assign n36258 = n35205 & n36195;
  assign n36259 = ~n36256 & ~n36257;
  assign n36260 = ~n36258 & n36259;
  assign n36261 = n35199 & n36200;
  assign n36262 = n36260 & ~n36261;
  assign n36263 = P1_P2_INSTQUEUE_REG_3__1_ & ~n36208;
  assign n6371 = ~n36262 | n36263;
  assign n36265 = n35213 & n36187;
  assign n36266 = n35215 & n36190;
  assign n36267 = n35227 & n36195;
  assign n36268 = ~n36265 & ~n36266;
  assign n36269 = ~n36267 & n36268;
  assign n36270 = n35221 & n36200;
  assign n36271 = n36269 & ~n36270;
  assign n36272 = P1_P2_INSTQUEUE_REG_3__0_ & ~n36208;
  assign n6376 = ~n36271 | n36272;
  assign n36274 = n35019 & n36186;
  assign n36275 = n35055 & n36274;
  assign n36276 = n35585 & n35927;
  assign n36277 = n35058 & n36276;
  assign n36278 = n35016 & n36192;
  assign n36279 = ~n36276 & ~n36278;
  assign n36280 = ~n36106 & ~n36279;
  assign n36281 = n35073 & n36280;
  assign n36282 = ~n36275 & ~n36277;
  assign n36283 = ~n36281 & n36282;
  assign n36284 = n35238 & n36199;
  assign n36285 = n35064 & n36284;
  assign n36286 = n36283 & ~n36285;
  assign n36287 = P1_P2_STATE2_REG_3_ & ~n36276;
  assign n36288 = n34998 & ~n36287;
  assign n36289 = ~n36274 & ~n36284;
  assign n36290 = n35015 & ~n36289;
  assign n36291 = n36279 & ~n36290;
  assign n36292 = n36288 & ~n36291;
  assign n36293 = P1_P2_INSTQUEUE_REG_2__7_ & ~n36292;
  assign n6381 = ~n36286 | n36293;
  assign n36295 = n35081 & n36274;
  assign n36296 = n35083 & n36276;
  assign n36297 = n35095 & n36280;
  assign n36298 = ~n36295 & ~n36296;
  assign n36299 = ~n36297 & n36298;
  assign n36300 = n35089 & n36284;
  assign n36301 = n36299 & ~n36300;
  assign n36302 = P1_P2_INSTQUEUE_REG_2__6_ & ~n36292;
  assign n6386 = ~n36301 | n36302;
  assign n36304 = n35103 & n36274;
  assign n36305 = n35105 & n36276;
  assign n36306 = n35117 & n36280;
  assign n36307 = ~n36304 & ~n36305;
  assign n36308 = ~n36306 & n36307;
  assign n36309 = n35111 & n36284;
  assign n36310 = n36308 & ~n36309;
  assign n36311 = P1_P2_INSTQUEUE_REG_2__5_ & ~n36292;
  assign n6391 = ~n36310 | n36311;
  assign n36313 = n35125 & n36274;
  assign n36314 = n35127 & n36276;
  assign n36315 = n35139 & n36280;
  assign n36316 = ~n36313 & ~n36314;
  assign n36317 = ~n36315 & n36316;
  assign n36318 = n35133 & n36284;
  assign n36319 = n36317 & ~n36318;
  assign n36320 = P1_P2_INSTQUEUE_REG_2__4_ & ~n36292;
  assign n6396 = ~n36319 | n36320;
  assign n36322 = n35147 & n36274;
  assign n36323 = n35149 & n36276;
  assign n36324 = n35161 & n36280;
  assign n36325 = ~n36322 & ~n36323;
  assign n36326 = ~n36324 & n36325;
  assign n36327 = n35155 & n36284;
  assign n36328 = n36326 & ~n36327;
  assign n36329 = P1_P2_INSTQUEUE_REG_2__3_ & ~n36292;
  assign n6401 = ~n36328 | n36329;
  assign n36331 = n35169 & n36274;
  assign n36332 = n35171 & n36276;
  assign n36333 = n35183 & n36280;
  assign n36334 = ~n36331 & ~n36332;
  assign n36335 = ~n36333 & n36334;
  assign n36336 = n35177 & n36284;
  assign n36337 = n36335 & ~n36336;
  assign n36338 = P1_P2_INSTQUEUE_REG_2__2_ & ~n36292;
  assign n6406 = ~n36337 | n36338;
  assign n36340 = n35191 & n36274;
  assign n36341 = n35193 & n36276;
  assign n36342 = n35205 & n36280;
  assign n36343 = ~n36340 & ~n36341;
  assign n36344 = ~n36342 & n36343;
  assign n36345 = n35199 & n36284;
  assign n36346 = n36344 & ~n36345;
  assign n36347 = P1_P2_INSTQUEUE_REG_2__1_ & ~n36292;
  assign n6411 = ~n36346 | n36347;
  assign n36349 = n35213 & n36274;
  assign n36350 = n35215 & n36276;
  assign n36351 = n35227 & n36280;
  assign n36352 = ~n36349 & ~n36350;
  assign n36353 = ~n36351 & n36352;
  assign n36354 = n35221 & n36284;
  assign n36355 = n36353 & ~n36354;
  assign n36356 = P1_P2_INSTQUEUE_REG_2__0_ & ~n36292;
  assign n6416 = ~n36355 | n36356;
  assign n36358 = n35020 & n36186;
  assign n36359 = n35055 & n36358;
  assign n36360 = n35007 & n36189;
  assign n36361 = n35058 & n36360;
  assign n36362 = n35017 & n36192;
  assign n36363 = ~n36360 & ~n36362;
  assign n36364 = ~n36106 & ~n36363;
  assign n36365 = n35073 & n36364;
  assign n36366 = ~n36359 & ~n36361;
  assign n36367 = ~n36365 & n36366;
  assign n36368 = n35326 & n36199;
  assign n36369 = n35064 & n36368;
  assign n36370 = n36367 & ~n36369;
  assign n36371 = P1_P2_STATE2_REG_3_ & ~n36360;
  assign n36372 = n34998 & ~n36371;
  assign n36373 = ~n36358 & ~n36368;
  assign n36374 = n35015 & ~n36373;
  assign n36375 = n36363 & ~n36374;
  assign n36376 = n36372 & ~n36375;
  assign n36377 = P1_P2_INSTQUEUE_REG_1__7_ & ~n36376;
  assign n6421 = ~n36370 | n36377;
  assign n36379 = n35081 & n36358;
  assign n36380 = n35083 & n36360;
  assign n36381 = n35095 & n36364;
  assign n36382 = ~n36379 & ~n36380;
  assign n36383 = ~n36381 & n36382;
  assign n36384 = n35089 & n36368;
  assign n36385 = n36383 & ~n36384;
  assign n36386 = P1_P2_INSTQUEUE_REG_1__6_ & ~n36376;
  assign n6426 = ~n36385 | n36386;
  assign n36388 = n35103 & n36358;
  assign n36389 = n35105 & n36360;
  assign n36390 = n35117 & n36364;
  assign n36391 = ~n36388 & ~n36389;
  assign n36392 = ~n36390 & n36391;
  assign n36393 = n35111 & n36368;
  assign n36394 = n36392 & ~n36393;
  assign n36395 = P1_P2_INSTQUEUE_REG_1__5_ & ~n36376;
  assign n6431 = ~n36394 | n36395;
  assign n36397 = n35125 & n36358;
  assign n36398 = n35127 & n36360;
  assign n36399 = n35139 & n36364;
  assign n36400 = ~n36397 & ~n36398;
  assign n36401 = ~n36399 & n36400;
  assign n36402 = n35133 & n36368;
  assign n36403 = n36401 & ~n36402;
  assign n36404 = P1_P2_INSTQUEUE_REG_1__4_ & ~n36376;
  assign n6436 = ~n36403 | n36404;
  assign n36406 = n35147 & n36358;
  assign n36407 = n35149 & n36360;
  assign n36408 = n35161 & n36364;
  assign n36409 = ~n36406 & ~n36407;
  assign n36410 = ~n36408 & n36409;
  assign n36411 = n35155 & n36368;
  assign n36412 = n36410 & ~n36411;
  assign n36413 = P1_P2_INSTQUEUE_REG_1__3_ & ~n36376;
  assign n6441 = ~n36412 | n36413;
  assign n36415 = n35169 & n36358;
  assign n36416 = n35171 & n36360;
  assign n36417 = n35183 & n36364;
  assign n36418 = ~n36415 & ~n36416;
  assign n36419 = ~n36417 & n36418;
  assign n36420 = n35177 & n36368;
  assign n36421 = n36419 & ~n36420;
  assign n36422 = P1_P2_INSTQUEUE_REG_1__2_ & ~n36376;
  assign n6446 = ~n36421 | n36422;
  assign n36424 = n35191 & n36358;
  assign n36425 = n35193 & n36360;
  assign n36426 = n35205 & n36364;
  assign n36427 = ~n36424 & ~n36425;
  assign n36428 = ~n36426 & n36427;
  assign n36429 = n35199 & n36368;
  assign n36430 = n36428 & ~n36429;
  assign n36431 = P1_P2_INSTQUEUE_REG_1__1_ & ~n36376;
  assign n6451 = ~n36430 | n36431;
  assign n36433 = n35213 & n36358;
  assign n36434 = n35215 & n36360;
  assign n36435 = n35227 & n36364;
  assign n36436 = ~n36433 & ~n36434;
  assign n36437 = ~n36435 & n36436;
  assign n36438 = n35221 & n36368;
  assign n36439 = n36437 & ~n36438;
  assign n36440 = P1_P2_INSTQUEUE_REG_1__0_ & ~n36376;
  assign n6456 = ~n36439 | n36440;
  assign n36442 = n35414 & n36186;
  assign n36443 = n35055 & n36442;
  assign n36444 = n35585 & n36103;
  assign n36445 = n35058 & n36444;
  assign n36446 = n35009 & n36192;
  assign n36447 = ~n36106 & n36446;
  assign n36448 = n35073 & n36447;
  assign n36449 = ~n36443 & ~n36445;
  assign n36450 = ~n36448 & n36449;
  assign n36451 = n35412 & n36199;
  assign n36452 = n35064 & n36451;
  assign n36453 = n36450 & ~n36452;
  assign n36454 = P1_P2_STATE2_REG_3_ & ~n36444;
  assign n36455 = n34998 & ~n36454;
  assign n36456 = ~n36442 & ~n36451;
  assign n36457 = n35015 & ~n36456;
  assign n36458 = ~n36446 & ~n36457;
  assign n36459 = n36455 & ~n36458;
  assign n36460 = P1_P2_INSTQUEUE_REG_0__7_ & ~n36459;
  assign n6461 = ~n36453 | n36460;
  assign n36462 = n35081 & n36442;
  assign n36463 = n35083 & n36444;
  assign n36464 = n35095 & n36447;
  assign n36465 = ~n36462 & ~n36463;
  assign n36466 = ~n36464 & n36465;
  assign n36467 = n35089 & n36451;
  assign n36468 = n36466 & ~n36467;
  assign n36469 = P1_P2_INSTQUEUE_REG_0__6_ & ~n36459;
  assign n6466 = ~n36468 | n36469;
  assign n36471 = n35103 & n36442;
  assign n36472 = n35105 & n36444;
  assign n36473 = n35117 & n36447;
  assign n36474 = ~n36471 & ~n36472;
  assign n36475 = ~n36473 & n36474;
  assign n36476 = n35111 & n36451;
  assign n36477 = n36475 & ~n36476;
  assign n36478 = P1_P2_INSTQUEUE_REG_0__5_ & ~n36459;
  assign n6471 = ~n36477 | n36478;
  assign n36480 = n35125 & n36442;
  assign n36481 = n35127 & n36444;
  assign n36482 = n35139 & n36447;
  assign n36483 = ~n36480 & ~n36481;
  assign n36484 = ~n36482 & n36483;
  assign n36485 = n35133 & n36451;
  assign n36486 = n36484 & ~n36485;
  assign n36487 = P1_P2_INSTQUEUE_REG_0__4_ & ~n36459;
  assign n6476 = ~n36486 | n36487;
  assign n36489 = n35147 & n36442;
  assign n36490 = n35149 & n36444;
  assign n36491 = n35161 & n36447;
  assign n36492 = ~n36489 & ~n36490;
  assign n36493 = ~n36491 & n36492;
  assign n36494 = n35155 & n36451;
  assign n36495 = n36493 & ~n36494;
  assign n36496 = P1_P2_INSTQUEUE_REG_0__3_ & ~n36459;
  assign n6481 = ~n36495 | n36496;
  assign n36498 = n35169 & n36442;
  assign n36499 = n35171 & n36444;
  assign n36500 = n35183 & n36447;
  assign n36501 = ~n36498 & ~n36499;
  assign n36502 = ~n36500 & n36501;
  assign n36503 = n35177 & n36451;
  assign n36504 = n36502 & ~n36503;
  assign n36505 = P1_P2_INSTQUEUE_REG_0__2_ & ~n36459;
  assign n6486 = ~n36504 | n36505;
  assign n36507 = n35191 & n36442;
  assign n36508 = n35193 & n36444;
  assign n36509 = n35205 & n36447;
  assign n36510 = ~n36507 & ~n36508;
  assign n36511 = ~n36509 & n36510;
  assign n36512 = n35199 & n36451;
  assign n36513 = n36511 & ~n36512;
  assign n36514 = P1_P2_INSTQUEUE_REG_0__1_ & ~n36459;
  assign n6491 = ~n36513 | n36514;
  assign n36516 = n35213 & n36442;
  assign n36517 = n35215 & n36444;
  assign n36518 = n35227 & n36447;
  assign n36519 = ~n36516 & ~n36517;
  assign n36520 = ~n36518 & n36519;
  assign n36521 = n35221 & n36451;
  assign n36522 = n36520 & ~n36521;
  assign n36523 = P1_P2_INSTQUEUE_REG_0__0_ & ~n36459;
  assign n6496 = ~n36522 | n36523;
  assign n36525 = P1_P2_STATE2_REG_3_ & ~P1_P2_STATE2_REG_0_;
  assign n36526 = P1_P2_STATE2_REG_0_ & P1_P2_FLUSH_REG;
  assign n36527 = n34293 & n36526;
  assign n36528 = ~n36525 & ~n36527;
  assign n36529 = ~n34825 & n34935;
  assign n36530 = n36528 & ~n36529;
  assign n36531 = P1_P2_INSTQUEUERD_ADDR_REG_4_ & n36530;
  assign n36532 = ~n34868 & n34941;
  assign n36533 = n34660 & n36532;
  assign n36534 = ~n36530 & n36533;
  assign n6501 = n36531 | n36534;
  assign n36536 = ~n34859 & n34941;
  assign n36537 = ~n34332 & ~n34832;
  assign n36538 = n34950 & ~n36537;
  assign n36539 = ~n36536 & ~n36538;
  assign n36540 = ~n36530 & ~n36539;
  assign n36541 = P1_P2_INSTQUEUERD_ADDR_REG_3_ & n36530;
  assign n6506 = n36540 | n36541;
  assign n36543 = ~n34783 & n34950;
  assign n36544 = P1_P2_STATE2_REG_1_ & ~n34957;
  assign n36545 = ~n34966 & n36544;
  assign n36546 = ~n36543 & ~n36545;
  assign n36547 = ~n34799 & n34941;
  assign n36548 = n36546 & ~n36547;
  assign n36549 = ~n36530 & ~n36548;
  assign n36550 = P1_P2_INSTQUEUERD_ADDR_REG_2_ & n36530;
  assign n6511 = n36549 | n36550;
  assign n36552 = n34895 & n34950;
  assign n36553 = n34966 & n36544;
  assign n36554 = ~n36552 & ~n36553;
  assign n36555 = ~n34900 & n34941;
  assign n36556 = n36554 & ~n36555;
  assign n36557 = ~n36530 & ~n36556;
  assign n36558 = P1_P2_INSTQUEUERD_ADDR_REG_1_ & n36530;
  assign n6516 = n36557 | n36558;
  assign n36560 = P1_P2_STATE2_REG_1_ & n34957;
  assign n36561 = ~P1_P2_INSTQUEUERD_ADDR_REG_0_ & n34950;
  assign n36562 = ~n36560 & ~n36561;
  assign n36563 = ~n34886 & n34941;
  assign n36564 = n36562 & ~n36563;
  assign n36565 = ~n36530 & ~n36564;
  assign n36566 = P1_P2_INSTQUEUERD_ADDR_REG_0_ & n36530;
  assign n6521 = n36565 | n36566;
  assign n36568 = P1_P2_STATE2_REG_0_ & n34293;
  assign n36569 = ~n34980 & n36568;
  assign n36570 = ~n34998 & ~n36527;
  assign n36571 = ~n36569 & n36570;
  assign n6526 = P1_P2_INSTQUEUEWR_ADDR_REG_4_ & n36571;
  assign n36573 = P1_P2_STATE2_REG_3_ & ~n34992;
  assign n36574 = ~n36571 & ~n36573;
  assign n36575 = P1_P2_INSTQUEUEWR_ADDR_REG_3_ & ~n36574;
  assign n36576 = ~n34941 & ~n35014;
  assign n36577 = ~n35034 & ~n36576;
  assign n36578 = P1_P2_STATE2_REG_3_ & n35003;
  assign n36579 = ~n36577 & ~n36578;
  assign n36580 = n35022 & ~n35029;
  assign n36581 = ~n35040 & ~n36580;
  assign n36582 = ~n35847 & ~n36581;
  assign n36583 = n35053 & ~n36582;
  assign n36584 = n36579 & ~n36583;
  assign n36585 = ~n36571 & ~n36584;
  assign n6531 = n36575 | n36585;
  assign n36587 = ~n35025 & ~n36576;
  assign n36588 = P1_P2_STATE2_REG_3_ & ~P1_P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n36589 = n34991 & n36588;
  assign n36590 = ~n36587 & ~n36589;
  assign n36591 = ~n35022 & ~n35029;
  assign n36592 = n35022 & n35029;
  assign n36593 = ~n36591 & ~n36592;
  assign n36594 = n35053 & ~n36593;
  assign n36595 = n36590 & ~n36594;
  assign n36596 = ~n36571 & ~n36595;
  assign n36597 = P1_P2_STATE2_REG_3_ & ~n34991;
  assign n36598 = ~n36571 & ~n36597;
  assign n36599 = P1_P2_INSTQUEUEWR_ADDR_REG_2_ & ~n36598;
  assign n6536 = n36596 | n36599;
  assign n36601 = ~n35018 & ~n36576;
  assign n36602 = P1_P2_STATE2_REG_3_ & ~P1_P2_INSTQUEUEWR_ADDR_REG_1_;
  assign n36603 = ~n35021 & n35053;
  assign n36604 = ~n36602 & ~n36603;
  assign n36605 = P1_P2_INSTQUEUEWR_ADDR_REG_0_ & ~n36604;
  assign n36606 = n35053 & n35326;
  assign n36607 = ~n36601 & ~n36605;
  assign n36608 = ~n36606 & n36607;
  assign n36609 = ~n36571 & ~n36608;
  assign n36610 = P1_P2_STATE2_REG_3_ & ~P1_P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n36611 = ~n36571 & ~n36610;
  assign n36612 = P1_P2_INSTQUEUEWR_ADDR_REG_1_ & ~n36611;
  assign n6541 = n36609 | n36612;
  assign n36614 = ~n34941 & ~n35013;
  assign n36615 = ~n36571 & n36614;
  assign n36616 = P1_P2_INSTQUEUEWR_ADDR_REG_0_ & ~n36615;
  assign n36617 = ~n34981 & ~n36610;
  assign n36618 = ~n36571 & ~n36617;
  assign n6546 = n36616 | n36618;
  assign n36620 = ~P1_P2_STATE2_REG_1_ & n35013;
  assign n36621 = ~P1_P2_STATE2_REG_0_ & n36620;
  assign n36622 = n34589 & n34633;
  assign n36623 = ~n34421 & ~n34580;
  assign n36624 = n34678 & n36623;
  assign n36625 = n34587 & n34633;
  assign n36626 = ~n34817 & ~n36624;
  assign n36627 = ~n36625 & n36626;
  assign n36628 = n34638 & n34686;
  assign n36629 = n34390 & n34585;
  assign n36630 = n34633 & n36629;
  assign n36631 = ~n36628 & ~n36630;
  assign n36632 = n34549 & ~n36631;
  assign n36633 = ~n34389 & n34692;
  assign n36634 = ~n34208 & n34358;
  assign n36635 = n34633 & n36634;
  assign n36636 = ~n36633 & ~n36635;
  assign n36637 = ~n34549 & ~n36636;
  assign n36638 = n34580 & n34678;
  assign n36639 = ~n36632 & ~n36637;
  assign n36640 = ~n36638 & n36639;
  assign n36641 = n34514 & ~n36640;
  assign n36642 = n34809 & ~n36622;
  assign n36643 = n36627 & n36642;
  assign n36644 = ~n36641 & n36643;
  assign n36645 = n34935 & ~n36644;
  assign n36646 = ~n36621 & ~n36645;
  assign n36647 = P1_P2_STATE2_REG_2_ & ~n36646;
  assign n36648 = ~P1_P2_INSTADDRPOINTER_REG_0_ & n34879;
  assign n36649 = ~P1_P2_INSTADDRPOINTER_REG_0_ & n34722;
  assign n36650 = ~n36648 & ~n36649;
  assign n36651 = ~P1_P2_INSTADDRPOINTER_REG_0_ & ~n34769;
  assign n36652 = P1_P2_INSTADDRPOINTER_REG_0_ & n34840;
  assign n36653 = P1_P2_INSTADDRPOINTER_REG_0_ & n34841;
  assign n36654 = n34581 & n34712;
  assign n36655 = n34718 & n36654;
  assign n36656 = ~P1_P2_INSTADDRPOINTER_REG_0_ & n36655;
  assign n36657 = n34658 & n34712;
  assign n36658 = n34718 & n36657;
  assign n36659 = ~P1_P2_INSTADDRPOINTER_REG_0_ & n36658;
  assign n36660 = ~n36656 & ~n36659;
  assign n36661 = P1_P2_INSTADDRPOINTER_REG_0_ & n34656;
  assign n36662 = n36660 & ~n36661;
  assign n36663 = n34783 & n36537;
  assign n36664 = P1_P2_INSTQUEUERD_ADDR_REG_0_ & ~n34895;
  assign n36665 = n36663 & n36664;
  assign n36666 = P1_P2_INSTQUEUE_REG_0__0_ & n36665;
  assign n36667 = ~P1_P2_INSTQUEUERD_ADDR_REG_0_ & ~n34895;
  assign n36668 = n36663 & n36667;
  assign n36669 = P1_P2_INSTQUEUE_REG_1__0_ & n36668;
  assign n36670 = P1_P2_INSTQUEUERD_ADDR_REG_0_ & n34895;
  assign n36671 = n36663 & n36670;
  assign n36672 = P1_P2_INSTQUEUE_REG_2__0_ & n36671;
  assign n36673 = ~P1_P2_INSTQUEUERD_ADDR_REG_0_ & n34895;
  assign n36674 = n36663 & n36673;
  assign n36675 = P1_P2_INSTQUEUE_REG_3__0_ & n36674;
  assign n36676 = ~n36666 & ~n36669;
  assign n36677 = ~n36672 & n36676;
  assign n36678 = ~n36675 & n36677;
  assign n36679 = ~n34783 & n36537;
  assign n36680 = n36664 & n36679;
  assign n36681 = P1_P2_INSTQUEUE_REG_4__0_ & n36680;
  assign n36682 = n36667 & n36679;
  assign n36683 = P1_P2_INSTQUEUE_REG_5__0_ & n36682;
  assign n36684 = n36670 & n36679;
  assign n36685 = P1_P2_INSTQUEUE_REG_6__0_ & n36684;
  assign n36686 = n36673 & n36679;
  assign n36687 = P1_P2_INSTQUEUE_REG_7__0_ & n36686;
  assign n36688 = ~n36681 & ~n36683;
  assign n36689 = ~n36685 & n36688;
  assign n36690 = ~n36687 & n36689;
  assign n36691 = n34783 & ~n36537;
  assign n36692 = n36664 & n36691;
  assign n36693 = P1_P2_INSTQUEUE_REG_8__0_ & n36692;
  assign n36694 = n36667 & n36691;
  assign n36695 = P1_P2_INSTQUEUE_REG_9__0_ & n36694;
  assign n36696 = n36670 & n36691;
  assign n36697 = P1_P2_INSTQUEUE_REG_10__0_ & n36696;
  assign n36698 = n36673 & n36691;
  assign n36699 = P1_P2_INSTQUEUE_REG_11__0_ & n36698;
  assign n36700 = ~n36693 & ~n36695;
  assign n36701 = ~n36697 & n36700;
  assign n36702 = ~n36699 & n36701;
  assign n36703 = ~n34783 & ~n36537;
  assign n36704 = n36664 & n36703;
  assign n36705 = P1_P2_INSTQUEUE_REG_12__0_ & n36704;
  assign n36706 = n36667 & n36703;
  assign n36707 = P1_P2_INSTQUEUE_REG_13__0_ & n36706;
  assign n36708 = n36670 & n36703;
  assign n36709 = P1_P2_INSTQUEUE_REG_14__0_ & n36708;
  assign n36710 = n36673 & n36703;
  assign n36711 = P1_P2_INSTQUEUE_REG_15__0_ & n36710;
  assign n36712 = ~n36705 & ~n36707;
  assign n36713 = ~n36709 & n36712;
  assign n36714 = ~n36711 & n36713;
  assign n36715 = n36678 & n36690;
  assign n36716 = n36702 & n36715;
  assign n36717 = n36714 & n36716;
  assign n36718 = P1_P2_INSTADDRPOINTER_REG_0_ & n36717;
  assign n36719 = ~P1_P2_INSTADDRPOINTER_REG_0_ & ~n36717;
  assign n36720 = ~n36718 & ~n36719;
  assign n36721 = P1_P2_INSTQUEUE_REG_0__7_ & n36665;
  assign n36722 = P1_P2_INSTQUEUE_REG_1__7_ & n36668;
  assign n36723 = P1_P2_INSTQUEUE_REG_2__7_ & n36671;
  assign n36724 = P1_P2_INSTQUEUE_REG_3__7_ & n36674;
  assign n36725 = ~n36721 & ~n36722;
  assign n36726 = ~n36723 & n36725;
  assign n36727 = ~n36724 & n36726;
  assign n36728 = P1_P2_INSTQUEUE_REG_4__7_ & n36680;
  assign n36729 = P1_P2_INSTQUEUE_REG_5__7_ & n36682;
  assign n36730 = P1_P2_INSTQUEUE_REG_6__7_ & n36684;
  assign n36731 = P1_P2_INSTQUEUE_REG_7__7_ & n36686;
  assign n36732 = ~n36728 & ~n36729;
  assign n36733 = ~n36730 & n36732;
  assign n36734 = ~n36731 & n36733;
  assign n36735 = P1_P2_INSTQUEUE_REG_8__7_ & n36692;
  assign n36736 = P1_P2_INSTQUEUE_REG_9__7_ & n36694;
  assign n36737 = P1_P2_INSTQUEUE_REG_10__7_ & n36696;
  assign n36738 = P1_P2_INSTQUEUE_REG_11__7_ & n36698;
  assign n36739 = ~n36735 & ~n36736;
  assign n36740 = ~n36737 & n36739;
  assign n36741 = ~n36738 & n36740;
  assign n36742 = P1_P2_INSTQUEUE_REG_12__7_ & n36704;
  assign n36743 = P1_P2_INSTQUEUE_REG_13__7_ & n36706;
  assign n36744 = P1_P2_INSTQUEUE_REG_14__7_ & n36708;
  assign n36745 = P1_P2_INSTQUEUE_REG_15__7_ & n36710;
  assign n36746 = ~n36742 & ~n36743;
  assign n36747 = ~n36744 & n36746;
  assign n36748 = ~n36745 & n36747;
  assign n36749 = n36727 & n36734;
  assign n36750 = n36741 & n36749;
  assign n36751 = n36748 & n36750;
  assign n36752 = n34688 & ~n36751;
  assign n36753 = ~n36720 & n36752;
  assign n36754 = n34688 & n36751;
  assign n36755 = ~n36720 & n36754;
  assign n36756 = ~n36652 & ~n36653;
  assign n36757 = n36662 & n36756;
  assign n36758 = ~n36753 & n36757;
  assign n36759 = ~n36755 & n36758;
  assign n36760 = n34654 & n34682;
  assign n36761 = ~P1_P2_INSTADDRPOINTER_REG_0_ & n36760;
  assign n36762 = ~P1_P2_INSTADDRPOINTER_REG_0_ & n34726;
  assign n36763 = n34483 & n34669;
  assign n36764 = n34715 & n36763;
  assign n36765 = ~P1_P2_INSTADDRPOINTER_REG_0_ & n36764;
  assign n36766 = ~P1_P2_INSTADDRPOINTER_REG_0_ & n36717;
  assign n36767 = P1_P2_INSTADDRPOINTER_REG_0_ & ~n36717;
  assign n36768 = ~n36766 & ~n36767;
  assign n36769 = n34683 & ~n36768;
  assign n36770 = n34358 & n34712;
  assign n36771 = n34715 & n36770;
  assign n36772 = ~P1_P2_INSTADDRPOINTER_REG_0_ & n36771;
  assign n36773 = ~n36761 & ~n36762;
  assign n36774 = ~n36765 & n36773;
  assign n36775 = ~n36769 & n36774;
  assign n36776 = ~n36772 & n36775;
  assign n36777 = P1_P2_INSTADDRPOINTER_REG_0_ & n34582;
  assign n36778 = P1_P2_INSTADDRPOINTER_REG_0_ & n34660;
  assign n36779 = P1_P2_INSTADDRPOINTER_REG_0_ & n34664;
  assign n36780 = ~P1_P2_INSTADDRPOINTER_REG_0_ & n34680;
  assign n36781 = ~P1_P2_INSTADDRPOINTER_REG_0_ & n34672;
  assign n36782 = ~n36777 & ~n36778;
  assign n36783 = ~n36779 & n36782;
  assign n36784 = ~n36780 & n36783;
  assign n36785 = ~n36781 & n36784;
  assign n36786 = n36776 & n36785;
  assign n36787 = n36650 & ~n36651;
  assign n36788 = n36759 & n36787;
  assign n36789 = n36786 & n36788;
  assign n36790 = n36647 & ~n36789;
  assign n36791 = ~P1_P2_STATE2_REG_2_ & ~n36646;
  assign n36792 = P1_P2_REIP_REG_0_ & n36791;
  assign n36793 = P1_P2_INSTADDRPOINTER_REG_0_ & n36646;
  assign n36794 = ~n36790 & ~n36792;
  assign n6551 = n36793 | ~n36794;
  assign n36796 = P1_P2_INSTADDRPOINTER_REG_1_ & n36646;
  assign n36797 = P1_P2_REIP_REG_1_ & n36791;
  assign n36798 = ~n34769 & ~n34963;
  assign n36799 = n34879 & ~n34963;
  assign n36800 = n34722 & ~n34963;
  assign n36801 = ~n36799 & ~n36800;
  assign n36802 = ~P1_P2_INSTADDRPOINTER_REG_1_ & n36767;
  assign n36803 = P1_P2_INSTADDRPOINTER_REG_1_ & ~n36767;
  assign n36804 = ~n36802 & ~n36803;
  assign n36805 = P1_P2_INSTQUEUE_REG_0__1_ & n36665;
  assign n36806 = P1_P2_INSTQUEUE_REG_1__1_ & n36668;
  assign n36807 = P1_P2_INSTQUEUE_REG_2__1_ & n36671;
  assign n36808 = P1_P2_INSTQUEUE_REG_3__1_ & n36674;
  assign n36809 = ~n36805 & ~n36806;
  assign n36810 = ~n36807 & n36809;
  assign n36811 = ~n36808 & n36810;
  assign n36812 = P1_P2_INSTQUEUE_REG_4__1_ & n36680;
  assign n36813 = P1_P2_INSTQUEUE_REG_5__1_ & n36682;
  assign n36814 = P1_P2_INSTQUEUE_REG_6__1_ & n36684;
  assign n36815 = P1_P2_INSTQUEUE_REG_7__1_ & n36686;
  assign n36816 = ~n36812 & ~n36813;
  assign n36817 = ~n36814 & n36816;
  assign n36818 = ~n36815 & n36817;
  assign n36819 = P1_P2_INSTQUEUE_REG_8__1_ & n36692;
  assign n36820 = P1_P2_INSTQUEUE_REG_9__1_ & n36694;
  assign n36821 = P1_P2_INSTQUEUE_REG_10__1_ & n36696;
  assign n36822 = P1_P2_INSTQUEUE_REG_11__1_ & n36698;
  assign n36823 = ~n36819 & ~n36820;
  assign n36824 = ~n36821 & n36823;
  assign n36825 = ~n36822 & n36824;
  assign n36826 = P1_P2_INSTQUEUE_REG_12__1_ & n36704;
  assign n36827 = P1_P2_INSTQUEUE_REG_13__1_ & n36706;
  assign n36828 = P1_P2_INSTQUEUE_REG_14__1_ & n36708;
  assign n36829 = P1_P2_INSTQUEUE_REG_15__1_ & n36710;
  assign n36830 = ~n36826 & ~n36827;
  assign n36831 = ~n36828 & n36830;
  assign n36832 = ~n36829 & n36831;
  assign n36833 = n36811 & n36818;
  assign n36834 = n36825 & n36833;
  assign n36835 = n36832 & n36834;
  assign n36836 = ~n36804 & ~n36835;
  assign n36837 = ~P1_P2_INSTADDRPOINTER_REG_1_ & ~n36767;
  assign n36838 = n36835 & n36837;
  assign n36839 = n36767 & n36835;
  assign n36840 = P1_P2_INSTADDRPOINTER_REG_1_ & n36839;
  assign n36841 = ~n36836 & ~n36838;
  assign n36842 = ~n36840 & n36841;
  assign n36843 = n36754 & ~n36842;
  assign n36844 = ~n34963 & n36771;
  assign n36845 = ~n34963 & n36764;
  assign n36846 = ~n34963 & n36760;
  assign n36847 = n34726 & ~n34963;
  assign n36848 = ~n36844 & ~n36845;
  assign n36849 = ~n36846 & n36848;
  assign n36850 = ~n36847 & n36849;
  assign n36851 = ~P1_P2_INSTADDRPOINTER_REG_1_ & n34582;
  assign n36852 = ~P1_P2_INSTADDRPOINTER_REG_1_ & n34660;
  assign n36853 = ~P1_P2_INSTADDRPOINTER_REG_1_ & n34664;
  assign n36854 = n34680 & ~n34963;
  assign n36855 = n34672 & ~n34963;
  assign n36856 = ~n36851 & ~n36852;
  assign n36857 = ~n36853 & n36856;
  assign n36858 = ~n36854 & n36857;
  assign n36859 = ~n36855 & n36858;
  assign n36860 = ~P1_P2_INSTADDRPOINTER_REG_1_ & n36718;
  assign n36861 = P1_P2_INSTADDRPOINTER_REG_1_ & ~n36718;
  assign n36862 = ~n36860 & ~n36861;
  assign n36863 = ~n36717 & n36835;
  assign n36864 = n36717 & ~n36835;
  assign n36865 = ~n36863 & ~n36864;
  assign n36866 = ~n36862 & n36865;
  assign n36867 = ~P1_P2_INSTADDRPOINTER_REG_1_ & ~n36718;
  assign n36868 = ~n36865 & n36867;
  assign n36869 = n36718 & ~n36865;
  assign n36870 = P1_P2_INSTADDRPOINTER_REG_1_ & n36869;
  assign n36871 = ~n36866 & ~n36868;
  assign n36872 = ~n36870 & n36871;
  assign n36873 = n34683 & ~n36872;
  assign n36874 = n36850 & n36859;
  assign n36875 = ~n36873 & n36874;
  assign n36876 = ~P1_P2_INSTADDRPOINTER_REG_1_ & n34840;
  assign n36877 = ~P1_P2_INSTADDRPOINTER_REG_1_ & n34841;
  assign n36878 = ~n34963 & n36655;
  assign n36879 = ~n34963 & n36658;
  assign n36880 = ~n36878 & ~n36879;
  assign n36881 = ~P1_P2_INSTADDRPOINTER_REG_1_ & n34656;
  assign n36882 = n36880 & ~n36881;
  assign n36883 = n36767 & ~n36835;
  assign n36884 = ~n36767 & n36835;
  assign n36885 = ~n36883 & ~n36884;
  assign n36886 = ~P1_P2_INSTADDRPOINTER_REG_1_ & ~n36885;
  assign n36887 = ~n36767 & ~n36835;
  assign n36888 = P1_P2_INSTADDRPOINTER_REG_1_ & n36887;
  assign n36889 = P1_P2_INSTADDRPOINTER_REG_1_ & n36767;
  assign n36890 = n36835 & n36889;
  assign n36891 = ~n36886 & ~n36888;
  assign n36892 = ~n36890 & n36891;
  assign n36893 = n36752 & ~n36892;
  assign n36894 = ~n36876 & ~n36877;
  assign n36895 = n36882 & n36894;
  assign n36896 = ~n36893 & n36895;
  assign n36897 = ~n36798 & n36801;
  assign n36898 = ~n36843 & n36897;
  assign n36899 = n36875 & n36898;
  assign n36900 = n36896 & n36899;
  assign n36901 = n36647 & ~n36900;
  assign n36902 = ~n36796 & ~n36797;
  assign n6556 = n36901 | ~n36902;
  assign n36904 = P1_P2_INSTADDRPOINTER_REG_2_ & n36646;
  assign n36905 = P1_P2_REIP_REG_2_ & n36791;
  assign n36906 = P1_P2_INSTADDRPOINTER_REG_0_ & P1_P2_INSTADDRPOINTER_REG_1_;
  assign n36907 = ~P1_P2_INSTADDRPOINTER_REG_2_ & n36906;
  assign n36908 = P1_P2_INSTADDRPOINTER_REG_2_ & ~n36906;
  assign n36909 = ~n36907 & ~n36908;
  assign n36910 = ~n34769 & ~n36909;
  assign n36911 = P1_P2_INSTADDRPOINTER_REG_1_ & ~P1_P2_INSTADDRPOINTER_REG_2_;
  assign n36912 = ~P1_P2_INSTADDRPOINTER_REG_1_ & P1_P2_INSTADDRPOINTER_REG_2_;
  assign n36913 = ~n36911 & ~n36912;
  assign n36914 = n34840 & ~n36913;
  assign n36915 = n34841 & ~n36913;
  assign n36916 = n36655 & ~n36909;
  assign n36917 = n36658 & ~n36909;
  assign n36918 = ~n36916 & ~n36917;
  assign n36919 = n34656 & ~n36913;
  assign n36920 = n36918 & ~n36919;
  assign n36921 = ~n36914 & ~n36915;
  assign n36922 = n36920 & n36921;
  assign n36923 = P1_P2_INSTADDRPOINTER_REG_1_ & ~n36887;
  assign n36924 = ~n36839 & ~n36923;
  assign n36925 = P1_P2_INSTQUEUE_REG_0__2_ & n36665;
  assign n36926 = P1_P2_INSTQUEUE_REG_1__2_ & n36668;
  assign n36927 = P1_P2_INSTQUEUE_REG_2__2_ & n36671;
  assign n36928 = P1_P2_INSTQUEUE_REG_3__2_ & n36674;
  assign n36929 = ~n36925 & ~n36926;
  assign n36930 = ~n36927 & n36929;
  assign n36931 = ~n36928 & n36930;
  assign n36932 = P1_P2_INSTQUEUE_REG_4__2_ & n36680;
  assign n36933 = P1_P2_INSTQUEUE_REG_5__2_ & n36682;
  assign n36934 = P1_P2_INSTQUEUE_REG_6__2_ & n36684;
  assign n36935 = P1_P2_INSTQUEUE_REG_7__2_ & n36686;
  assign n36936 = ~n36932 & ~n36933;
  assign n36937 = ~n36934 & n36936;
  assign n36938 = ~n36935 & n36937;
  assign n36939 = P1_P2_INSTQUEUE_REG_8__2_ & n36692;
  assign n36940 = P1_P2_INSTQUEUE_REG_9__2_ & n36694;
  assign n36941 = P1_P2_INSTQUEUE_REG_10__2_ & n36696;
  assign n36942 = P1_P2_INSTQUEUE_REG_11__2_ & n36698;
  assign n36943 = ~n36939 & ~n36940;
  assign n36944 = ~n36941 & n36943;
  assign n36945 = ~n36942 & n36944;
  assign n36946 = P1_P2_INSTQUEUE_REG_12__2_ & n36704;
  assign n36947 = P1_P2_INSTQUEUE_REG_13__2_ & n36706;
  assign n36948 = P1_P2_INSTQUEUE_REG_14__2_ & n36708;
  assign n36949 = P1_P2_INSTQUEUE_REG_15__2_ & n36710;
  assign n36950 = ~n36946 & ~n36947;
  assign n36951 = ~n36948 & n36950;
  assign n36952 = ~n36949 & n36951;
  assign n36953 = n36931 & n36938;
  assign n36954 = n36945 & n36953;
  assign n36955 = n36952 & n36954;
  assign n36956 = ~n36835 & n36955;
  assign n36957 = n36835 & ~n36955;
  assign n36958 = ~n36956 & ~n36957;
  assign n36959 = ~P1_P2_INSTADDRPOINTER_REG_2_ & ~n36958;
  assign n36960 = P1_P2_INSTADDRPOINTER_REG_2_ & n36958;
  assign n36961 = ~n36959 & ~n36960;
  assign n36962 = n36924 & ~n36961;
  assign n36963 = ~n36924 & n36961;
  assign n36964 = ~n36962 & ~n36963;
  assign n36965 = n36754 & ~n36964;
  assign n36966 = n34879 & ~n36909;
  assign n36967 = n34722 & ~n36909;
  assign n36968 = ~n36966 & ~n36967;
  assign n36969 = P1_P2_INSTADDRPOINTER_REG_1_ & n36835;
  assign n36970 = ~n36839 & ~n36889;
  assign n36971 = ~n36969 & n36970;
  assign n36972 = ~n36961 & n36971;
  assign n36973 = ~P1_P2_INSTADDRPOINTER_REG_2_ & n36958;
  assign n36974 = P1_P2_INSTADDRPOINTER_REG_2_ & ~n36958;
  assign n36975 = ~n36973 & ~n36974;
  assign n36976 = ~n36971 & ~n36975;
  assign n36977 = ~n36972 & ~n36976;
  assign n36978 = n36752 & ~n36977;
  assign n36979 = n36968 & ~n36978;
  assign n36980 = n36771 & ~n36909;
  assign n36981 = n36764 & ~n36909;
  assign n36982 = n36760 & ~n36909;
  assign n36983 = n34726 & ~n36909;
  assign n36984 = ~n36980 & ~n36981;
  assign n36985 = ~n36982 & n36984;
  assign n36986 = ~n36983 & n36985;
  assign n36987 = n34582 & ~n36913;
  assign n36988 = n34660 & ~n36913;
  assign n36989 = n34664 & ~n36913;
  assign n36990 = ~P1_P2_INSTADDRPOINTER_REG_2_ & ~n36906;
  assign n36991 = P1_P2_INSTADDRPOINTER_REG_2_ & n36906;
  assign n36992 = ~n36990 & ~n36991;
  assign n36993 = n34680 & ~n36992;
  assign n36994 = n34672 & ~n36992;
  assign n36995 = ~n36987 & ~n36988;
  assign n36996 = ~n36989 & n36995;
  assign n36997 = ~n36993 & n36996;
  assign n36998 = ~n36994 & n36997;
  assign n36999 = ~n36717 & ~n36835;
  assign n37000 = n36955 & ~n36999;
  assign n37001 = ~n36955 & n36999;
  assign n37002 = ~n37000 & ~n37001;
  assign n37003 = ~P1_P2_INSTADDRPOINTER_REG_2_ & ~n37002;
  assign n37004 = P1_P2_INSTADDRPOINTER_REG_2_ & n37002;
  assign n37005 = ~n37003 & ~n37004;
  assign n37006 = ~n36718 & n36865;
  assign n37007 = P1_P2_INSTADDRPOINTER_REG_1_ & ~n37006;
  assign n37008 = ~n36869 & ~n37007;
  assign n37009 = ~n37005 & n37008;
  assign n37010 = ~P1_P2_INSTADDRPOINTER_REG_2_ & n37002;
  assign n37011 = P1_P2_INSTADDRPOINTER_REG_2_ & ~n37002;
  assign n37012 = ~n37010 & ~n37011;
  assign n37013 = ~n37008 & ~n37012;
  assign n37014 = ~n37009 & ~n37013;
  assign n37015 = n34683 & ~n37014;
  assign n37016 = n36986 & n36998;
  assign n37017 = ~n37015 & n37016;
  assign n37018 = ~n36910 & n36922;
  assign n37019 = ~n36965 & n37018;
  assign n37020 = n36979 & n37019;
  assign n37021 = n37017 & n37020;
  assign n37022 = n36647 & ~n37021;
  assign n37023 = ~n36904 & ~n36905;
  assign n6561 = n37022 | ~n37023;
  assign n37025 = P1_P2_INSTADDRPOINTER_REG_3_ & n36646;
  assign n37026 = P1_P2_REIP_REG_3_ & n36791;
  assign n37027 = ~P1_P2_INSTADDRPOINTER_REG_3_ & n36991;
  assign n37028 = P1_P2_INSTADDRPOINTER_REG_3_ & ~n36991;
  assign n37029 = ~n37027 & ~n37028;
  assign n37030 = n34879 & ~n37029;
  assign n37031 = n34722 & ~n37029;
  assign n37032 = ~n37030 & ~n37031;
  assign n37033 = ~n34769 & ~n37029;
  assign n37034 = P1_P2_INSTADDRPOINTER_REG_1_ & P1_P2_INSTADDRPOINTER_REG_2_;
  assign n37035 = ~P1_P2_INSTADDRPOINTER_REG_3_ & n37034;
  assign n37036 = P1_P2_INSTADDRPOINTER_REG_3_ & ~n37034;
  assign n37037 = ~n37035 & ~n37036;
  assign n37038 = n34840 & ~n37037;
  assign n37039 = n34841 & ~n37037;
  assign n37040 = n36655 & ~n37029;
  assign n37041 = n36658 & ~n37029;
  assign n37042 = ~n37040 & ~n37041;
  assign n37043 = n34656 & ~n37037;
  assign n37044 = n37042 & ~n37043;
  assign n37045 = ~n37038 & ~n37039;
  assign n37046 = n37044 & n37045;
  assign n37047 = ~n36971 & ~n36973;
  assign n37048 = ~n36974 & ~n37047;
  assign n37049 = P1_P2_INSTQUEUE_REG_0__3_ & n36665;
  assign n37050 = P1_P2_INSTQUEUE_REG_1__3_ & n36668;
  assign n37051 = P1_P2_INSTQUEUE_REG_2__3_ & n36671;
  assign n37052 = P1_P2_INSTQUEUE_REG_3__3_ & n36674;
  assign n37053 = ~n37049 & ~n37050;
  assign n37054 = ~n37051 & n37053;
  assign n37055 = ~n37052 & n37054;
  assign n37056 = P1_P2_INSTQUEUE_REG_4__3_ & n36680;
  assign n37057 = P1_P2_INSTQUEUE_REG_5__3_ & n36682;
  assign n37058 = P1_P2_INSTQUEUE_REG_6__3_ & n36684;
  assign n37059 = P1_P2_INSTQUEUE_REG_7__3_ & n36686;
  assign n37060 = ~n37056 & ~n37057;
  assign n37061 = ~n37058 & n37060;
  assign n37062 = ~n37059 & n37061;
  assign n37063 = P1_P2_INSTQUEUE_REG_8__3_ & n36692;
  assign n37064 = P1_P2_INSTQUEUE_REG_9__3_ & n36694;
  assign n37065 = P1_P2_INSTQUEUE_REG_10__3_ & n36696;
  assign n37066 = P1_P2_INSTQUEUE_REG_11__3_ & n36698;
  assign n37067 = ~n37063 & ~n37064;
  assign n37068 = ~n37065 & n37067;
  assign n37069 = ~n37066 & n37068;
  assign n37070 = P1_P2_INSTQUEUE_REG_12__3_ & n36704;
  assign n37071 = P1_P2_INSTQUEUE_REG_13__3_ & n36706;
  assign n37072 = P1_P2_INSTQUEUE_REG_14__3_ & n36708;
  assign n37073 = P1_P2_INSTQUEUE_REG_15__3_ & n36710;
  assign n37074 = ~n37070 & ~n37071;
  assign n37075 = ~n37072 & n37074;
  assign n37076 = ~n37073 & n37075;
  assign n37077 = n37055 & n37062;
  assign n37078 = n37069 & n37077;
  assign n37079 = n37076 & n37078;
  assign n37080 = ~n36835 & ~n36955;
  assign n37081 = n37079 & ~n37080;
  assign n37082 = ~n37079 & n37080;
  assign n37083 = ~n37081 & ~n37082;
  assign n37084 = P1_P2_INSTADDRPOINTER_REG_3_ & ~n37083;
  assign n37085 = ~P1_P2_INSTADDRPOINTER_REG_3_ & n37083;
  assign n37086 = ~n37084 & ~n37085;
  assign n37087 = n37048 & ~n37086;
  assign n37088 = P1_P2_INSTADDRPOINTER_REG_3_ & n37083;
  assign n37089 = ~P1_P2_INSTADDRPOINTER_REG_3_ & ~n37083;
  assign n37090 = ~n37088 & ~n37089;
  assign n37091 = ~n37048 & ~n37090;
  assign n37092 = ~n37087 & ~n37091;
  assign n37093 = n36752 & ~n37092;
  assign n37094 = ~n36924 & ~n36973;
  assign n37095 = ~n36974 & ~n37094;
  assign n37096 = n37079 & n37080;
  assign n37097 = ~n37079 & ~n37080;
  assign n37098 = ~n37096 & ~n37097;
  assign n37099 = ~P1_P2_INSTADDRPOINTER_REG_3_ & n37098;
  assign n37100 = ~n37095 & ~n37099;
  assign n37101 = P1_P2_INSTADDRPOINTER_REG_3_ & ~n37098;
  assign n37102 = n37100 & ~n37101;
  assign n37103 = ~P1_P2_INSTADDRPOINTER_REG_3_ & ~n37098;
  assign n37104 = P1_P2_INSTADDRPOINTER_REG_3_ & n37098;
  assign n37105 = ~n37103 & ~n37104;
  assign n37106 = n37095 & n37105;
  assign n37107 = ~n37102 & ~n37106;
  assign n37108 = n36754 & n37107;
  assign n37109 = ~n37093 & ~n37108;
  assign n37110 = n36771 & ~n37029;
  assign n37111 = n36764 & ~n37029;
  assign n37112 = n36760 & ~n37029;
  assign n37113 = n34726 & ~n37029;
  assign n37114 = ~n37110 & ~n37111;
  assign n37115 = ~n37112 & n37114;
  assign n37116 = ~n37113 & n37115;
  assign n37117 = n34582 & ~n37037;
  assign n37118 = n34660 & ~n37037;
  assign n37119 = n34664 & ~n37037;
  assign n37120 = ~P1_P2_INSTADDRPOINTER_REG_3_ & n36990;
  assign n37121 = P1_P2_INSTADDRPOINTER_REG_3_ & ~n36990;
  assign n37122 = ~n37120 & ~n37121;
  assign n37123 = n34680 & n37122;
  assign n37124 = n34672 & n37122;
  assign n37125 = ~n37117 & ~n37118;
  assign n37126 = ~n37119 & n37125;
  assign n37127 = ~n37123 & n37126;
  assign n37128 = ~n37124 & n37127;
  assign n37129 = n37008 & ~n37011;
  assign n37130 = n37000 & n37079;
  assign n37131 = ~n37000 & ~n37079;
  assign n37132 = ~n37130 & ~n37131;
  assign n37133 = P1_P2_INSTADDRPOINTER_REG_3_ & n37132;
  assign n37134 = ~n37010 & n37132;
  assign n37135 = P1_P2_INSTADDRPOINTER_REG_3_ & ~n37010;
  assign n37136 = ~n37134 & ~n37135;
  assign n37137 = ~n37129 & ~n37133;
  assign n37138 = ~n37136 & n37137;
  assign n37139 = ~P1_P2_INSTADDRPOINTER_REG_3_ & n37132;
  assign n37140 = P1_P2_INSTADDRPOINTER_REG_3_ & ~n37132;
  assign n37141 = ~n37139 & ~n37140;
  assign n37142 = ~n37011 & n37141;
  assign n37143 = ~n37008 & ~n37010;
  assign n37144 = n37142 & ~n37143;
  assign n37145 = ~n37138 & ~n37144;
  assign n37146 = n34683 & n37145;
  assign n37147 = n37116 & n37128;
  assign n37148 = ~n37146 & n37147;
  assign n37149 = n37032 & ~n37033;
  assign n37150 = n37046 & n37149;
  assign n37151 = n37109 & n37150;
  assign n37152 = n37148 & n37151;
  assign n37153 = n36647 & ~n37152;
  assign n37154 = ~n37025 & ~n37026;
  assign n6566 = n37153 | ~n37154;
  assign n37156 = P1_P2_INSTADDRPOINTER_REG_4_ & n36646;
  assign n37157 = P1_P2_REIP_REG_4_ & n36791;
  assign n37158 = P1_P2_INSTADDRPOINTER_REG_3_ & n36991;
  assign n37159 = ~P1_P2_INSTADDRPOINTER_REG_4_ & n37158;
  assign n37160 = P1_P2_INSTADDRPOINTER_REG_4_ & ~n37158;
  assign n37161 = ~n37159 & ~n37160;
  assign n37162 = ~n34769 & ~n37161;
  assign n37163 = P1_P2_INSTADDRPOINTER_REG_3_ & n37034;
  assign n37164 = ~P1_P2_INSTADDRPOINTER_REG_4_ & n37163;
  assign n37165 = P1_P2_INSTADDRPOINTER_REG_4_ & ~n37163;
  assign n37166 = ~n37164 & ~n37165;
  assign n37167 = n34840 & ~n37166;
  assign n37168 = n34841 & ~n37166;
  assign n37169 = n36655 & ~n37161;
  assign n37170 = n36658 & ~n37161;
  assign n37171 = ~n37169 & ~n37170;
  assign n37172 = n34656 & ~n37166;
  assign n37173 = n37171 & ~n37172;
  assign n37174 = ~n37167 & ~n37168;
  assign n37175 = n37173 & n37174;
  assign n37176 = P1_P2_INSTQUEUE_REG_0__4_ & n36665;
  assign n37177 = P1_P2_INSTQUEUE_REG_1__4_ & n36668;
  assign n37178 = P1_P2_INSTQUEUE_REG_2__4_ & n36671;
  assign n37179 = P1_P2_INSTQUEUE_REG_3__4_ & n36674;
  assign n37180 = ~n37176 & ~n37177;
  assign n37181 = ~n37178 & n37180;
  assign n37182 = ~n37179 & n37181;
  assign n37183 = P1_P2_INSTQUEUE_REG_4__4_ & n36680;
  assign n37184 = P1_P2_INSTQUEUE_REG_5__4_ & n36682;
  assign n37185 = P1_P2_INSTQUEUE_REG_6__4_ & n36684;
  assign n37186 = P1_P2_INSTQUEUE_REG_7__4_ & n36686;
  assign n37187 = ~n37183 & ~n37184;
  assign n37188 = ~n37185 & n37187;
  assign n37189 = ~n37186 & n37188;
  assign n37190 = P1_P2_INSTQUEUE_REG_8__4_ & n36692;
  assign n37191 = P1_P2_INSTQUEUE_REG_9__4_ & n36694;
  assign n37192 = P1_P2_INSTQUEUE_REG_10__4_ & n36696;
  assign n37193 = P1_P2_INSTQUEUE_REG_11__4_ & n36698;
  assign n37194 = ~n37190 & ~n37191;
  assign n37195 = ~n37192 & n37194;
  assign n37196 = ~n37193 & n37195;
  assign n37197 = P1_P2_INSTQUEUE_REG_12__4_ & n36704;
  assign n37198 = P1_P2_INSTQUEUE_REG_13__4_ & n36706;
  assign n37199 = P1_P2_INSTQUEUE_REG_14__4_ & n36708;
  assign n37200 = P1_P2_INSTQUEUE_REG_15__4_ & n36710;
  assign n37201 = ~n37197 & ~n37198;
  assign n37202 = ~n37199 & n37201;
  assign n37203 = ~n37200 & n37202;
  assign n37204 = n37182 & n37189;
  assign n37205 = n37196 & n37204;
  assign n37206 = n37203 & n37205;
  assign n37207 = n37082 & n37206;
  assign n37208 = ~n37082 & ~n37206;
  assign n37209 = ~n37207 & ~n37208;
  assign n37210 = P1_P2_INSTADDRPOINTER_REG_4_ & ~n37209;
  assign n37211 = ~P1_P2_INSTADDRPOINTER_REG_4_ & n37209;
  assign n37212 = ~n37210 & ~n37211;
  assign n37213 = ~n37100 & ~n37101;
  assign n37214 = n37212 & ~n37213;
  assign n37215 = ~P1_P2_INSTADDRPOINTER_REG_4_ & ~n37209;
  assign n37216 = P1_P2_INSTADDRPOINTER_REG_4_ & n37209;
  assign n37217 = ~n37215 & ~n37216;
  assign n37218 = ~n37101 & n37217;
  assign n37219 = ~n37100 & n37218;
  assign n37220 = ~n37214 & ~n37219;
  assign n37221 = n36754 & n37220;
  assign n37222 = n34879 & ~n37161;
  assign n37223 = n34722 & ~n37161;
  assign n37224 = ~n37222 & ~n37223;
  assign n37225 = ~n36973 & ~n37089;
  assign n37226 = ~n36839 & ~n36969;
  assign n37227 = ~n36974 & n37226;
  assign n37228 = ~n36889 & n37227;
  assign n37229 = n37225 & ~n37228;
  assign n37230 = ~n37088 & ~n37229;
  assign n37231 = n37082 & ~n37206;
  assign n37232 = ~n37082 & n37206;
  assign n37233 = ~n37231 & ~n37232;
  assign n37234 = P1_P2_INSTADDRPOINTER_REG_4_ & ~n37233;
  assign n37235 = ~P1_P2_INSTADDRPOINTER_REG_4_ & n37233;
  assign n37236 = ~n37234 & ~n37235;
  assign n37237 = n37230 & ~n37236;
  assign n37238 = P1_P2_INSTADDRPOINTER_REG_4_ & n37233;
  assign n37239 = ~P1_P2_INSTADDRPOINTER_REG_4_ & ~n37233;
  assign n37240 = ~n37238 & ~n37239;
  assign n37241 = ~n37230 & ~n37240;
  assign n37242 = ~n37237 & ~n37241;
  assign n37243 = n36752 & ~n37242;
  assign n37244 = n37224 & ~n37243;
  assign n37245 = n36771 & ~n37161;
  assign n37246 = n36764 & ~n37161;
  assign n37247 = n36760 & ~n37161;
  assign n37248 = n34726 & ~n37161;
  assign n37249 = ~n37245 & ~n37246;
  assign n37250 = ~n37247 & n37249;
  assign n37251 = ~n37248 & n37250;
  assign n37252 = n34582 & ~n37166;
  assign n37253 = n34660 & ~n37166;
  assign n37254 = n34664 & ~n37166;
  assign n37255 = ~P1_P2_INSTADDRPOINTER_REG_4_ & n37121;
  assign n37256 = P1_P2_INSTADDRPOINTER_REG_4_ & ~n37121;
  assign n37257 = ~n37255 & ~n37256;
  assign n37258 = n34680 & ~n37257;
  assign n37259 = n34672 & ~n37257;
  assign n37260 = ~n37252 & ~n37253;
  assign n37261 = ~n37254 & n37260;
  assign n37262 = ~n37258 & n37261;
  assign n37263 = ~n37259 & n37262;
  assign n37264 = n37131 & n37206;
  assign n37265 = ~n37131 & ~n37206;
  assign n37266 = ~n37264 & ~n37265;
  assign n37267 = ~P1_P2_INSTADDRPOINTER_REG_4_ & ~n37266;
  assign n37268 = P1_P2_INSTADDRPOINTER_REG_4_ & n37266;
  assign n37269 = ~n37267 & ~n37268;
  assign n37270 = n37011 & n37132;
  assign n37271 = ~n37011 & ~n37132;
  assign n37272 = P1_P2_INSTADDRPOINTER_REG_3_ & ~n37271;
  assign n37273 = ~n37270 & ~n37272;
  assign n37274 = ~n37008 & ~n37136;
  assign n37275 = n37273 & ~n37274;
  assign n37276 = ~n37269 & n37275;
  assign n37277 = ~P1_P2_INSTADDRPOINTER_REG_4_ & n37266;
  assign n37278 = P1_P2_INSTADDRPOINTER_REG_4_ & ~n37266;
  assign n37279 = ~n37277 & ~n37278;
  assign n37280 = ~n37275 & ~n37279;
  assign n37281 = ~n37276 & ~n37280;
  assign n37282 = n34683 & ~n37281;
  assign n37283 = n37251 & n37263;
  assign n37284 = ~n37282 & n37283;
  assign n37285 = ~n37162 & n37175;
  assign n37286 = ~n37221 & n37285;
  assign n37287 = n37244 & n37286;
  assign n37288 = n37284 & n37287;
  assign n37289 = n36647 & ~n37288;
  assign n37290 = ~n37156 & ~n37157;
  assign n6571 = n37289 | ~n37290;
  assign n37292 = P1_P2_INSTADDRPOINTER_REG_5_ & n36646;
  assign n37293 = P1_P2_REIP_REG_5_ & n36791;
  assign n37294 = P1_P2_INSTADDRPOINTER_REG_4_ & n37163;
  assign n37295 = ~P1_P2_INSTADDRPOINTER_REG_5_ & n37294;
  assign n37296 = P1_P2_INSTADDRPOINTER_REG_5_ & ~n37294;
  assign n37297 = ~n37295 & ~n37296;
  assign n37298 = n34840 & ~n37297;
  assign n37299 = n34841 & ~n37297;
  assign n37300 = P1_P2_INSTADDRPOINTER_REG_4_ & n37158;
  assign n37301 = ~P1_P2_INSTADDRPOINTER_REG_5_ & n37300;
  assign n37302 = P1_P2_INSTADDRPOINTER_REG_5_ & ~n37300;
  assign n37303 = ~n37301 & ~n37302;
  assign n37304 = n36655 & ~n37303;
  assign n37305 = n36658 & ~n37303;
  assign n37306 = ~n37304 & ~n37305;
  assign n37307 = n34656 & ~n37297;
  assign n37308 = n37306 & ~n37307;
  assign n37309 = ~n37298 & ~n37299;
  assign n37310 = n37308 & n37309;
  assign n37311 = ~n34769 & ~n37303;
  assign n37312 = n37088 & ~n37239;
  assign n37313 = ~n37238 & ~n37312;
  assign n37314 = n37225 & ~n37239;
  assign n37315 = ~n37228 & n37314;
  assign n37316 = n37313 & ~n37315;
  assign n37317 = P1_P2_INSTQUEUE_REG_0__5_ & n36665;
  assign n37318 = P1_P2_INSTQUEUE_REG_1__5_ & n36668;
  assign n37319 = P1_P2_INSTQUEUE_REG_2__5_ & n36671;
  assign n37320 = P1_P2_INSTQUEUE_REG_3__5_ & n36674;
  assign n37321 = ~n37317 & ~n37318;
  assign n37322 = ~n37319 & n37321;
  assign n37323 = ~n37320 & n37322;
  assign n37324 = P1_P2_INSTQUEUE_REG_4__5_ & n36680;
  assign n37325 = P1_P2_INSTQUEUE_REG_5__5_ & n36682;
  assign n37326 = P1_P2_INSTQUEUE_REG_6__5_ & n36684;
  assign n37327 = P1_P2_INSTQUEUE_REG_7__5_ & n36686;
  assign n37328 = ~n37324 & ~n37325;
  assign n37329 = ~n37326 & n37328;
  assign n37330 = ~n37327 & n37329;
  assign n37331 = P1_P2_INSTQUEUE_REG_8__5_ & n36692;
  assign n37332 = P1_P2_INSTQUEUE_REG_9__5_ & n36694;
  assign n37333 = P1_P2_INSTQUEUE_REG_10__5_ & n36696;
  assign n37334 = P1_P2_INSTQUEUE_REG_11__5_ & n36698;
  assign n37335 = ~n37331 & ~n37332;
  assign n37336 = ~n37333 & n37335;
  assign n37337 = ~n37334 & n37336;
  assign n37338 = P1_P2_INSTQUEUE_REG_12__5_ & n36704;
  assign n37339 = P1_P2_INSTQUEUE_REG_13__5_ & n36706;
  assign n37340 = P1_P2_INSTQUEUE_REG_14__5_ & n36708;
  assign n37341 = P1_P2_INSTQUEUE_REG_15__5_ & n36710;
  assign n37342 = ~n37338 & ~n37339;
  assign n37343 = ~n37340 & n37342;
  assign n37344 = ~n37341 & n37343;
  assign n37345 = n37323 & n37330;
  assign n37346 = n37337 & n37345;
  assign n37347 = n37344 & n37346;
  assign n37348 = ~n37231 & n37347;
  assign n37349 = ~n37206 & ~n37347;
  assign n37350 = n37082 & n37349;
  assign n37351 = ~n37348 & ~n37350;
  assign n37352 = P1_P2_INSTADDRPOINTER_REG_5_ & ~n37351;
  assign n37353 = ~P1_P2_INSTADDRPOINTER_REG_5_ & n37351;
  assign n37354 = ~n37352 & ~n37353;
  assign n37355 = n37316 & ~n37354;
  assign n37356 = ~n37316 & n37354;
  assign n37357 = ~n37355 & ~n37356;
  assign n37358 = n36752 & ~n37357;
  assign n37359 = n34879 & ~n37303;
  assign n37360 = n34722 & ~n37303;
  assign n37361 = ~n37359 & ~n37360;
  assign n37362 = n37101 & ~n37211;
  assign n37363 = ~n37210 & ~n37362;
  assign n37364 = ~n37099 & ~n37211;
  assign n37365 = ~n37095 & n37364;
  assign n37366 = n37363 & ~n37365;
  assign n37367 = n37231 & n37347;
  assign n37368 = ~n37231 & ~n37347;
  assign n37369 = ~n37367 & ~n37368;
  assign n37370 = ~P1_P2_INSTADDRPOINTER_REG_5_ & ~n37369;
  assign n37371 = P1_P2_INSTADDRPOINTER_REG_5_ & n37369;
  assign n37372 = ~n37370 & ~n37371;
  assign n37373 = n37366 & ~n37372;
  assign n37374 = ~n37366 & n37372;
  assign n37375 = ~n37373 & ~n37374;
  assign n37376 = n36754 & ~n37375;
  assign n37377 = n37361 & ~n37376;
  assign n37378 = n36771 & ~n37303;
  assign n37379 = n36764 & ~n37303;
  assign n37380 = n36760 & ~n37303;
  assign n37381 = n34726 & ~n37303;
  assign n37382 = ~n37378 & ~n37379;
  assign n37383 = ~n37380 & n37382;
  assign n37384 = ~n37381 & n37383;
  assign n37385 = n34582 & ~n37297;
  assign n37386 = n34660 & ~n37297;
  assign n37387 = n34664 & ~n37297;
  assign n37388 = P1_P2_INSTADDRPOINTER_REG_4_ & n37121;
  assign n37389 = ~P1_P2_INSTADDRPOINTER_REG_5_ & n37388;
  assign n37390 = P1_P2_INSTADDRPOINTER_REG_5_ & ~n37388;
  assign n37391 = ~n37389 & ~n37390;
  assign n37392 = n34680 & ~n37391;
  assign n37393 = n34672 & ~n37391;
  assign n37394 = ~n37385 & ~n37386;
  assign n37395 = ~n37387 & n37394;
  assign n37396 = ~n37392 & n37395;
  assign n37397 = ~n37393 & n37396;
  assign n37398 = n37131 & ~n37206;
  assign n37399 = n37347 & n37398;
  assign n37400 = ~n37347 & ~n37398;
  assign n37401 = ~n37399 & ~n37400;
  assign n37402 = P1_P2_INSTADDRPOINTER_REG_5_ & ~n37401;
  assign n37403 = ~P1_P2_INSTADDRPOINTER_REG_5_ & n37401;
  assign n37404 = ~n37277 & ~n37403;
  assign n37405 = ~n37402 & n37404;
  assign n37406 = n37275 & ~n37278;
  assign n37407 = n37405 & ~n37406;
  assign n37408 = ~P1_P2_INSTADDRPOINTER_REG_5_ & ~n37401;
  assign n37409 = P1_P2_INSTADDRPOINTER_REG_5_ & n37401;
  assign n37410 = ~n37408 & ~n37409;
  assign n37411 = ~n37278 & n37410;
  assign n37412 = ~n37275 & ~n37277;
  assign n37413 = n37411 & ~n37412;
  assign n37414 = ~n37407 & ~n37413;
  assign n37415 = n34683 & n37414;
  assign n37416 = n37384 & n37397;
  assign n37417 = ~n37415 & n37416;
  assign n37418 = n37310 & ~n37311;
  assign n37419 = ~n37358 & n37418;
  assign n37420 = n37377 & n37419;
  assign n37421 = n37417 & n37420;
  assign n37422 = n36647 & ~n37421;
  assign n37423 = ~n37292 & ~n37293;
  assign n6576 = n37422 | ~n37423;
  assign n37425 = P1_P2_INSTADDRPOINTER_REG_6_ & n36646;
  assign n37426 = P1_P2_REIP_REG_6_ & n36791;
  assign n37427 = P1_P2_INSTADDRPOINTER_REG_5_ & n37294;
  assign n37428 = ~P1_P2_INSTADDRPOINTER_REG_6_ & n37427;
  assign n37429 = P1_P2_INSTADDRPOINTER_REG_6_ & ~n37427;
  assign n37430 = ~n37428 & ~n37429;
  assign n37431 = n34840 & ~n37430;
  assign n37432 = n34841 & ~n37430;
  assign n37433 = P1_P2_INSTADDRPOINTER_REG_5_ & n37300;
  assign n37434 = ~P1_P2_INSTADDRPOINTER_REG_6_ & n37433;
  assign n37435 = P1_P2_INSTADDRPOINTER_REG_6_ & ~n37433;
  assign n37436 = ~n37434 & ~n37435;
  assign n37437 = n36655 & ~n37436;
  assign n37438 = n36658 & ~n37436;
  assign n37439 = ~n37437 & ~n37438;
  assign n37440 = n34656 & ~n37430;
  assign n37441 = n37439 & ~n37440;
  assign n37442 = ~n37431 & ~n37432;
  assign n37443 = n37441 & n37442;
  assign n37444 = ~n34769 & ~n37436;
  assign n37445 = ~P1_P2_INSTADDRPOINTER_REG_5_ & ~n37351;
  assign n37446 = ~n37316 & ~n37445;
  assign n37447 = P1_P2_INSTADDRPOINTER_REG_5_ & n37351;
  assign n37448 = ~n37446 & ~n37447;
  assign n37449 = P1_P2_INSTQUEUE_REG_0__6_ & n36665;
  assign n37450 = P1_P2_INSTQUEUE_REG_1__6_ & n36668;
  assign n37451 = P1_P2_INSTQUEUE_REG_2__6_ & n36671;
  assign n37452 = P1_P2_INSTQUEUE_REG_3__6_ & n36674;
  assign n37453 = ~n37449 & ~n37450;
  assign n37454 = ~n37451 & n37453;
  assign n37455 = ~n37452 & n37454;
  assign n37456 = P1_P2_INSTQUEUE_REG_4__6_ & n36680;
  assign n37457 = P1_P2_INSTQUEUE_REG_5__6_ & n36682;
  assign n37458 = P1_P2_INSTQUEUE_REG_6__6_ & n36684;
  assign n37459 = P1_P2_INSTQUEUE_REG_7__6_ & n36686;
  assign n37460 = ~n37456 & ~n37457;
  assign n37461 = ~n37458 & n37460;
  assign n37462 = ~n37459 & n37461;
  assign n37463 = P1_P2_INSTQUEUE_REG_8__6_ & n36692;
  assign n37464 = P1_P2_INSTQUEUE_REG_9__6_ & n36694;
  assign n37465 = P1_P2_INSTQUEUE_REG_10__6_ & n36696;
  assign n37466 = P1_P2_INSTQUEUE_REG_11__6_ & n36698;
  assign n37467 = ~n37463 & ~n37464;
  assign n37468 = ~n37465 & n37467;
  assign n37469 = ~n37466 & n37468;
  assign n37470 = P1_P2_INSTQUEUE_REG_12__6_ & n36704;
  assign n37471 = P1_P2_INSTQUEUE_REG_13__6_ & n36706;
  assign n37472 = P1_P2_INSTQUEUE_REG_14__6_ & n36708;
  assign n37473 = P1_P2_INSTQUEUE_REG_15__6_ & n36710;
  assign n37474 = ~n37470 & ~n37471;
  assign n37475 = ~n37472 & n37474;
  assign n37476 = ~n37473 & n37475;
  assign n37477 = n37455 & n37462;
  assign n37478 = n37469 & n37477;
  assign n37479 = n37476 & n37478;
  assign n37480 = n37350 & ~n37479;
  assign n37481 = ~n37350 & n37479;
  assign n37482 = ~n37480 & ~n37481;
  assign n37483 = P1_P2_INSTADDRPOINTER_REG_6_ & ~n37482;
  assign n37484 = ~P1_P2_INSTADDRPOINTER_REG_6_ & n37482;
  assign n37485 = ~n37483 & ~n37484;
  assign n37486 = n37448 & ~n37485;
  assign n37487 = ~n37448 & n37485;
  assign n37488 = ~n37486 & ~n37487;
  assign n37489 = n36752 & ~n37488;
  assign n37490 = n34879 & ~n37436;
  assign n37491 = n34722 & ~n37436;
  assign n37492 = ~n37490 & ~n37491;
  assign n37493 = ~n37366 & ~n37369;
  assign n37494 = P1_P2_INSTADDRPOINTER_REG_5_ & ~n37366;
  assign n37495 = P1_P2_INSTADDRPOINTER_REG_5_ & ~n37369;
  assign n37496 = ~n37493 & ~n37494;
  assign n37497 = ~n37495 & n37496;
  assign n37498 = n37231 & ~n37347;
  assign n37499 = n37479 & n37498;
  assign n37500 = ~n37479 & ~n37498;
  assign n37501 = ~n37499 & ~n37500;
  assign n37502 = ~P1_P2_INSTADDRPOINTER_REG_6_ & ~n37501;
  assign n37503 = P1_P2_INSTADDRPOINTER_REG_6_ & n37501;
  assign n37504 = ~n37502 & ~n37503;
  assign n37505 = n37497 & ~n37504;
  assign n37506 = ~n37497 & n37504;
  assign n37507 = ~n37505 & ~n37506;
  assign n37508 = n36754 & ~n37507;
  assign n37509 = n37492 & ~n37508;
  assign n37510 = n36771 & ~n37436;
  assign n37511 = n36764 & ~n37436;
  assign n37512 = n36760 & ~n37436;
  assign n37513 = n34726 & ~n37436;
  assign n37514 = ~n37510 & ~n37511;
  assign n37515 = ~n37512 & n37514;
  assign n37516 = ~n37513 & n37515;
  assign n37517 = n34582 & ~n37430;
  assign n37518 = n34660 & ~n37430;
  assign n37519 = n34664 & ~n37430;
  assign n37520 = P1_P2_INSTADDRPOINTER_REG_5_ & n37388;
  assign n37521 = ~P1_P2_INSTADDRPOINTER_REG_6_ & n37520;
  assign n37522 = P1_P2_INSTADDRPOINTER_REG_6_ & ~n37520;
  assign n37523 = ~n37521 & ~n37522;
  assign n37524 = n34680 & ~n37523;
  assign n37525 = n34672 & ~n37523;
  assign n37526 = ~n37517 & ~n37518;
  assign n37527 = ~n37519 & n37526;
  assign n37528 = ~n37524 & n37527;
  assign n37529 = ~n37525 & n37528;
  assign n37530 = n37278 & ~n37401;
  assign n37531 = ~n37278 & n37401;
  assign n37532 = P1_P2_INSTADDRPOINTER_REG_5_ & ~n37531;
  assign n37533 = ~n37530 & ~n37532;
  assign n37534 = ~n37275 & n37404;
  assign n37535 = n37533 & ~n37534;
  assign n37536 = ~n37347 & n37398;
  assign n37537 = n37479 & n37536;
  assign n37538 = ~n37479 & ~n37536;
  assign n37539 = ~n37537 & ~n37538;
  assign n37540 = ~P1_P2_INSTADDRPOINTER_REG_6_ & ~n37539;
  assign n37541 = P1_P2_INSTADDRPOINTER_REG_6_ & n37539;
  assign n37542 = ~n37540 & ~n37541;
  assign n37543 = n37535 & ~n37542;
  assign n37544 = ~n37535 & n37542;
  assign n37545 = ~n37543 & ~n37544;
  assign n37546 = n34683 & ~n37545;
  assign n37547 = n37516 & n37529;
  assign n37548 = ~n37546 & n37547;
  assign n37549 = n37443 & ~n37444;
  assign n37550 = ~n37489 & n37549;
  assign n37551 = n37509 & n37550;
  assign n37552 = n37548 & n37551;
  assign n37553 = n36647 & ~n37552;
  assign n37554 = ~n37425 & ~n37426;
  assign n6581 = n37553 | ~n37554;
  assign n37556 = P1_P2_INSTADDRPOINTER_REG_7_ & n36646;
  assign n37557 = P1_P2_REIP_REG_7_ & n36791;
  assign n37558 = P1_P2_INSTADDRPOINTER_REG_6_ & n37427;
  assign n37559 = ~P1_P2_INSTADDRPOINTER_REG_7_ & n37558;
  assign n37560 = P1_P2_INSTADDRPOINTER_REG_7_ & ~n37558;
  assign n37561 = ~n37559 & ~n37560;
  assign n37562 = n34840 & ~n37561;
  assign n37563 = n34841 & ~n37561;
  assign n37564 = P1_P2_INSTADDRPOINTER_REG_6_ & n37433;
  assign n37565 = ~P1_P2_INSTADDRPOINTER_REG_7_ & n37564;
  assign n37566 = P1_P2_INSTADDRPOINTER_REG_7_ & ~n37564;
  assign n37567 = ~n37565 & ~n37566;
  assign n37568 = n36655 & ~n37567;
  assign n37569 = n36658 & ~n37567;
  assign n37570 = ~n37568 & ~n37569;
  assign n37571 = n34656 & ~n37561;
  assign n37572 = n37570 & ~n37571;
  assign n37573 = ~n37562 & ~n37563;
  assign n37574 = n37572 & n37573;
  assign n37575 = ~n34769 & ~n37567;
  assign n37576 = P1_P2_INSTADDRPOINTER_REG_6_ & n37482;
  assign n37577 = ~P1_P2_INSTADDRPOINTER_REG_6_ & ~n37482;
  assign n37578 = ~n37448 & ~n37577;
  assign n37579 = ~n37576 & ~n37578;
  assign n37580 = n36751 & ~n37480;
  assign n37581 = ~n36751 & ~n37479;
  assign n37582 = n37350 & n37581;
  assign n37583 = ~n37580 & ~n37582;
  assign n37584 = P1_P2_INSTADDRPOINTER_REG_7_ & ~n37583;
  assign n37585 = ~P1_P2_INSTADDRPOINTER_REG_7_ & n37583;
  assign n37586 = ~n37584 & ~n37585;
  assign n37587 = n37579 & ~n37586;
  assign n37588 = ~n37579 & n37586;
  assign n37589 = ~n37587 & ~n37588;
  assign n37590 = n36752 & ~n37589;
  assign n37591 = n34879 & ~n37567;
  assign n37592 = n34722 & ~n37567;
  assign n37593 = ~n37591 & ~n37592;
  assign n37594 = P1_P2_INSTADDRPOINTER_REG_6_ & ~n37501;
  assign n37595 = ~P1_P2_INSTADDRPOINTER_REG_6_ & n37501;
  assign n37596 = ~n37497 & ~n37595;
  assign n37597 = ~n37594 & ~n37596;
  assign n37598 = ~n37479 & n37498;
  assign n37599 = n36751 & n37598;
  assign n37600 = ~n36751 & ~n37598;
  assign n37601 = ~n37599 & ~n37600;
  assign n37602 = ~P1_P2_INSTADDRPOINTER_REG_7_ & ~n37601;
  assign n37603 = P1_P2_INSTADDRPOINTER_REG_7_ & n37601;
  assign n37604 = ~n37602 & ~n37603;
  assign n37605 = n37597 & ~n37604;
  assign n37606 = ~n37597 & n37604;
  assign n37607 = ~n37605 & ~n37606;
  assign n37608 = n36754 & ~n37607;
  assign n37609 = n37593 & ~n37608;
  assign n37610 = n36771 & ~n37567;
  assign n37611 = n36764 & ~n37567;
  assign n37612 = n36760 & ~n37567;
  assign n37613 = n34726 & ~n37567;
  assign n37614 = ~n37610 & ~n37611;
  assign n37615 = ~n37612 & n37614;
  assign n37616 = ~n37613 & n37615;
  assign n37617 = n34582 & ~n37561;
  assign n37618 = n34660 & ~n37561;
  assign n37619 = n34664 & ~n37561;
  assign n37620 = P1_P2_INSTADDRPOINTER_REG_6_ & n37520;
  assign n37621 = ~P1_P2_INSTADDRPOINTER_REG_7_ & n37620;
  assign n37622 = P1_P2_INSTADDRPOINTER_REG_7_ & ~n37620;
  assign n37623 = ~n37621 & ~n37622;
  assign n37624 = n34680 & ~n37623;
  assign n37625 = n34672 & ~n37623;
  assign n37626 = ~n37617 & ~n37618;
  assign n37627 = ~n37619 & n37626;
  assign n37628 = ~n37624 & n37627;
  assign n37629 = ~n37625 & n37628;
  assign n37630 = P1_P2_INSTADDRPOINTER_REG_6_ & ~n37539;
  assign n37631 = ~P1_P2_INSTADDRPOINTER_REG_6_ & n37539;
  assign n37632 = ~n37535 & ~n37631;
  assign n37633 = ~n37630 & ~n37632;
  assign n37634 = ~n37479 & n37536;
  assign n37635 = n36751 & n37634;
  assign n37636 = ~n36751 & ~n37634;
  assign n37637 = ~n37635 & ~n37636;
  assign n37638 = ~P1_P2_INSTADDRPOINTER_REG_7_ & ~n37637;
  assign n37639 = P1_P2_INSTADDRPOINTER_REG_7_ & n37637;
  assign n37640 = ~n37638 & ~n37639;
  assign n37641 = n37633 & ~n37640;
  assign n37642 = ~n37633 & n37640;
  assign n37643 = ~n37641 & ~n37642;
  assign n37644 = n34683 & ~n37643;
  assign n37645 = n37616 & n37629;
  assign n37646 = ~n37644 & n37645;
  assign n37647 = n37574 & ~n37575;
  assign n37648 = ~n37590 & n37647;
  assign n37649 = n37609 & n37648;
  assign n37650 = n37646 & n37649;
  assign n37651 = n36647 & ~n37650;
  assign n37652 = ~n37556 & ~n37557;
  assign n6586 = n37651 | ~n37652;
  assign n37654 = P1_P2_INSTADDRPOINTER_REG_8_ & n36646;
  assign n37655 = P1_P2_REIP_REG_8_ & n36791;
  assign n37656 = P1_P2_INSTADDRPOINTER_REG_7_ & n37558;
  assign n37657 = ~P1_P2_INSTADDRPOINTER_REG_8_ & n37656;
  assign n37658 = P1_P2_INSTADDRPOINTER_REG_8_ & ~n37656;
  assign n37659 = ~n37657 & ~n37658;
  assign n37660 = n34840 & ~n37659;
  assign n37661 = n34841 & ~n37659;
  assign n37662 = n34656 & ~n37659;
  assign n37663 = P1_P2_INSTADDRPOINTER_REG_7_ & n37564;
  assign n37664 = ~P1_P2_INSTADDRPOINTER_REG_8_ & n37663;
  assign n37665 = P1_P2_INSTADDRPOINTER_REG_8_ & ~n37663;
  assign n37666 = ~n37664 & ~n37665;
  assign n37667 = n36658 & ~n37666;
  assign n37668 = n36655 & ~n37666;
  assign n37669 = ~n37662 & ~n37667;
  assign n37670 = ~n37668 & n37669;
  assign n37671 = ~n37660 & ~n37661;
  assign n37672 = n37670 & n37671;
  assign n37673 = ~n34769 & ~n37666;
  assign n37674 = ~P1_P2_INSTADDRPOINTER_REG_7_ & ~n37583;
  assign n37675 = ~n37579 & ~n37674;
  assign n37676 = P1_P2_INSTADDRPOINTER_REG_7_ & n37583;
  assign n37677 = ~n37675 & ~n37676;
  assign n37678 = ~P1_P2_INSTADDRPOINTER_REG_8_ & ~n37582;
  assign n37679 = P1_P2_INSTADDRPOINTER_REG_8_ & n37582;
  assign n37680 = ~n37678 & ~n37679;
  assign n37681 = n37677 & ~n37680;
  assign n37682 = ~n37677 & n37680;
  assign n37683 = ~n37681 & ~n37682;
  assign n37684 = n36752 & ~n37683;
  assign n37685 = n34879 & ~n37666;
  assign n37686 = n34722 & ~n37666;
  assign n37687 = ~n37685 & ~n37686;
  assign n37688 = ~n37597 & ~n37601;
  assign n37689 = P1_P2_INSTADDRPOINTER_REG_7_ & ~n37597;
  assign n37690 = P1_P2_INSTADDRPOINTER_REG_7_ & ~n37601;
  assign n37691 = ~n37688 & ~n37689;
  assign n37692 = ~n37690 & n37691;
  assign n37693 = n37498 & n37581;
  assign n37694 = ~P1_P2_INSTADDRPOINTER_REG_8_ & n37693;
  assign n37695 = P1_P2_INSTADDRPOINTER_REG_8_ & ~n37693;
  assign n37696 = ~n37694 & ~n37695;
  assign n37697 = n37692 & ~n37696;
  assign n37698 = ~n37692 & n37696;
  assign n37699 = ~n37697 & ~n37698;
  assign n37700 = n36754 & ~n37699;
  assign n37701 = n37687 & ~n37700;
  assign n37702 = n36771 & ~n37666;
  assign n37703 = n34726 & ~n37666;
  assign n37704 = n36760 & ~n37666;
  assign n37705 = n36764 & ~n37666;
  assign n37706 = ~n37702 & ~n37703;
  assign n37707 = ~n37704 & n37706;
  assign n37708 = ~n37705 & n37707;
  assign n37709 = n34582 & ~n37659;
  assign n37710 = n34660 & ~n37659;
  assign n37711 = n34664 & ~n37659;
  assign n37712 = P1_P2_INSTADDRPOINTER_REG_7_ & n37620;
  assign n37713 = ~P1_P2_INSTADDRPOINTER_REG_8_ & n37712;
  assign n37714 = P1_P2_INSTADDRPOINTER_REG_8_ & ~n37712;
  assign n37715 = ~n37713 & ~n37714;
  assign n37716 = n34680 & ~n37715;
  assign n37717 = n34672 & ~n37715;
  assign n37718 = ~n37709 & ~n37710;
  assign n37719 = ~n37711 & n37718;
  assign n37720 = ~n37716 & n37719;
  assign n37721 = ~n37717 & n37720;
  assign n37722 = ~n37633 & ~n37637;
  assign n37723 = P1_P2_INSTADDRPOINTER_REG_7_ & ~n37633;
  assign n37724 = P1_P2_INSTADDRPOINTER_REG_7_ & ~n37637;
  assign n37725 = ~n37722 & ~n37723;
  assign n37726 = ~n37724 & n37725;
  assign n37727 = n37536 & n37581;
  assign n37728 = ~P1_P2_INSTADDRPOINTER_REG_8_ & n37727;
  assign n37729 = P1_P2_INSTADDRPOINTER_REG_8_ & ~n37727;
  assign n37730 = ~n37728 & ~n37729;
  assign n37731 = n37726 & ~n37730;
  assign n37732 = ~n37726 & n37730;
  assign n37733 = ~n37731 & ~n37732;
  assign n37734 = n34683 & ~n37733;
  assign n37735 = n37708 & n37721;
  assign n37736 = ~n37734 & n37735;
  assign n37737 = n37672 & ~n37673;
  assign n37738 = ~n37684 & n37737;
  assign n37739 = n37701 & n37738;
  assign n37740 = n37736 & n37739;
  assign n37741 = n36647 & ~n37740;
  assign n37742 = ~n37654 & ~n37655;
  assign n6591 = n37741 | ~n37742;
  assign n37744 = P1_P2_INSTADDRPOINTER_REG_9_ & n36646;
  assign n37745 = P1_P2_REIP_REG_9_ & n36791;
  assign n37746 = P1_P2_INSTADDRPOINTER_REG_8_ & n37656;
  assign n37747 = ~P1_P2_INSTADDRPOINTER_REG_9_ & n37746;
  assign n37748 = P1_P2_INSTADDRPOINTER_REG_9_ & ~n37746;
  assign n37749 = ~n37747 & ~n37748;
  assign n37750 = n34840 & ~n37749;
  assign n37751 = n34841 & ~n37749;
  assign n37752 = P1_P2_INSTADDRPOINTER_REG_8_ & n37663;
  assign n37753 = ~P1_P2_INSTADDRPOINTER_REG_9_ & n37752;
  assign n37754 = P1_P2_INSTADDRPOINTER_REG_9_ & ~n37752;
  assign n37755 = ~n37753 & ~n37754;
  assign n37756 = n36655 & ~n37755;
  assign n37757 = n34656 & ~n37749;
  assign n37758 = n36658 & ~n37755;
  assign n37759 = ~n37757 & ~n37758;
  assign n37760 = ~n37750 & ~n37751;
  assign n37761 = ~n37756 & n37760;
  assign n37762 = n37759 & n37761;
  assign n37763 = ~n34769 & ~n37755;
  assign n37764 = ~P1_P2_INSTADDRPOINTER_REG_8_ & n37582;
  assign n37765 = ~n37677 & ~n37764;
  assign n37766 = P1_P2_INSTADDRPOINTER_REG_8_ & ~n37582;
  assign n37767 = ~n37765 & ~n37766;
  assign n37768 = P1_P2_INSTADDRPOINTER_REG_9_ & n37582;
  assign n37769 = ~P1_P2_INSTADDRPOINTER_REG_9_ & ~n37582;
  assign n37770 = ~n37768 & ~n37769;
  assign n37771 = n37767 & ~n37770;
  assign n37772 = P1_P2_INSTADDRPOINTER_REG_9_ & ~n37582;
  assign n37773 = ~P1_P2_INSTADDRPOINTER_REG_9_ & n37582;
  assign n37774 = ~n37772 & ~n37773;
  assign n37775 = ~n37767 & ~n37774;
  assign n37776 = ~n37771 & ~n37775;
  assign n37777 = n36752 & ~n37776;
  assign n37778 = n34879 & ~n37755;
  assign n37779 = n34722 & ~n37755;
  assign n37780 = ~n37778 & ~n37779;
  assign n37781 = P1_P2_INSTADDRPOINTER_REG_8_ & n37693;
  assign n37782 = ~P1_P2_INSTADDRPOINTER_REG_8_ & ~n37693;
  assign n37783 = ~n37692 & ~n37782;
  assign n37784 = ~n37781 & ~n37783;
  assign n37785 = ~P1_P2_INSTADDRPOINTER_REG_9_ & n37784;
  assign n37786 = P1_P2_INSTADDRPOINTER_REG_9_ & ~n37784;
  assign n37787 = ~n37785 & ~n37786;
  assign n37788 = n36754 & n37787;
  assign n37789 = n37780 & ~n37788;
  assign n37790 = n36771 & ~n37755;
  assign n37791 = n34726 & ~n37755;
  assign n37792 = n36760 & ~n37755;
  assign n37793 = n36764 & ~n37755;
  assign n37794 = ~n37790 & ~n37791;
  assign n37795 = ~n37792 & n37794;
  assign n37796 = ~n37793 & n37795;
  assign n37797 = n34582 & ~n37749;
  assign n37798 = n34660 & ~n37749;
  assign n37799 = n34664 & ~n37749;
  assign n37800 = P1_P2_INSTADDRPOINTER_REG_8_ & n37712;
  assign n37801 = ~P1_P2_INSTADDRPOINTER_REG_9_ & n37800;
  assign n37802 = P1_P2_INSTADDRPOINTER_REG_9_ & ~n37800;
  assign n37803 = ~n37801 & ~n37802;
  assign n37804 = n34680 & ~n37803;
  assign n37805 = n34672 & ~n37803;
  assign n37806 = ~n37797 & ~n37798;
  assign n37807 = ~n37799 & n37806;
  assign n37808 = ~n37804 & n37807;
  assign n37809 = ~n37805 & n37808;
  assign n37810 = P1_P2_INSTADDRPOINTER_REG_8_ & n37727;
  assign n37811 = ~P1_P2_INSTADDRPOINTER_REG_8_ & ~n37727;
  assign n37812 = ~n37726 & ~n37811;
  assign n37813 = ~n37810 & ~n37812;
  assign n37814 = ~P1_P2_INSTADDRPOINTER_REG_9_ & n37813;
  assign n37815 = P1_P2_INSTADDRPOINTER_REG_9_ & ~n37813;
  assign n37816 = ~n37814 & ~n37815;
  assign n37817 = n34683 & n37816;
  assign n37818 = n37796 & n37809;
  assign n37819 = ~n37817 & n37818;
  assign n37820 = n37762 & ~n37763;
  assign n37821 = ~n37777 & n37820;
  assign n37822 = n37789 & n37821;
  assign n37823 = n37819 & n37822;
  assign n37824 = n36647 & ~n37823;
  assign n37825 = ~n37744 & ~n37745;
  assign n6596 = n37824 | ~n37825;
  assign n37827 = P1_P2_INSTADDRPOINTER_REG_10_ & n36646;
  assign n37828 = P1_P2_REIP_REG_10_ & n36791;
  assign n37829 = P1_P2_INSTADDRPOINTER_REG_9_ & n37746;
  assign n37830 = ~P1_P2_INSTADDRPOINTER_REG_10_ & n37829;
  assign n37831 = P1_P2_INSTADDRPOINTER_REG_10_ & ~n37829;
  assign n37832 = ~n37830 & ~n37831;
  assign n37833 = n34840 & ~n37832;
  assign n37834 = n34841 & ~n37832;
  assign n37835 = P1_P2_INSTADDRPOINTER_REG_9_ & n37752;
  assign n37836 = ~P1_P2_INSTADDRPOINTER_REG_10_ & n37835;
  assign n37837 = P1_P2_INSTADDRPOINTER_REG_10_ & ~n37835;
  assign n37838 = ~n37836 & ~n37837;
  assign n37839 = n36655 & ~n37838;
  assign n37840 = n34656 & ~n37832;
  assign n37841 = n36658 & ~n37838;
  assign n37842 = ~n37840 & ~n37841;
  assign n37843 = ~n37833 & ~n37834;
  assign n37844 = ~n37839 & n37843;
  assign n37845 = n37842 & n37844;
  assign n37846 = ~n34769 & ~n37838;
  assign n37847 = ~n37764 & ~n37773;
  assign n37848 = ~n37677 & n37847;
  assign n37849 = ~n37766 & ~n37772;
  assign n37850 = ~n37848 & n37849;
  assign n37851 = ~P1_P2_INSTADDRPOINTER_REG_10_ & ~n37582;
  assign n37852 = P1_P2_INSTADDRPOINTER_REG_10_ & n37582;
  assign n37853 = ~n37851 & ~n37852;
  assign n37854 = n37850 & ~n37853;
  assign n37855 = P1_P2_INSTADDRPOINTER_REG_10_ & ~n37582;
  assign n37856 = ~P1_P2_INSTADDRPOINTER_REG_10_ & n37582;
  assign n37857 = ~n37855 & ~n37856;
  assign n37858 = ~n37850 & ~n37857;
  assign n37859 = ~n37854 & ~n37858;
  assign n37860 = n36752 & ~n37859;
  assign n37861 = n34879 & ~n37838;
  assign n37862 = n34722 & ~n37838;
  assign n37863 = ~n37861 & ~n37862;
  assign n37864 = ~P1_P2_INSTADDRPOINTER_REG_10_ & ~n37786;
  assign n37865 = P1_P2_INSTADDRPOINTER_REG_9_ & P1_P2_INSTADDRPOINTER_REG_10_;
  assign n37866 = ~n37784 & n37865;
  assign n37867 = ~n37864 & ~n37866;
  assign n37868 = n36754 & n37867;
  assign n37869 = n37863 & ~n37868;
  assign n37870 = n36771 & ~n37838;
  assign n37871 = n34726 & ~n37838;
  assign n37872 = n36760 & ~n37838;
  assign n37873 = n36764 & ~n37838;
  assign n37874 = ~n37870 & ~n37871;
  assign n37875 = ~n37872 & n37874;
  assign n37876 = ~n37873 & n37875;
  assign n37877 = n34582 & ~n37832;
  assign n37878 = n34660 & ~n37832;
  assign n37879 = n34664 & ~n37832;
  assign n37880 = P1_P2_INSTADDRPOINTER_REG_9_ & n37800;
  assign n37881 = ~P1_P2_INSTADDRPOINTER_REG_10_ & n37880;
  assign n37882 = P1_P2_INSTADDRPOINTER_REG_10_ & ~n37880;
  assign n37883 = ~n37881 & ~n37882;
  assign n37884 = n34680 & ~n37883;
  assign n37885 = n34672 & ~n37883;
  assign n37886 = ~n37877 & ~n37878;
  assign n37887 = ~n37879 & n37886;
  assign n37888 = ~n37884 & n37887;
  assign n37889 = ~n37885 & n37888;
  assign n37890 = ~P1_P2_INSTADDRPOINTER_REG_10_ & ~n37815;
  assign n37891 = ~n37813 & n37865;
  assign n37892 = ~n37890 & ~n37891;
  assign n37893 = n34683 & n37892;
  assign n37894 = n37876 & n37889;
  assign n37895 = ~n37893 & n37894;
  assign n37896 = n37845 & ~n37846;
  assign n37897 = ~n37860 & n37896;
  assign n37898 = n37869 & n37897;
  assign n37899 = n37895 & n37898;
  assign n37900 = n36647 & ~n37899;
  assign n37901 = ~n37827 & ~n37828;
  assign n6601 = n37900 | ~n37901;
  assign n37903 = P1_P2_INSTADDRPOINTER_REG_11_ & n36646;
  assign n37904 = P1_P2_REIP_REG_11_ & n36791;
  assign n37905 = ~n37903 & ~n37904;
  assign n37906 = P1_P2_INSTADDRPOINTER_REG_10_ & n37835;
  assign n37907 = ~P1_P2_INSTADDRPOINTER_REG_11_ & n37906;
  assign n37908 = P1_P2_INSTADDRPOINTER_REG_11_ & ~n37906;
  assign n37909 = ~n37907 & ~n37908;
  assign n37910 = n36771 & ~n37909;
  assign n37911 = n34726 & ~n37909;
  assign n37912 = n36760 & ~n37909;
  assign n37913 = n36764 & ~n37909;
  assign n37914 = ~n37910 & ~n37911;
  assign n37915 = ~n37912 & n37914;
  assign n37916 = ~n37913 & n37915;
  assign n37917 = P1_P2_INSTADDRPOINTER_REG_10_ & n37829;
  assign n37918 = ~P1_P2_INSTADDRPOINTER_REG_11_ & n37917;
  assign n37919 = P1_P2_INSTADDRPOINTER_REG_11_ & ~n37917;
  assign n37920 = ~n37918 & ~n37919;
  assign n37921 = n34582 & ~n37920;
  assign n37922 = n34660 & ~n37920;
  assign n37923 = n34664 & ~n37920;
  assign n37924 = P1_P2_INSTADDRPOINTER_REG_10_ & n37880;
  assign n37925 = ~P1_P2_INSTADDRPOINTER_REG_11_ & n37924;
  assign n37926 = P1_P2_INSTADDRPOINTER_REG_11_ & ~n37924;
  assign n37927 = ~n37925 & ~n37926;
  assign n37928 = n34680 & ~n37927;
  assign n37929 = n34672 & ~n37927;
  assign n37930 = ~n37921 & ~n37922;
  assign n37931 = ~n37923 & n37930;
  assign n37932 = ~n37928 & n37931;
  assign n37933 = ~n37929 & n37932;
  assign n37934 = P1_P2_INSTADDRPOINTER_REG_11_ & ~n37891;
  assign n37935 = ~P1_P2_INSTADDRPOINTER_REG_11_ & n37891;
  assign n37936 = ~n37934 & ~n37935;
  assign n37937 = n34683 & ~n37936;
  assign n37938 = n37916 & n37933;
  assign n37939 = ~n37937 & n37938;
  assign n37940 = n34879 & ~n37909;
  assign n37941 = n34722 & ~n37909;
  assign n37942 = ~n37940 & ~n37941;
  assign n37943 = ~n34769 & ~n37909;
  assign n37944 = n37849 & ~n37855;
  assign n37945 = n37847 & ~n37856;
  assign n37946 = ~n37677 & n37945;
  assign n37947 = n37944 & ~n37946;
  assign n37948 = ~P1_P2_INSTADDRPOINTER_REG_11_ & ~n37582;
  assign n37949 = P1_P2_INSTADDRPOINTER_REG_11_ & n37582;
  assign n37950 = ~n37948 & ~n37949;
  assign n37951 = n37947 & ~n37950;
  assign n37952 = ~n37947 & n37950;
  assign n37953 = ~n37951 & ~n37952;
  assign n37954 = n36752 & ~n37953;
  assign n37955 = n34840 & ~n37920;
  assign n37956 = n34841 & ~n37920;
  assign n37957 = n36655 & ~n37909;
  assign n37958 = n34656 & ~n37920;
  assign n37959 = n36658 & ~n37909;
  assign n37960 = ~n37958 & ~n37959;
  assign n37961 = ~n37955 & ~n37956;
  assign n37962 = ~n37957 & n37961;
  assign n37963 = n37960 & n37962;
  assign n37964 = P1_P2_INSTADDRPOINTER_REG_11_ & ~n37866;
  assign n37965 = ~P1_P2_INSTADDRPOINTER_REG_11_ & n37866;
  assign n37966 = ~n37964 & ~n37965;
  assign n37967 = n36754 & ~n37966;
  assign n37968 = n37942 & ~n37943;
  assign n37969 = ~n37954 & n37968;
  assign n37970 = n37963 & n37969;
  assign n37971 = ~n37967 & n37970;
  assign n37972 = n37939 & n37971;
  assign n37973 = n36647 & ~n37972;
  assign n6606 = ~n37905 | n37973;
  assign n37975 = P1_P2_INSTADDRPOINTER_REG_12_ & n36646;
  assign n37976 = P1_P2_REIP_REG_12_ & n36791;
  assign n37977 = P1_P2_INSTADDRPOINTER_REG_11_ & n37917;
  assign n37978 = ~P1_P2_INSTADDRPOINTER_REG_12_ & n37977;
  assign n37979 = P1_P2_INSTADDRPOINTER_REG_12_ & ~n37977;
  assign n37980 = ~n37978 & ~n37979;
  assign n37981 = n34840 & ~n37980;
  assign n37982 = n34841 & ~n37980;
  assign n37983 = P1_P2_INSTADDRPOINTER_REG_11_ & n37906;
  assign n37984 = ~P1_P2_INSTADDRPOINTER_REG_12_ & n37983;
  assign n37985 = P1_P2_INSTADDRPOINTER_REG_12_ & ~n37983;
  assign n37986 = ~n37984 & ~n37985;
  assign n37987 = n36655 & ~n37986;
  assign n37988 = n34656 & ~n37980;
  assign n37989 = n36658 & ~n37986;
  assign n37990 = ~n37988 & ~n37989;
  assign n37991 = ~n37981 & ~n37982;
  assign n37992 = ~n37987 & n37991;
  assign n37993 = n37990 & n37992;
  assign n37994 = ~n34769 & ~n37986;
  assign n37995 = ~P1_P2_INSTADDRPOINTER_REG_12_ & ~n37582;
  assign n37996 = P1_P2_INSTADDRPOINTER_REG_12_ & n37582;
  assign n37997 = ~n37995 & ~n37996;
  assign n37998 = P1_P2_INSTADDRPOINTER_REG_11_ & ~n37582;
  assign n37999 = ~P1_P2_INSTADDRPOINTER_REG_11_ & n37582;
  assign n38000 = ~n37947 & ~n37999;
  assign n38001 = ~n37998 & ~n38000;
  assign n38002 = ~n37997 & n38001;
  assign n38003 = ~P1_P2_INSTADDRPOINTER_REG_12_ & n37582;
  assign n38004 = P1_P2_INSTADDRPOINTER_REG_12_ & ~n37582;
  assign n38005 = ~n38003 & ~n38004;
  assign n38006 = ~n38001 & ~n38005;
  assign n38007 = ~n38002 & ~n38006;
  assign n38008 = n36752 & ~n38007;
  assign n38009 = n34879 & ~n37986;
  assign n38010 = n34722 & ~n37986;
  assign n38011 = ~n38009 & ~n38010;
  assign n38012 = P1_P2_INSTADDRPOINTER_REG_11_ & n37866;
  assign n38013 = ~P1_P2_INSTADDRPOINTER_REG_12_ & ~n38012;
  assign n38014 = P1_P2_INSTADDRPOINTER_REG_11_ & P1_P2_INSTADDRPOINTER_REG_12_;
  assign n38015 = n37866 & n38014;
  assign n38016 = ~n38013 & ~n38015;
  assign n38017 = n36754 & n38016;
  assign n38018 = n38011 & ~n38017;
  assign n38019 = n36771 & ~n37986;
  assign n38020 = n34726 & ~n37986;
  assign n38021 = n36760 & ~n37986;
  assign n38022 = n36764 & ~n37986;
  assign n38023 = ~n38019 & ~n38020;
  assign n38024 = ~n38021 & n38023;
  assign n38025 = ~n38022 & n38024;
  assign n38026 = n34582 & ~n37980;
  assign n38027 = n34660 & ~n37980;
  assign n38028 = n34664 & ~n37980;
  assign n38029 = P1_P2_INSTADDRPOINTER_REG_11_ & n37924;
  assign n38030 = ~P1_P2_INSTADDRPOINTER_REG_12_ & n38029;
  assign n38031 = P1_P2_INSTADDRPOINTER_REG_12_ & ~n38029;
  assign n38032 = ~n38030 & ~n38031;
  assign n38033 = n34680 & ~n38032;
  assign n38034 = n34672 & ~n38032;
  assign n38035 = ~n38026 & ~n38027;
  assign n38036 = ~n38028 & n38035;
  assign n38037 = ~n38033 & n38036;
  assign n38038 = ~n38034 & n38037;
  assign n38039 = P1_P2_INSTADDRPOINTER_REG_11_ & n37891;
  assign n38040 = ~P1_P2_INSTADDRPOINTER_REG_12_ & ~n38039;
  assign n38041 = n37891 & n38014;
  assign n38042 = ~n38040 & ~n38041;
  assign n38043 = n34683 & n38042;
  assign n38044 = n38025 & n38038;
  assign n38045 = ~n38043 & n38044;
  assign n38046 = n37993 & ~n37994;
  assign n38047 = ~n38008 & n38046;
  assign n38048 = n38018 & n38047;
  assign n38049 = n38045 & n38048;
  assign n38050 = n36647 & ~n38049;
  assign n38051 = ~n37975 & ~n37976;
  assign n6611 = n38050 | ~n38051;
  assign n38053 = P1_P2_INSTADDRPOINTER_REG_13_ & n36646;
  assign n38054 = P1_P2_REIP_REG_13_ & n36791;
  assign n38055 = P1_P2_INSTADDRPOINTER_REG_12_ & n37977;
  assign n38056 = ~P1_P2_INSTADDRPOINTER_REG_13_ & n38055;
  assign n38057 = P1_P2_INSTADDRPOINTER_REG_13_ & ~n38055;
  assign n38058 = ~n38056 & ~n38057;
  assign n38059 = n34840 & ~n38058;
  assign n38060 = n34841 & ~n38058;
  assign n38061 = P1_P2_INSTADDRPOINTER_REG_12_ & n37983;
  assign n38062 = ~P1_P2_INSTADDRPOINTER_REG_13_ & n38061;
  assign n38063 = P1_P2_INSTADDRPOINTER_REG_13_ & ~n38061;
  assign n38064 = ~n38062 & ~n38063;
  assign n38065 = n36655 & ~n38064;
  assign n38066 = n34656 & ~n38058;
  assign n38067 = n36658 & ~n38064;
  assign n38068 = ~n38066 & ~n38067;
  assign n38069 = ~n38059 & ~n38060;
  assign n38070 = ~n38065 & n38069;
  assign n38071 = n38068 & n38070;
  assign n38072 = ~n34769 & ~n38064;
  assign n38073 = P1_P2_INSTADDRPOINTER_REG_13_ & ~n37582;
  assign n38074 = P1_P2_INSTADDRPOINTER_REG_12_ & P1_P2_INSTADDRPOINTER_REG_13_;
  assign n38075 = n37582 & ~n38074;
  assign n38076 = ~n38073 & ~n38075;
  assign n38077 = n38001 & ~n38004;
  assign n38078 = n38076 & ~n38077;
  assign n38079 = ~P1_P2_INSTADDRPOINTER_REG_13_ & ~n37582;
  assign n38080 = P1_P2_INSTADDRPOINTER_REG_13_ & n37582;
  assign n38081 = ~n38079 & ~n38080;
  assign n38082 = ~n38004 & n38081;
  assign n38083 = ~n38001 & ~n38003;
  assign n38084 = n38082 & ~n38083;
  assign n38085 = ~n38078 & ~n38084;
  assign n38086 = n36752 & n38085;
  assign n38087 = n34879 & ~n38064;
  assign n38088 = n34722 & ~n38064;
  assign n38089 = ~n38087 & ~n38088;
  assign n38090 = ~P1_P2_INSTADDRPOINTER_REG_13_ & ~n38015;
  assign n38091 = P1_P2_INSTADDRPOINTER_REG_13_ & n38015;
  assign n38092 = ~n38090 & ~n38091;
  assign n38093 = n36754 & n38092;
  assign n38094 = n38089 & ~n38093;
  assign n38095 = n36771 & ~n38064;
  assign n38096 = n34726 & ~n38064;
  assign n38097 = n36760 & ~n38064;
  assign n38098 = n36764 & ~n38064;
  assign n38099 = ~n38095 & ~n38096;
  assign n38100 = ~n38097 & n38099;
  assign n38101 = ~n38098 & n38100;
  assign n38102 = n34582 & ~n38058;
  assign n38103 = n34660 & ~n38058;
  assign n38104 = n34664 & ~n38058;
  assign n38105 = P1_P2_INSTADDRPOINTER_REG_12_ & n38029;
  assign n38106 = ~P1_P2_INSTADDRPOINTER_REG_13_ & n38105;
  assign n38107 = P1_P2_INSTADDRPOINTER_REG_13_ & ~n38105;
  assign n38108 = ~n38106 & ~n38107;
  assign n38109 = n34680 & ~n38108;
  assign n38110 = n34672 & ~n38108;
  assign n38111 = ~n38102 & ~n38103;
  assign n38112 = ~n38104 & n38111;
  assign n38113 = ~n38109 & n38112;
  assign n38114 = ~n38110 & n38113;
  assign n38115 = ~P1_P2_INSTADDRPOINTER_REG_13_ & ~n38041;
  assign n38116 = P1_P2_INSTADDRPOINTER_REG_13_ & n38041;
  assign n38117 = ~n38115 & ~n38116;
  assign n38118 = n34683 & n38117;
  assign n38119 = n38101 & n38114;
  assign n38120 = ~n38118 & n38119;
  assign n38121 = n38071 & ~n38072;
  assign n38122 = ~n38086 & n38121;
  assign n38123 = n38094 & n38122;
  assign n38124 = n38120 & n38123;
  assign n38125 = n36647 & ~n38124;
  assign n38126 = ~n38053 & ~n38054;
  assign n6616 = n38125 | ~n38126;
  assign n38128 = P1_P2_INSTADDRPOINTER_REG_14_ & n36646;
  assign n38129 = P1_P2_REIP_REG_14_ & n36791;
  assign n38130 = ~n38128 & ~n38129;
  assign n38131 = P1_P2_INSTADDRPOINTER_REG_13_ & n38061;
  assign n38132 = ~P1_P2_INSTADDRPOINTER_REG_14_ & n38131;
  assign n38133 = P1_P2_INSTADDRPOINTER_REG_14_ & ~n38131;
  assign n38134 = ~n38132 & ~n38133;
  assign n38135 = n36771 & ~n38134;
  assign n38136 = n34726 & ~n38134;
  assign n38137 = n36760 & ~n38134;
  assign n38138 = n36764 & ~n38134;
  assign n38139 = ~n38135 & ~n38136;
  assign n38140 = ~n38137 & n38139;
  assign n38141 = ~n38138 & n38140;
  assign n38142 = P1_P2_INSTADDRPOINTER_REG_13_ & n38055;
  assign n38143 = ~P1_P2_INSTADDRPOINTER_REG_14_ & n38142;
  assign n38144 = P1_P2_INSTADDRPOINTER_REG_14_ & ~n38142;
  assign n38145 = ~n38143 & ~n38144;
  assign n38146 = n34582 & ~n38145;
  assign n38147 = n34660 & ~n38145;
  assign n38148 = n34664 & ~n38145;
  assign n38149 = P1_P2_INSTADDRPOINTER_REG_13_ & n38105;
  assign n38150 = ~P1_P2_INSTADDRPOINTER_REG_14_ & n38149;
  assign n38151 = P1_P2_INSTADDRPOINTER_REG_14_ & ~n38149;
  assign n38152 = ~n38150 & ~n38151;
  assign n38153 = n34680 & ~n38152;
  assign n38154 = n34672 & ~n38152;
  assign n38155 = ~n38146 & ~n38147;
  assign n38156 = ~n38148 & n38155;
  assign n38157 = ~n38153 & n38156;
  assign n38158 = ~n38154 & n38157;
  assign n38159 = ~P1_P2_INSTADDRPOINTER_REG_14_ & n38116;
  assign n38160 = P1_P2_INSTADDRPOINTER_REG_14_ & ~n38116;
  assign n38161 = ~n38159 & ~n38160;
  assign n38162 = n34683 & ~n38161;
  assign n38163 = n38141 & n38158;
  assign n38164 = ~n38162 & n38163;
  assign n38165 = n34879 & ~n38134;
  assign n38166 = n34722 & ~n38134;
  assign n38167 = ~n38165 & ~n38166;
  assign n38168 = ~n34769 & ~n38134;
  assign n38169 = n34840 & ~n38145;
  assign n38170 = n34841 & ~n38145;
  assign n38171 = n36655 & ~n38134;
  assign n38172 = n34656 & ~n38145;
  assign n38173 = n36658 & ~n38134;
  assign n38174 = ~n38172 & ~n38173;
  assign n38175 = ~n38169 & ~n38170;
  assign n38176 = ~n38171 & n38175;
  assign n38177 = n38174 & n38176;
  assign n38178 = ~n38004 & ~n38073;
  assign n38179 = ~n37998 & n38178;
  assign n38180 = ~n37999 & ~n38075;
  assign n38181 = ~n37947 & n38180;
  assign n38182 = n38179 & ~n38181;
  assign n38183 = ~P1_P2_INSTADDRPOINTER_REG_14_ & ~n37582;
  assign n38184 = P1_P2_INSTADDRPOINTER_REG_14_ & n37582;
  assign n38185 = ~n38183 & ~n38184;
  assign n38186 = n38182 & ~n38185;
  assign n38187 = ~n38182 & n38185;
  assign n38188 = ~n38186 & ~n38187;
  assign n38189 = n36752 & ~n38188;
  assign n38190 = ~P1_P2_INSTADDRPOINTER_REG_14_ & n38091;
  assign n38191 = P1_P2_INSTADDRPOINTER_REG_14_ & ~n38091;
  assign n38192 = ~n38190 & ~n38191;
  assign n38193 = n36754 & ~n38192;
  assign n38194 = n38167 & ~n38168;
  assign n38195 = n38177 & n38194;
  assign n38196 = ~n38189 & n38195;
  assign n38197 = ~n38193 & n38196;
  assign n38198 = n38164 & n38197;
  assign n38199 = n36647 & ~n38198;
  assign n6621 = ~n38130 | n38199;
  assign n38201 = P1_P2_INSTADDRPOINTER_REG_15_ & n36646;
  assign n38202 = P1_P2_REIP_REG_15_ & n36791;
  assign n38203 = ~n38201 & ~n38202;
  assign n38204 = P1_P2_INSTADDRPOINTER_REG_14_ & n38131;
  assign n38205 = ~P1_P2_INSTADDRPOINTER_REG_15_ & n38204;
  assign n38206 = P1_P2_INSTADDRPOINTER_REG_15_ & ~n38204;
  assign n38207 = ~n38205 & ~n38206;
  assign n38208 = n36771 & ~n38207;
  assign n38209 = n34726 & ~n38207;
  assign n38210 = n36760 & ~n38207;
  assign n38211 = n36764 & ~n38207;
  assign n38212 = ~n38208 & ~n38209;
  assign n38213 = ~n38210 & n38212;
  assign n38214 = ~n38211 & n38213;
  assign n38215 = P1_P2_INSTADDRPOINTER_REG_14_ & n38142;
  assign n38216 = ~P1_P2_INSTADDRPOINTER_REG_15_ & n38215;
  assign n38217 = P1_P2_INSTADDRPOINTER_REG_15_ & ~n38215;
  assign n38218 = ~n38216 & ~n38217;
  assign n38219 = n34582 & ~n38218;
  assign n38220 = n34660 & ~n38218;
  assign n38221 = n34664 & ~n38218;
  assign n38222 = P1_P2_INSTADDRPOINTER_REG_14_ & n38149;
  assign n38223 = ~P1_P2_INSTADDRPOINTER_REG_15_ & n38222;
  assign n38224 = P1_P2_INSTADDRPOINTER_REG_15_ & ~n38222;
  assign n38225 = ~n38223 & ~n38224;
  assign n38226 = n34680 & ~n38225;
  assign n38227 = n34672 & ~n38225;
  assign n38228 = ~n38219 & ~n38220;
  assign n38229 = ~n38221 & n38228;
  assign n38230 = ~n38226 & n38229;
  assign n38231 = ~n38227 & n38230;
  assign n38232 = P1_P2_INSTADDRPOINTER_REG_14_ & n38116;
  assign n38233 = ~P1_P2_INSTADDRPOINTER_REG_15_ & ~n38232;
  assign n38234 = P1_P2_INSTADDRPOINTER_REG_14_ & P1_P2_INSTADDRPOINTER_REG_15_;
  assign n38235 = P1_P2_INSTADDRPOINTER_REG_13_ & n38234;
  assign n38236 = n38041 & n38235;
  assign n38237 = ~n38233 & ~n38236;
  assign n38238 = n34683 & n38237;
  assign n38239 = n38214 & n38231;
  assign n38240 = ~n38238 & n38239;
  assign n38241 = n34879 & ~n38207;
  assign n38242 = n34722 & ~n38207;
  assign n38243 = ~n38241 & ~n38242;
  assign n38244 = ~n34769 & ~n38207;
  assign n38245 = n34840 & ~n38218;
  assign n38246 = n34841 & ~n38218;
  assign n38247 = n36655 & ~n38207;
  assign n38248 = n34656 & ~n38218;
  assign n38249 = n36658 & ~n38207;
  assign n38250 = ~n38248 & ~n38249;
  assign n38251 = ~n38245 & ~n38246;
  assign n38252 = ~n38247 & n38251;
  assign n38253 = n38250 & n38252;
  assign n38254 = P1_P2_INSTADDRPOINTER_REG_14_ & ~n37582;
  assign n38255 = n38179 & ~n38254;
  assign n38256 = ~P1_P2_INSTADDRPOINTER_REG_14_ & n37582;
  assign n38257 = n38180 & ~n38256;
  assign n38258 = ~n37947 & n38257;
  assign n38259 = n38255 & ~n38258;
  assign n38260 = ~P1_P2_INSTADDRPOINTER_REG_15_ & ~n37582;
  assign n38261 = P1_P2_INSTADDRPOINTER_REG_15_ & n37582;
  assign n38262 = ~n38260 & ~n38261;
  assign n38263 = n38259 & ~n38262;
  assign n38264 = ~n38259 & n38262;
  assign n38265 = ~n38263 & ~n38264;
  assign n38266 = n36752 & ~n38265;
  assign n38267 = P1_P2_INSTADDRPOINTER_REG_14_ & n38091;
  assign n38268 = ~P1_P2_INSTADDRPOINTER_REG_15_ & ~n38267;
  assign n38269 = n38015 & n38235;
  assign n38270 = ~n38268 & ~n38269;
  assign n38271 = n36754 & n38270;
  assign n38272 = n38243 & ~n38244;
  assign n38273 = n38253 & n38272;
  assign n38274 = ~n38266 & n38273;
  assign n38275 = ~n38271 & n38274;
  assign n38276 = n38240 & n38275;
  assign n38277 = n36647 & ~n38276;
  assign n6626 = ~n38203 | n38277;
  assign n38279 = P1_P2_INSTADDRPOINTER_REG_16_ & n36646;
  assign n38280 = P1_P2_REIP_REG_16_ & n36791;
  assign n38281 = ~n38279 & ~n38280;
  assign n38282 = P1_P2_INSTADDRPOINTER_REG_15_ & n38204;
  assign n38283 = ~P1_P2_INSTADDRPOINTER_REG_16_ & n38282;
  assign n38284 = P1_P2_INSTADDRPOINTER_REG_16_ & ~n38282;
  assign n38285 = ~n38283 & ~n38284;
  assign n38286 = n36771 & ~n38285;
  assign n38287 = n34726 & ~n38285;
  assign n38288 = n36760 & ~n38285;
  assign n38289 = n36764 & ~n38285;
  assign n38290 = ~n38286 & ~n38287;
  assign n38291 = ~n38288 & n38290;
  assign n38292 = ~n38289 & n38291;
  assign n38293 = P1_P2_INSTADDRPOINTER_REG_15_ & n38215;
  assign n38294 = ~P1_P2_INSTADDRPOINTER_REG_16_ & n38293;
  assign n38295 = P1_P2_INSTADDRPOINTER_REG_16_ & ~n38293;
  assign n38296 = ~n38294 & ~n38295;
  assign n38297 = n34582 & ~n38296;
  assign n38298 = n34660 & ~n38296;
  assign n38299 = n34664 & ~n38296;
  assign n38300 = P1_P2_INSTADDRPOINTER_REG_15_ & n38222;
  assign n38301 = ~P1_P2_INSTADDRPOINTER_REG_16_ & n38300;
  assign n38302 = P1_P2_INSTADDRPOINTER_REG_16_ & ~n38300;
  assign n38303 = ~n38301 & ~n38302;
  assign n38304 = n34680 & ~n38303;
  assign n38305 = n34672 & ~n38303;
  assign n38306 = ~n38297 & ~n38298;
  assign n38307 = ~n38299 & n38306;
  assign n38308 = ~n38304 & n38307;
  assign n38309 = ~n38305 & n38308;
  assign n38310 = ~P1_P2_INSTADDRPOINTER_REG_16_ & n38236;
  assign n38311 = P1_P2_INSTADDRPOINTER_REG_16_ & ~n38236;
  assign n38312 = ~n38310 & ~n38311;
  assign n38313 = n34683 & ~n38312;
  assign n38314 = n38292 & n38309;
  assign n38315 = ~n38313 & n38314;
  assign n38316 = n34879 & ~n38285;
  assign n38317 = n34722 & ~n38285;
  assign n38318 = ~n38316 & ~n38317;
  assign n38319 = ~n34769 & ~n38285;
  assign n38320 = P1_P2_INSTADDRPOINTER_REG_15_ & ~n37582;
  assign n38321 = ~P1_P2_INSTADDRPOINTER_REG_15_ & n37582;
  assign n38322 = ~n38259 & ~n38321;
  assign n38323 = ~n38320 & ~n38322;
  assign n38324 = ~P1_P2_INSTADDRPOINTER_REG_16_ & ~n37582;
  assign n38325 = P1_P2_INSTADDRPOINTER_REG_16_ & n37582;
  assign n38326 = ~n38324 & ~n38325;
  assign n38327 = n38323 & ~n38326;
  assign n38328 = ~n38323 & n38326;
  assign n38329 = ~n38327 & ~n38328;
  assign n38330 = n36752 & ~n38329;
  assign n38331 = n34840 & ~n38296;
  assign n38332 = n34841 & ~n38296;
  assign n38333 = n36655 & ~n38285;
  assign n38334 = n34656 & ~n38296;
  assign n38335 = n36658 & ~n38285;
  assign n38336 = ~n38334 & ~n38335;
  assign n38337 = ~n38331 & ~n38332;
  assign n38338 = ~n38333 & n38337;
  assign n38339 = n38336 & n38338;
  assign n38340 = ~P1_P2_INSTADDRPOINTER_REG_16_ & n38269;
  assign n38341 = P1_P2_INSTADDRPOINTER_REG_16_ & ~n38269;
  assign n38342 = ~n38340 & ~n38341;
  assign n38343 = n36754 & ~n38342;
  assign n38344 = n38318 & ~n38319;
  assign n38345 = ~n38330 & n38344;
  assign n38346 = n38339 & n38345;
  assign n38347 = ~n38343 & n38346;
  assign n38348 = n38315 & n38347;
  assign n38349 = n36647 & ~n38348;
  assign n6631 = ~n38281 | n38349;
  assign n38351 = P1_P2_INSTADDRPOINTER_REG_17_ & n36646;
  assign n38352 = P1_P2_REIP_REG_17_ & n36791;
  assign n38353 = P1_P2_INSTADDRPOINTER_REG_16_ & n38293;
  assign n38354 = ~P1_P2_INSTADDRPOINTER_REG_17_ & n38353;
  assign n38355 = P1_P2_INSTADDRPOINTER_REG_17_ & ~n38353;
  assign n38356 = ~n38354 & ~n38355;
  assign n38357 = n34840 & ~n38356;
  assign n38358 = n34841 & ~n38356;
  assign n38359 = P1_P2_INSTADDRPOINTER_REG_16_ & n38282;
  assign n38360 = ~P1_P2_INSTADDRPOINTER_REG_17_ & n38359;
  assign n38361 = P1_P2_INSTADDRPOINTER_REG_17_ & ~n38359;
  assign n38362 = ~n38360 & ~n38361;
  assign n38363 = n36655 & ~n38362;
  assign n38364 = n34656 & ~n38356;
  assign n38365 = n36658 & ~n38362;
  assign n38366 = ~n38364 & ~n38365;
  assign n38367 = ~n38357 & ~n38358;
  assign n38368 = ~n38363 & n38367;
  assign n38369 = n38366 & n38368;
  assign n38370 = ~n34769 & ~n38362;
  assign n38371 = P1_P2_INSTADDRPOINTER_REG_16_ & P1_P2_INSTADDRPOINTER_REG_17_;
  assign n38372 = ~n38323 & n38371;
  assign n38373 = n37582 & ~n38372;
  assign n38374 = P1_P2_INSTADDRPOINTER_REG_17_ & ~n37582;
  assign n38375 = ~P1_P2_INSTADDRPOINTER_REG_16_ & ~n38320;
  assign n38376 = ~n38322 & n38375;
  assign n38377 = ~n38373 & ~n38374;
  assign n38378 = ~n38376 & n38377;
  assign n38379 = P1_P2_INSTADDRPOINTER_REG_17_ & n38376;
  assign n38380 = ~n37582 & ~n38379;
  assign n38381 = P1_P2_INSTADDRPOINTER_REG_17_ & n37582;
  assign n38382 = P1_P2_INSTADDRPOINTER_REG_16_ & ~n38323;
  assign n38383 = ~n38380 & ~n38381;
  assign n38384 = ~n38382 & n38383;
  assign n38385 = ~n38378 & ~n38384;
  assign n38386 = n36752 & n38385;
  assign n38387 = n34879 & ~n38362;
  assign n38388 = n34722 & ~n38362;
  assign n38389 = ~n38387 & ~n38388;
  assign n38390 = P1_P2_INSTADDRPOINTER_REG_16_ & n38269;
  assign n38391 = ~P1_P2_INSTADDRPOINTER_REG_17_ & ~n38390;
  assign n38392 = n38269 & n38371;
  assign n38393 = ~n38391 & ~n38392;
  assign n38394 = n36754 & n38393;
  assign n38395 = n38389 & ~n38394;
  assign n38396 = n36771 & ~n38362;
  assign n38397 = n34726 & ~n38362;
  assign n38398 = n36760 & ~n38362;
  assign n38399 = n36764 & ~n38362;
  assign n38400 = ~n38396 & ~n38397;
  assign n38401 = ~n38398 & n38400;
  assign n38402 = ~n38399 & n38401;
  assign n38403 = n34582 & ~n38356;
  assign n38404 = n34660 & ~n38356;
  assign n38405 = n34664 & ~n38356;
  assign n38406 = P1_P2_INSTADDRPOINTER_REG_16_ & n38300;
  assign n38407 = ~P1_P2_INSTADDRPOINTER_REG_17_ & n38406;
  assign n38408 = P1_P2_INSTADDRPOINTER_REG_17_ & ~n38406;
  assign n38409 = ~n38407 & ~n38408;
  assign n38410 = n34680 & ~n38409;
  assign n38411 = n34672 & ~n38409;
  assign n38412 = ~n38403 & ~n38404;
  assign n38413 = ~n38405 & n38412;
  assign n38414 = ~n38410 & n38413;
  assign n38415 = ~n38411 & n38414;
  assign n38416 = P1_P2_INSTADDRPOINTER_REG_16_ & n38236;
  assign n38417 = ~P1_P2_INSTADDRPOINTER_REG_17_ & ~n38416;
  assign n38418 = n38236 & n38371;
  assign n38419 = ~n38417 & ~n38418;
  assign n38420 = n34683 & n38419;
  assign n38421 = n38402 & n38415;
  assign n38422 = ~n38420 & n38421;
  assign n38423 = n38369 & ~n38370;
  assign n38424 = ~n38386 & n38423;
  assign n38425 = n38395 & n38424;
  assign n38426 = n38422 & n38425;
  assign n38427 = n36647 & ~n38426;
  assign n38428 = ~n38351 & ~n38352;
  assign n6636 = n38427 | ~n38428;
  assign n38430 = P1_P2_INSTADDRPOINTER_REG_18_ & n36646;
  assign n38431 = P1_P2_REIP_REG_18_ & n36791;
  assign n38432 = ~n38430 & ~n38431;
  assign n38433 = P1_P2_INSTADDRPOINTER_REG_17_ & n38359;
  assign n38434 = ~P1_P2_INSTADDRPOINTER_REG_18_ & n38433;
  assign n38435 = P1_P2_INSTADDRPOINTER_REG_18_ & ~n38433;
  assign n38436 = ~n38434 & ~n38435;
  assign n38437 = n36771 & ~n38436;
  assign n38438 = n34726 & ~n38436;
  assign n38439 = n36760 & ~n38436;
  assign n38440 = n36764 & ~n38436;
  assign n38441 = ~n38437 & ~n38438;
  assign n38442 = ~n38439 & n38441;
  assign n38443 = ~n38440 & n38442;
  assign n38444 = P1_P2_INSTADDRPOINTER_REG_17_ & n38353;
  assign n38445 = ~P1_P2_INSTADDRPOINTER_REG_18_ & n38444;
  assign n38446 = P1_P2_INSTADDRPOINTER_REG_18_ & ~n38444;
  assign n38447 = ~n38445 & ~n38446;
  assign n38448 = n34582 & ~n38447;
  assign n38449 = n34660 & ~n38447;
  assign n38450 = n34664 & ~n38447;
  assign n38451 = P1_P2_INSTADDRPOINTER_REG_17_ & n38406;
  assign n38452 = ~P1_P2_INSTADDRPOINTER_REG_18_ & n38451;
  assign n38453 = P1_P2_INSTADDRPOINTER_REG_18_ & ~n38451;
  assign n38454 = ~n38452 & ~n38453;
  assign n38455 = n34680 & ~n38454;
  assign n38456 = n34672 & ~n38454;
  assign n38457 = ~n38448 & ~n38449;
  assign n38458 = ~n38450 & n38457;
  assign n38459 = ~n38455 & n38458;
  assign n38460 = ~n38456 & n38459;
  assign n38461 = ~P1_P2_INSTADDRPOINTER_REG_18_ & n38418;
  assign n38462 = P1_P2_INSTADDRPOINTER_REG_18_ & ~n38418;
  assign n38463 = ~n38461 & ~n38462;
  assign n38464 = n34683 & ~n38463;
  assign n38465 = n38443 & n38460;
  assign n38466 = ~n38464 & n38465;
  assign n38467 = n34879 & ~n38436;
  assign n38468 = n34722 & ~n38436;
  assign n38469 = ~n38467 & ~n38468;
  assign n38470 = ~n34769 & ~n38436;
  assign n38471 = ~n37582 & ~n38376;
  assign n38472 = ~n38372 & ~n38471;
  assign n38473 = ~n38374 & n38472;
  assign n38474 = ~P1_P2_INSTADDRPOINTER_REG_18_ & ~n37582;
  assign n38475 = P1_P2_INSTADDRPOINTER_REG_18_ & n37582;
  assign n38476 = ~n38474 & ~n38475;
  assign n38477 = n38473 & ~n38476;
  assign n38478 = ~n38473 & n38476;
  assign n38479 = ~n38477 & ~n38478;
  assign n38480 = n36752 & ~n38479;
  assign n38481 = n34840 & ~n38447;
  assign n38482 = n34841 & ~n38447;
  assign n38483 = n36655 & ~n38436;
  assign n38484 = n34656 & ~n38447;
  assign n38485 = n36658 & ~n38436;
  assign n38486 = ~n38484 & ~n38485;
  assign n38487 = ~n38481 & ~n38482;
  assign n38488 = ~n38483 & n38487;
  assign n38489 = n38486 & n38488;
  assign n38490 = ~P1_P2_INSTADDRPOINTER_REG_18_ & n38392;
  assign n38491 = P1_P2_INSTADDRPOINTER_REG_18_ & ~n38392;
  assign n38492 = ~n38490 & ~n38491;
  assign n38493 = n36754 & ~n38492;
  assign n38494 = n38469 & ~n38470;
  assign n38495 = ~n38480 & n38494;
  assign n38496 = n38489 & n38495;
  assign n38497 = ~n38493 & n38496;
  assign n38498 = n38466 & n38497;
  assign n38499 = n36647 & ~n38498;
  assign n6641 = ~n38432 | n38499;
  assign n38501 = P1_P2_INSTADDRPOINTER_REG_19_ & n36646;
  assign n38502 = P1_P2_REIP_REG_19_ & n36791;
  assign n38503 = P1_P2_INSTADDRPOINTER_REG_18_ & n38444;
  assign n38504 = ~P1_P2_INSTADDRPOINTER_REG_19_ & n38503;
  assign n38505 = P1_P2_INSTADDRPOINTER_REG_19_ & ~n38503;
  assign n38506 = ~n38504 & ~n38505;
  assign n38507 = n34840 & ~n38506;
  assign n38508 = n34841 & ~n38506;
  assign n38509 = P1_P2_INSTADDRPOINTER_REG_18_ & n38433;
  assign n38510 = ~P1_P2_INSTADDRPOINTER_REG_19_ & n38509;
  assign n38511 = P1_P2_INSTADDRPOINTER_REG_19_ & ~n38509;
  assign n38512 = ~n38510 & ~n38511;
  assign n38513 = n36655 & ~n38512;
  assign n38514 = n34656 & ~n38506;
  assign n38515 = n36658 & ~n38512;
  assign n38516 = ~n38514 & ~n38515;
  assign n38517 = ~n38507 & ~n38508;
  assign n38518 = ~n38513 & n38517;
  assign n38519 = n38516 & n38518;
  assign n38520 = ~n34769 & ~n38512;
  assign n38521 = ~P1_P2_INSTADDRPOINTER_REG_19_ & ~n37582;
  assign n38522 = P1_P2_INSTADDRPOINTER_REG_19_ & n37582;
  assign n38523 = ~n38521 & ~n38522;
  assign n38524 = ~P1_P2_INSTADDRPOINTER_REG_18_ & n37582;
  assign n38525 = ~n38473 & ~n38524;
  assign n38526 = P1_P2_INSTADDRPOINTER_REG_18_ & ~n37582;
  assign n38527 = ~n38525 & ~n38526;
  assign n38528 = ~n38523 & n38527;
  assign n38529 = ~P1_P2_INSTADDRPOINTER_REG_19_ & n37582;
  assign n38530 = P1_P2_INSTADDRPOINTER_REG_19_ & ~n37582;
  assign n38531 = ~n38529 & ~n38530;
  assign n38532 = ~n38527 & ~n38531;
  assign n38533 = ~n38528 & ~n38532;
  assign n38534 = n36752 & ~n38533;
  assign n38535 = n34879 & ~n38512;
  assign n38536 = n34722 & ~n38512;
  assign n38537 = ~n38535 & ~n38536;
  assign n38538 = P1_P2_INSTADDRPOINTER_REG_18_ & n38392;
  assign n38539 = ~P1_P2_INSTADDRPOINTER_REG_19_ & ~n38538;
  assign n38540 = P1_P2_INSTADDRPOINTER_REG_18_ & P1_P2_INSTADDRPOINTER_REG_19_;
  assign n38541 = n38392 & n38540;
  assign n38542 = ~n38539 & ~n38541;
  assign n38543 = n36754 & n38542;
  assign n38544 = n38537 & ~n38543;
  assign n38545 = n36771 & ~n38512;
  assign n38546 = n34726 & ~n38512;
  assign n38547 = n36760 & ~n38512;
  assign n38548 = n36764 & ~n38512;
  assign n38549 = ~n38545 & ~n38546;
  assign n38550 = ~n38547 & n38549;
  assign n38551 = ~n38548 & n38550;
  assign n38552 = n34582 & ~n38506;
  assign n38553 = n34660 & ~n38506;
  assign n38554 = n34664 & ~n38506;
  assign n38555 = P1_P2_INSTADDRPOINTER_REG_18_ & n38451;
  assign n38556 = ~P1_P2_INSTADDRPOINTER_REG_19_ & n38555;
  assign n38557 = P1_P2_INSTADDRPOINTER_REG_19_ & ~n38555;
  assign n38558 = ~n38556 & ~n38557;
  assign n38559 = n34680 & ~n38558;
  assign n38560 = n34672 & ~n38558;
  assign n38561 = ~n38552 & ~n38553;
  assign n38562 = ~n38554 & n38561;
  assign n38563 = ~n38559 & n38562;
  assign n38564 = ~n38560 & n38563;
  assign n38565 = P1_P2_INSTADDRPOINTER_REG_18_ & n38418;
  assign n38566 = ~P1_P2_INSTADDRPOINTER_REG_19_ & ~n38565;
  assign n38567 = n38418 & n38540;
  assign n38568 = ~n38566 & ~n38567;
  assign n38569 = n34683 & n38568;
  assign n38570 = n38551 & n38564;
  assign n38571 = ~n38569 & n38570;
  assign n38572 = n38519 & ~n38520;
  assign n38573 = ~n38534 & n38572;
  assign n38574 = n38544 & n38573;
  assign n38575 = n38571 & n38574;
  assign n38576 = n36647 & ~n38575;
  assign n38577 = ~n38501 & ~n38502;
  assign n6646 = n38576 | ~n38577;
  assign n38579 = P1_P2_INSTADDRPOINTER_REG_20_ & n36646;
  assign n38580 = P1_P2_REIP_REG_20_ & n36791;
  assign n38581 = ~n38579 & ~n38580;
  assign n38582 = P1_P2_INSTADDRPOINTER_REG_19_ & P1_P2_INSTADDRPOINTER_REG_20_;
  assign n38583 = n37582 & ~n38582;
  assign n38584 = P1_P2_INSTADDRPOINTER_REG_20_ & ~n37582;
  assign n38585 = ~n38583 & ~n38584;
  assign n38586 = n38527 & ~n38530;
  assign n38587 = n38585 & ~n38586;
  assign n38588 = ~P1_P2_INSTADDRPOINTER_REG_19_ & n38527;
  assign n38589 = P1_P2_INSTADDRPOINTER_REG_20_ & n38588;
  assign n38590 = ~n37582 & ~n38589;
  assign n38591 = P1_P2_INSTADDRPOINTER_REG_20_ & n37582;
  assign n38592 = P1_P2_INSTADDRPOINTER_REG_19_ & ~n38527;
  assign n38593 = ~n38590 & ~n38591;
  assign n38594 = ~n38592 & n38593;
  assign n38595 = ~n38587 & ~n38594;
  assign n38596 = n36752 & n38595;
  assign n38597 = P1_P2_INSTADDRPOINTER_REG_19_ & n38509;
  assign n38598 = ~P1_P2_INSTADDRPOINTER_REG_20_ & n38597;
  assign n38599 = P1_P2_INSTADDRPOINTER_REG_20_ & ~n38597;
  assign n38600 = ~n38598 & ~n38599;
  assign n38601 = ~n34769 & ~n38600;
  assign n38602 = n34879 & ~n38600;
  assign n38603 = n34722 & ~n38600;
  assign n38604 = ~n38602 & ~n38603;
  assign n38605 = P1_P2_INSTADDRPOINTER_REG_19_ & n38503;
  assign n38606 = ~P1_P2_INSTADDRPOINTER_REG_20_ & n38605;
  assign n38607 = P1_P2_INSTADDRPOINTER_REG_20_ & ~n38605;
  assign n38608 = ~n38606 & ~n38607;
  assign n38609 = n34840 & ~n38608;
  assign n38610 = n34841 & ~n38608;
  assign n38611 = n36655 & ~n38600;
  assign n38612 = n34656 & ~n38608;
  assign n38613 = n36658 & ~n38600;
  assign n38614 = ~n38612 & ~n38613;
  assign n38615 = ~n38609 & ~n38610;
  assign n38616 = ~n38611 & n38615;
  assign n38617 = n38614 & n38616;
  assign n38618 = ~P1_P2_INSTADDRPOINTER_REG_20_ & ~n38541;
  assign n38619 = P1_P2_INSTADDRPOINTER_REG_20_ & n38541;
  assign n38620 = ~n38618 & ~n38619;
  assign n38621 = n36754 & n38620;
  assign n38622 = n36771 & ~n38600;
  assign n38623 = n34726 & ~n38600;
  assign n38624 = n36760 & ~n38600;
  assign n38625 = n36764 & ~n38600;
  assign n38626 = ~n38622 & ~n38623;
  assign n38627 = ~n38624 & n38626;
  assign n38628 = ~n38625 & n38627;
  assign n38629 = n34582 & ~n38608;
  assign n38630 = n34660 & ~n38608;
  assign n38631 = n34664 & ~n38608;
  assign n38632 = P1_P2_INSTADDRPOINTER_REG_19_ & n38555;
  assign n38633 = ~P1_P2_INSTADDRPOINTER_REG_20_ & n38632;
  assign n38634 = P1_P2_INSTADDRPOINTER_REG_20_ & ~n38632;
  assign n38635 = ~n38633 & ~n38634;
  assign n38636 = n34680 & ~n38635;
  assign n38637 = n34672 & ~n38635;
  assign n38638 = ~n38629 & ~n38630;
  assign n38639 = ~n38631 & n38638;
  assign n38640 = ~n38636 & n38639;
  assign n38641 = ~n38637 & n38640;
  assign n38642 = ~P1_P2_INSTADDRPOINTER_REG_20_ & ~n38567;
  assign n38643 = P1_P2_INSTADDRPOINTER_REG_20_ & n38567;
  assign n38644 = ~n38642 & ~n38643;
  assign n38645 = n34683 & n38644;
  assign n38646 = n38628 & n38641;
  assign n38647 = ~n38645 & n38646;
  assign n38648 = ~n38601 & n38604;
  assign n38649 = n38617 & n38648;
  assign n38650 = ~n38621 & n38649;
  assign n38651 = n38647 & n38650;
  assign n38652 = ~n38596 & n38651;
  assign n38653 = n36647 & ~n38652;
  assign n6651 = ~n38581 | n38653;
  assign n38655 = P1_P2_INSTADDRPOINTER_REG_21_ & n36646;
  assign n38656 = P1_P2_REIP_REG_21_ & n36791;
  assign n38657 = P1_P2_INSTADDRPOINTER_REG_20_ & n38597;
  assign n38658 = ~P1_P2_INSTADDRPOINTER_REG_21_ & n38657;
  assign n38659 = P1_P2_INSTADDRPOINTER_REG_21_ & ~n38657;
  assign n38660 = ~n38658 & ~n38659;
  assign n38661 = ~n34769 & ~n38660;
  assign n38662 = P1_P2_INSTADDRPOINTER_REG_20_ & n38605;
  assign n38663 = ~P1_P2_INSTADDRPOINTER_REG_21_ & n38662;
  assign n38664 = P1_P2_INSTADDRPOINTER_REG_21_ & ~n38662;
  assign n38665 = ~n38663 & ~n38664;
  assign n38666 = n34840 & ~n38665;
  assign n38667 = n34841 & ~n38665;
  assign n38668 = n36655 & ~n38660;
  assign n38669 = n34656 & ~n38665;
  assign n38670 = n36658 & ~n38660;
  assign n38671 = ~n38669 & ~n38670;
  assign n38672 = ~n38666 & ~n38667;
  assign n38673 = ~n38668 & n38672;
  assign n38674 = n38671 & n38673;
  assign n38675 = ~P1_P2_INSTADDRPOINTER_REG_21_ & ~n38619;
  assign n38676 = P1_P2_INSTADDRPOINTER_REG_21_ & n38619;
  assign n38677 = ~n38675 & ~n38676;
  assign n38678 = n36754 & n38677;
  assign n38679 = n34582 & ~n38665;
  assign n38680 = n34660 & ~n38665;
  assign n38681 = n34664 & ~n38665;
  assign n38682 = P1_P2_INSTADDRPOINTER_REG_20_ & n38632;
  assign n38683 = ~P1_P2_INSTADDRPOINTER_REG_21_ & n38682;
  assign n38684 = P1_P2_INSTADDRPOINTER_REG_21_ & ~n38682;
  assign n38685 = ~n38683 & ~n38684;
  assign n38686 = n34680 & ~n38685;
  assign n38687 = n34672 & ~n38685;
  assign n38688 = ~n38679 & ~n38680;
  assign n38689 = ~n38681 & n38688;
  assign n38690 = ~n38686 & n38689;
  assign n38691 = ~n38687 & n38690;
  assign n38692 = n36771 & ~n38660;
  assign n38693 = n34726 & ~n38660;
  assign n38694 = n36760 & ~n38660;
  assign n38695 = n36764 & ~n38660;
  assign n38696 = ~n38692 & ~n38693;
  assign n38697 = ~n38694 & n38696;
  assign n38698 = ~n38695 & n38697;
  assign n38699 = ~P1_P2_INSTADDRPOINTER_REG_21_ & ~n38643;
  assign n38700 = P1_P2_INSTADDRPOINTER_REG_20_ & P1_P2_INSTADDRPOINTER_REG_21_;
  assign n38701 = n38567 & n38700;
  assign n38702 = ~n38699 & ~n38701;
  assign n38703 = n34683 & n38702;
  assign n38704 = n38691 & n38698;
  assign n38705 = ~n38703 & n38704;
  assign n38706 = n34879 & ~n38660;
  assign n38707 = n34722 & ~n38660;
  assign n38708 = ~n38706 & ~n38707;
  assign n38709 = ~n38527 & n38582;
  assign n38710 = ~n38584 & ~n38709;
  assign n38711 = ~n37582 & ~n38588;
  assign n38712 = n38710 & ~n38711;
  assign n38713 = ~P1_P2_INSTADDRPOINTER_REG_21_ & ~n37582;
  assign n38714 = P1_P2_INSTADDRPOINTER_REG_21_ & n37582;
  assign n38715 = ~n38713 & ~n38714;
  assign n38716 = n38712 & ~n38715;
  assign n38717 = ~n38712 & n38715;
  assign n38718 = ~n38716 & ~n38717;
  assign n38719 = n36752 & ~n38718;
  assign n38720 = n38708 & ~n38719;
  assign n38721 = ~n38661 & n38674;
  assign n38722 = ~n38678 & n38721;
  assign n38723 = n38705 & n38722;
  assign n38724 = n38720 & n38723;
  assign n38725 = n36647 & ~n38724;
  assign n38726 = ~n38655 & ~n38656;
  assign n6656 = n38725 | ~n38726;
  assign n38728 = P1_P2_INSTADDRPOINTER_REG_22_ & n36646;
  assign n38729 = P1_P2_REIP_REG_22_ & n36791;
  assign n38730 = ~n38728 & ~n38729;
  assign n38731 = P1_P2_INSTADDRPOINTER_REG_21_ & n38682;
  assign n38732 = ~P1_P2_INSTADDRPOINTER_REG_22_ & n38731;
  assign n38733 = P1_P2_INSTADDRPOINTER_REG_22_ & ~n38731;
  assign n38734 = ~n38732 & ~n38733;
  assign n38735 = n34680 & ~n38734;
  assign n38736 = n34672 & ~n38734;
  assign n38737 = ~n38735 & ~n38736;
  assign n38738 = P1_P2_INSTADDRPOINTER_REG_21_ & n38662;
  assign n38739 = ~P1_P2_INSTADDRPOINTER_REG_22_ & n38738;
  assign n38740 = P1_P2_INSTADDRPOINTER_REG_22_ & ~n38738;
  assign n38741 = ~n38739 & ~n38740;
  assign n38742 = n34582 & ~n38741;
  assign n38743 = n34660 & ~n38741;
  assign n38744 = n34664 & ~n38741;
  assign n38745 = ~n38742 & ~n38743;
  assign n38746 = ~n38744 & n38745;
  assign n38747 = P1_P2_INSTADDRPOINTER_REG_21_ & n38657;
  assign n38748 = ~P1_P2_INSTADDRPOINTER_REG_22_ & n38747;
  assign n38749 = P1_P2_INSTADDRPOINTER_REG_22_ & ~n38747;
  assign n38750 = ~n38748 & ~n38749;
  assign n38751 = n36760 & ~n38750;
  assign n38752 = n36764 & ~n38750;
  assign n38753 = n34726 & ~n38750;
  assign n38754 = ~n38751 & ~n38752;
  assign n38755 = ~n38753 & n38754;
  assign n38756 = ~P1_P2_INSTADDRPOINTER_REG_22_ & n38701;
  assign n38757 = P1_P2_INSTADDRPOINTER_REG_22_ & ~n38701;
  assign n38758 = ~n38756 & ~n38757;
  assign n38759 = n34683 & ~n38758;
  assign n38760 = n36771 & ~n38750;
  assign n38761 = ~n38759 & ~n38760;
  assign n38762 = n38737 & n38746;
  assign n38763 = n38755 & n38762;
  assign n38764 = n38761 & n38763;
  assign n38765 = P1_P2_INSTADDRPOINTER_REG_21_ & n38582;
  assign n38766 = n37582 & ~n38765;
  assign n38767 = ~n38524 & ~n38766;
  assign n38768 = ~n38473 & n38767;
  assign n38769 = P1_P2_INSTADDRPOINTER_REG_21_ & ~n37582;
  assign n38770 = ~n38526 & ~n38769;
  assign n38771 = ~n38530 & n38770;
  assign n38772 = ~n38584 & n38771;
  assign n38773 = ~n38768 & n38772;
  assign n38774 = ~P1_P2_INSTADDRPOINTER_REG_22_ & ~n37582;
  assign n38775 = P1_P2_INSTADDRPOINTER_REG_22_ & n37582;
  assign n38776 = ~n38774 & ~n38775;
  assign n38777 = n38773 & ~n38776;
  assign n38778 = ~n38773 & n38776;
  assign n38779 = ~n38777 & ~n38778;
  assign n38780 = n36752 & ~n38779;
  assign n38781 = ~n34769 & ~n38750;
  assign n38782 = n34879 & ~n38750;
  assign n38783 = n34722 & ~n38750;
  assign n38784 = ~n38782 & ~n38783;
  assign n38785 = n34840 & ~n38741;
  assign n38786 = n34841 & ~n38741;
  assign n38787 = n36655 & ~n38750;
  assign n38788 = n34656 & ~n38741;
  assign n38789 = n36658 & ~n38750;
  assign n38790 = ~n38788 & ~n38789;
  assign n38791 = ~n38785 & ~n38786;
  assign n38792 = ~n38787 & n38791;
  assign n38793 = n38790 & n38792;
  assign n38794 = ~P1_P2_INSTADDRPOINTER_REG_22_ & n38676;
  assign n38795 = P1_P2_INSTADDRPOINTER_REG_22_ & ~n38676;
  assign n38796 = ~n38794 & ~n38795;
  assign n38797 = n36754 & ~n38796;
  assign n38798 = ~n38780 & ~n38781;
  assign n38799 = n38784 & n38798;
  assign n38800 = n38793 & n38799;
  assign n38801 = ~n38797 & n38800;
  assign n38802 = n38764 & n38801;
  assign n38803 = n36647 & ~n38802;
  assign n6661 = ~n38730 | n38803;
  assign n38805 = P1_P2_INSTADDRPOINTER_REG_23_ & n36646;
  assign n38806 = P1_P2_REIP_REG_23_ & n36791;
  assign n38807 = ~n38805 & ~n38806;
  assign n38808 = P1_P2_INSTADDRPOINTER_REG_22_ & n38731;
  assign n38809 = ~P1_P2_INSTADDRPOINTER_REG_23_ & n38808;
  assign n38810 = P1_P2_INSTADDRPOINTER_REG_23_ & ~n38808;
  assign n38811 = ~n38809 & ~n38810;
  assign n38812 = n34680 & ~n38811;
  assign n38813 = n34672 & ~n38811;
  assign n38814 = ~n38812 & ~n38813;
  assign n38815 = P1_P2_INSTADDRPOINTER_REG_22_ & n38738;
  assign n38816 = ~P1_P2_INSTADDRPOINTER_REG_23_ & n38815;
  assign n38817 = P1_P2_INSTADDRPOINTER_REG_23_ & ~n38815;
  assign n38818 = ~n38816 & ~n38817;
  assign n38819 = n34582 & ~n38818;
  assign n38820 = n34660 & ~n38818;
  assign n38821 = n34664 & ~n38818;
  assign n38822 = ~n38819 & ~n38820;
  assign n38823 = ~n38821 & n38822;
  assign n38824 = P1_P2_INSTADDRPOINTER_REG_22_ & n38747;
  assign n38825 = ~P1_P2_INSTADDRPOINTER_REG_23_ & n38824;
  assign n38826 = P1_P2_INSTADDRPOINTER_REG_23_ & ~n38824;
  assign n38827 = ~n38825 & ~n38826;
  assign n38828 = n36760 & ~n38827;
  assign n38829 = n36764 & ~n38827;
  assign n38830 = n34726 & ~n38827;
  assign n38831 = ~n38828 & ~n38829;
  assign n38832 = ~n38830 & n38831;
  assign n38833 = P1_P2_INSTADDRPOINTER_REG_22_ & n38701;
  assign n38834 = ~P1_P2_INSTADDRPOINTER_REG_23_ & ~n38833;
  assign n38835 = P1_P2_INSTADDRPOINTER_REG_22_ & P1_P2_INSTADDRPOINTER_REG_23_;
  assign n38836 = n38701 & n38835;
  assign n38837 = ~n38834 & ~n38836;
  assign n38838 = n34683 & n38837;
  assign n38839 = n36771 & ~n38827;
  assign n38840 = ~n38838 & ~n38839;
  assign n38841 = n38814 & n38823;
  assign n38842 = n38832 & n38841;
  assign n38843 = n38840 & n38842;
  assign n38844 = ~P1_P2_INSTADDRPOINTER_REG_22_ & n37582;
  assign n38845 = n38767 & ~n38844;
  assign n38846 = ~n38473 & n38845;
  assign n38847 = P1_P2_INSTADDRPOINTER_REG_22_ & ~n37582;
  assign n38848 = n38772 & ~n38847;
  assign n38849 = ~n38846 & n38848;
  assign n38850 = ~P1_P2_INSTADDRPOINTER_REG_23_ & ~n37582;
  assign n38851 = P1_P2_INSTADDRPOINTER_REG_23_ & n37582;
  assign n38852 = ~n38850 & ~n38851;
  assign n38853 = n38849 & ~n38852;
  assign n38854 = ~n38849 & n38852;
  assign n38855 = ~n38853 & ~n38854;
  assign n38856 = n36752 & ~n38855;
  assign n38857 = ~n34769 & ~n38827;
  assign n38858 = n34879 & ~n38827;
  assign n38859 = n34722 & ~n38827;
  assign n38860 = ~n38858 & ~n38859;
  assign n38861 = n34840 & ~n38818;
  assign n38862 = n34841 & ~n38818;
  assign n38863 = n36655 & ~n38827;
  assign n38864 = n34656 & ~n38818;
  assign n38865 = n36658 & ~n38827;
  assign n38866 = ~n38864 & ~n38865;
  assign n38867 = ~n38861 & ~n38862;
  assign n38868 = ~n38863 & n38867;
  assign n38869 = n38866 & n38868;
  assign n38870 = P1_P2_INSTADDRPOINTER_REG_22_ & n38676;
  assign n38871 = ~P1_P2_INSTADDRPOINTER_REG_23_ & ~n38870;
  assign n38872 = n38676 & n38835;
  assign n38873 = ~n38871 & ~n38872;
  assign n38874 = n36754 & n38873;
  assign n38875 = ~n38856 & ~n38857;
  assign n38876 = n38860 & n38875;
  assign n38877 = n38869 & n38876;
  assign n38878 = ~n38874 & n38877;
  assign n38879 = n38843 & n38878;
  assign n38880 = n36647 & ~n38879;
  assign n6666 = ~n38807 | n38880;
  assign n38882 = P1_P2_INSTADDRPOINTER_REG_24_ & n36646;
  assign n38883 = P1_P2_REIP_REG_24_ & n36791;
  assign n38884 = ~n38882 & ~n38883;
  assign n38885 = P1_P2_INSTADDRPOINTER_REG_23_ & n38808;
  assign n38886 = ~P1_P2_INSTADDRPOINTER_REG_24_ & n38885;
  assign n38887 = P1_P2_INSTADDRPOINTER_REG_24_ & ~n38885;
  assign n38888 = ~n38886 & ~n38887;
  assign n38889 = n34680 & ~n38888;
  assign n38890 = n34672 & ~n38888;
  assign n38891 = ~n38889 & ~n38890;
  assign n38892 = P1_P2_INSTADDRPOINTER_REG_23_ & n38815;
  assign n38893 = ~P1_P2_INSTADDRPOINTER_REG_24_ & n38892;
  assign n38894 = P1_P2_INSTADDRPOINTER_REG_24_ & ~n38892;
  assign n38895 = ~n38893 & ~n38894;
  assign n38896 = n34582 & ~n38895;
  assign n38897 = n34660 & ~n38895;
  assign n38898 = n34664 & ~n38895;
  assign n38899 = ~n38896 & ~n38897;
  assign n38900 = ~n38898 & n38899;
  assign n38901 = ~P1_P2_INSTADDRPOINTER_REG_24_ & n38836;
  assign n38902 = P1_P2_INSTADDRPOINTER_REG_24_ & ~n38836;
  assign n38903 = ~n38901 & ~n38902;
  assign n38904 = n34683 & ~n38903;
  assign n38905 = P1_P2_INSTADDRPOINTER_REG_23_ & n38824;
  assign n38906 = ~P1_P2_INSTADDRPOINTER_REG_24_ & n38905;
  assign n38907 = P1_P2_INSTADDRPOINTER_REG_24_ & ~n38905;
  assign n38908 = ~n38906 & ~n38907;
  assign n38909 = n36771 & ~n38908;
  assign n38910 = ~n38904 & ~n38909;
  assign n38911 = n36760 & ~n38908;
  assign n38912 = n36764 & ~n38908;
  assign n38913 = n34726 & ~n38908;
  assign n38914 = ~n38911 & ~n38912;
  assign n38915 = ~n38913 & n38914;
  assign n38916 = n38891 & n38900;
  assign n38917 = n38910 & n38916;
  assign n38918 = n38915 & n38917;
  assign n38919 = P1_P2_INSTADDRPOINTER_REG_23_ & ~n37582;
  assign n38920 = n38848 & ~n38919;
  assign n38921 = ~P1_P2_INSTADDRPOINTER_REG_23_ & n37582;
  assign n38922 = n38845 & ~n38921;
  assign n38923 = ~n38473 & n38922;
  assign n38924 = n38920 & ~n38923;
  assign n38925 = ~P1_P2_INSTADDRPOINTER_REG_24_ & ~n37582;
  assign n38926 = P1_P2_INSTADDRPOINTER_REG_24_ & n37582;
  assign n38927 = ~n38925 & ~n38926;
  assign n38928 = n38924 & ~n38927;
  assign n38929 = ~n38924 & n38927;
  assign n38930 = ~n38928 & ~n38929;
  assign n38931 = n36752 & ~n38930;
  assign n38932 = ~n34769 & ~n38908;
  assign n38933 = n34879 & ~n38908;
  assign n38934 = n34722 & ~n38908;
  assign n38935 = ~n38933 & ~n38934;
  assign n38936 = ~P1_P2_INSTADDRPOINTER_REG_24_ & n38872;
  assign n38937 = P1_P2_INSTADDRPOINTER_REG_24_ & ~n38872;
  assign n38938 = ~n38936 & ~n38937;
  assign n38939 = n36754 & ~n38938;
  assign n38940 = n34840 & ~n38895;
  assign n38941 = n34841 & ~n38895;
  assign n38942 = n36655 & ~n38908;
  assign n38943 = n34656 & ~n38895;
  assign n38944 = n36658 & ~n38908;
  assign n38945 = ~n38943 & ~n38944;
  assign n38946 = ~n38940 & ~n38941;
  assign n38947 = ~n38942 & n38946;
  assign n38948 = n38945 & n38947;
  assign n38949 = ~n38931 & ~n38932;
  assign n38950 = n38935 & n38949;
  assign n38951 = ~n38939 & n38950;
  assign n38952 = n38948 & n38951;
  assign n38953 = n38918 & n38952;
  assign n38954 = n36647 & ~n38953;
  assign n6671 = ~n38884 | n38954;
  assign n38956 = P1_P2_INSTADDRPOINTER_REG_25_ & n36646;
  assign n38957 = P1_P2_REIP_REG_25_ & n36791;
  assign n38958 = ~n38956 & ~n38957;
  assign n38959 = P1_P2_INSTADDRPOINTER_REG_24_ & n38885;
  assign n38960 = ~P1_P2_INSTADDRPOINTER_REG_25_ & n38959;
  assign n38961 = P1_P2_INSTADDRPOINTER_REG_25_ & ~n38959;
  assign n38962 = ~n38960 & ~n38961;
  assign n38963 = n34680 & ~n38962;
  assign n38964 = n34672 & ~n38962;
  assign n38965 = ~n38963 & ~n38964;
  assign n38966 = P1_P2_INSTADDRPOINTER_REG_24_ & n38892;
  assign n38967 = ~P1_P2_INSTADDRPOINTER_REG_25_ & n38966;
  assign n38968 = P1_P2_INSTADDRPOINTER_REG_25_ & ~n38966;
  assign n38969 = ~n38967 & ~n38968;
  assign n38970 = n34582 & ~n38969;
  assign n38971 = n34660 & ~n38969;
  assign n38972 = n34664 & ~n38969;
  assign n38973 = ~n38970 & ~n38971;
  assign n38974 = ~n38972 & n38973;
  assign n38975 = P1_P2_INSTADDRPOINTER_REG_24_ & n38836;
  assign n38976 = ~P1_P2_INSTADDRPOINTER_REG_25_ & ~n38975;
  assign n38977 = P1_P2_INSTADDRPOINTER_REG_24_ & P1_P2_INSTADDRPOINTER_REG_25_;
  assign n38978 = n38836 & n38977;
  assign n38979 = ~n38976 & ~n38978;
  assign n38980 = n34683 & n38979;
  assign n38981 = P1_P2_INSTADDRPOINTER_REG_24_ & n38905;
  assign n38982 = ~P1_P2_INSTADDRPOINTER_REG_25_ & n38981;
  assign n38983 = P1_P2_INSTADDRPOINTER_REG_25_ & ~n38981;
  assign n38984 = ~n38982 & ~n38983;
  assign n38985 = n36771 & ~n38984;
  assign n38986 = ~n38980 & ~n38985;
  assign n38987 = n36760 & ~n38984;
  assign n38988 = n36764 & ~n38984;
  assign n38989 = n34726 & ~n38984;
  assign n38990 = ~n38987 & ~n38988;
  assign n38991 = ~n38989 & n38990;
  assign n38992 = n38965 & n38974;
  assign n38993 = n38986 & n38992;
  assign n38994 = n38991 & n38993;
  assign n38995 = ~P1_P2_INSTADDRPOINTER_REG_25_ & ~n37582;
  assign n38996 = P1_P2_INSTADDRPOINTER_REG_25_ & n37582;
  assign n38997 = ~n38995 & ~n38996;
  assign n38998 = P1_P2_INSTADDRPOINTER_REG_24_ & ~n37582;
  assign n38999 = ~P1_P2_INSTADDRPOINTER_REG_24_ & n37582;
  assign n39000 = ~n38924 & ~n38999;
  assign n39001 = ~n38998 & ~n39000;
  assign n39002 = ~n38997 & n39001;
  assign n39003 = ~P1_P2_INSTADDRPOINTER_REG_25_ & n37582;
  assign n39004 = P1_P2_INSTADDRPOINTER_REG_25_ & ~n37582;
  assign n39005 = ~n39003 & ~n39004;
  assign n39006 = ~n39001 & ~n39005;
  assign n39007 = ~n39002 & ~n39006;
  assign n39008 = n36752 & ~n39007;
  assign n39009 = ~n34769 & ~n38984;
  assign n39010 = P1_P2_INSTADDRPOINTER_REG_24_ & n38872;
  assign n39011 = ~P1_P2_INSTADDRPOINTER_REG_25_ & ~n39010;
  assign n39012 = n38872 & n38977;
  assign n39013 = ~n39011 & ~n39012;
  assign n39014 = n36754 & n39013;
  assign n39015 = n34879 & ~n38984;
  assign n39016 = n34722 & ~n38984;
  assign n39017 = ~n39015 & ~n39016;
  assign n39018 = n34840 & ~n38969;
  assign n39019 = n34841 & ~n38969;
  assign n39020 = n36655 & ~n38984;
  assign n39021 = n34656 & ~n38969;
  assign n39022 = n36658 & ~n38984;
  assign n39023 = ~n39021 & ~n39022;
  assign n39024 = ~n39018 & ~n39019;
  assign n39025 = ~n39020 & n39024;
  assign n39026 = n39023 & n39025;
  assign n39027 = ~n39008 & ~n39009;
  assign n39028 = ~n39014 & n39027;
  assign n39029 = n39017 & n39028;
  assign n39030 = n39026 & n39029;
  assign n39031 = n38994 & n39030;
  assign n39032 = n36647 & ~n39031;
  assign n6676 = ~n38958 | n39032;
  assign n39034 = P1_P2_INSTADDRPOINTER_REG_26_ & n36646;
  assign n39035 = P1_P2_REIP_REG_26_ & n36791;
  assign n39036 = P1_P2_INSTADDRPOINTER_REG_26_ & ~n37582;
  assign n39037 = P1_P2_INSTADDRPOINTER_REG_25_ & P1_P2_INSTADDRPOINTER_REG_26_;
  assign n39038 = n37582 & ~n39037;
  assign n39039 = ~n39036 & ~n39038;
  assign n39040 = n39001 & ~n39004;
  assign n39041 = n39039 & ~n39040;
  assign n39042 = ~P1_P2_INSTADDRPOINTER_REG_26_ & ~n37582;
  assign n39043 = P1_P2_INSTADDRPOINTER_REG_26_ & n37582;
  assign n39044 = ~n39042 & ~n39043;
  assign n39045 = ~n39004 & n39044;
  assign n39046 = ~n39001 & ~n39003;
  assign n39047 = n39045 & ~n39046;
  assign n39048 = ~n39041 & ~n39047;
  assign n39049 = n36752 & n39048;
  assign n39050 = ~P1_P2_INSTADDRPOINTER_REG_26_ & ~n39012;
  assign n39051 = P1_P2_INSTADDRPOINTER_REG_26_ & n39012;
  assign n39052 = ~n39050 & ~n39051;
  assign n39053 = n36754 & n39052;
  assign n39054 = ~n39049 & ~n39053;
  assign n39055 = P1_P2_INSTADDRPOINTER_REG_25_ & n38981;
  assign n39056 = ~P1_P2_INSTADDRPOINTER_REG_26_ & n39055;
  assign n39057 = P1_P2_INSTADDRPOINTER_REG_26_ & ~n39055;
  assign n39058 = ~n39056 & ~n39057;
  assign n39059 = ~n34769 & ~n39058;
  assign n39060 = n34879 & ~n39058;
  assign n39061 = n34722 & ~n39058;
  assign n39062 = ~n39060 & ~n39061;
  assign n39063 = P1_P2_INSTADDRPOINTER_REG_25_ & n38966;
  assign n39064 = ~P1_P2_INSTADDRPOINTER_REG_26_ & n39063;
  assign n39065 = P1_P2_INSTADDRPOINTER_REG_26_ & ~n39063;
  assign n39066 = ~n39064 & ~n39065;
  assign n39067 = n34840 & ~n39066;
  assign n39068 = n34841 & ~n39066;
  assign n39069 = n36655 & ~n39058;
  assign n39070 = n34656 & ~n39066;
  assign n39071 = n36658 & ~n39058;
  assign n39072 = ~n39070 & ~n39071;
  assign n39073 = ~n39067 & ~n39068;
  assign n39074 = ~n39069 & n39073;
  assign n39075 = n39072 & n39074;
  assign n39076 = P1_P2_INSTADDRPOINTER_REG_25_ & n38959;
  assign n39077 = ~P1_P2_INSTADDRPOINTER_REG_26_ & n39076;
  assign n39078 = P1_P2_INSTADDRPOINTER_REG_26_ & ~n39076;
  assign n39079 = ~n39077 & ~n39078;
  assign n39080 = n34680 & ~n39079;
  assign n39081 = n34672 & ~n39079;
  assign n39082 = ~n39080 & ~n39081;
  assign n39083 = n34582 & ~n39066;
  assign n39084 = n34660 & ~n39066;
  assign n39085 = n34664 & ~n39066;
  assign n39086 = ~n39083 & ~n39084;
  assign n39087 = ~n39085 & n39086;
  assign n39088 = ~P1_P2_INSTADDRPOINTER_REG_26_ & ~n38978;
  assign n39089 = P1_P2_INSTADDRPOINTER_REG_26_ & n38978;
  assign n39090 = ~n39088 & ~n39089;
  assign n39091 = n34683 & n39090;
  assign n39092 = n36771 & ~n39058;
  assign n39093 = ~n39091 & ~n39092;
  assign n39094 = n36760 & ~n39058;
  assign n39095 = n36764 & ~n39058;
  assign n39096 = n34726 & ~n39058;
  assign n39097 = ~n39094 & ~n39095;
  assign n39098 = ~n39096 & n39097;
  assign n39099 = n39082 & n39087;
  assign n39100 = n39093 & n39099;
  assign n39101 = n39098 & n39100;
  assign n39102 = n39054 & ~n39059;
  assign n39103 = n39062 & n39102;
  assign n39104 = n39075 & n39103;
  assign n39105 = n39101 & n39104;
  assign n39106 = n36647 & ~n39105;
  assign n39107 = ~n39034 & ~n39035;
  assign n6681 = n39106 | ~n39107;
  assign n39109 = P1_P2_INSTADDRPOINTER_REG_27_ & n36646;
  assign n39110 = P1_P2_REIP_REG_27_ & n36791;
  assign n39111 = ~n39004 & ~n39036;
  assign n39112 = ~n39001 & ~n39038;
  assign n39113 = n39111 & ~n39112;
  assign n39114 = ~P1_P2_INSTADDRPOINTER_REG_27_ & ~n37582;
  assign n39115 = P1_P2_INSTADDRPOINTER_REG_27_ & n37582;
  assign n39116 = ~n39114 & ~n39115;
  assign n39117 = n39113 & ~n39116;
  assign n39118 = ~n39113 & n39116;
  assign n39119 = ~n39117 & ~n39118;
  assign n39120 = n36752 & ~n39119;
  assign n39121 = ~P1_P2_INSTADDRPOINTER_REG_27_ & n39051;
  assign n39122 = P1_P2_INSTADDRPOINTER_REG_27_ & ~n39051;
  assign n39123 = ~n39121 & ~n39122;
  assign n39124 = n36754 & ~n39123;
  assign n39125 = ~n39120 & ~n39124;
  assign n39126 = P1_P2_INSTADDRPOINTER_REG_26_ & n39055;
  assign n39127 = ~P1_P2_INSTADDRPOINTER_REG_27_ & n39126;
  assign n39128 = P1_P2_INSTADDRPOINTER_REG_27_ & ~n39126;
  assign n39129 = ~n39127 & ~n39128;
  assign n39130 = ~n34769 & ~n39129;
  assign n39131 = n34879 & ~n39129;
  assign n39132 = n34722 & ~n39129;
  assign n39133 = ~n39131 & ~n39132;
  assign n39134 = P1_P2_INSTADDRPOINTER_REG_26_ & n39063;
  assign n39135 = ~P1_P2_INSTADDRPOINTER_REG_27_ & n39134;
  assign n39136 = P1_P2_INSTADDRPOINTER_REG_27_ & ~n39134;
  assign n39137 = ~n39135 & ~n39136;
  assign n39138 = n34840 & ~n39137;
  assign n39139 = n34841 & ~n39137;
  assign n39140 = n36655 & ~n39129;
  assign n39141 = n34656 & ~n39137;
  assign n39142 = n36658 & ~n39129;
  assign n39143 = ~n39141 & ~n39142;
  assign n39144 = ~n39138 & ~n39139;
  assign n39145 = ~n39140 & n39144;
  assign n39146 = n39143 & n39145;
  assign n39147 = P1_P2_INSTADDRPOINTER_REG_26_ & n39076;
  assign n39148 = ~P1_P2_INSTADDRPOINTER_REG_27_ & n39147;
  assign n39149 = P1_P2_INSTADDRPOINTER_REG_27_ & ~n39147;
  assign n39150 = ~n39148 & ~n39149;
  assign n39151 = n34680 & ~n39150;
  assign n39152 = n34672 & ~n39150;
  assign n39153 = ~n39151 & ~n39152;
  assign n39154 = n34582 & ~n39137;
  assign n39155 = n34660 & ~n39137;
  assign n39156 = n34664 & ~n39137;
  assign n39157 = ~n39154 & ~n39155;
  assign n39158 = ~n39156 & n39157;
  assign n39159 = ~P1_P2_INSTADDRPOINTER_REG_27_ & n39089;
  assign n39160 = P1_P2_INSTADDRPOINTER_REG_27_ & ~n39089;
  assign n39161 = ~n39159 & ~n39160;
  assign n39162 = n34683 & ~n39161;
  assign n39163 = n36771 & ~n39129;
  assign n39164 = ~n39162 & ~n39163;
  assign n39165 = n36760 & ~n39129;
  assign n39166 = n36764 & ~n39129;
  assign n39167 = n34726 & ~n39129;
  assign n39168 = ~n39165 & ~n39166;
  assign n39169 = ~n39167 & n39168;
  assign n39170 = n39153 & n39158;
  assign n39171 = n39164 & n39170;
  assign n39172 = n39169 & n39171;
  assign n39173 = n39125 & ~n39130;
  assign n39174 = n39133 & n39173;
  assign n39175 = n39146 & n39174;
  assign n39176 = n39172 & n39175;
  assign n39177 = n36647 & ~n39176;
  assign n39178 = ~n39109 & ~n39110;
  assign n6686 = n39177 | ~n39178;
  assign n39180 = P1_P2_INSTADDRPOINTER_REG_28_ & n36646;
  assign n39181 = P1_P2_REIP_REG_28_ & n36791;
  assign n39182 = P1_P2_INSTADDRPOINTER_REG_27_ & P1_P2_INSTADDRPOINTER_REG_28_;
  assign n39183 = ~n39113 & n39182;
  assign n39184 = n37582 & ~n39183;
  assign n39185 = P1_P2_INSTADDRPOINTER_REG_28_ & ~n37582;
  assign n39186 = ~P1_P2_INSTADDRPOINTER_REG_27_ & ~n39004;
  assign n39187 = ~n39036 & n39186;
  assign n39188 = ~n39112 & n39187;
  assign n39189 = ~n39184 & ~n39185;
  assign n39190 = ~n39188 & n39189;
  assign n39191 = P1_P2_INSTADDRPOINTER_REG_28_ & n39188;
  assign n39192 = ~n37582 & ~n39191;
  assign n39193 = P1_P2_INSTADDRPOINTER_REG_28_ & n37582;
  assign n39194 = P1_P2_INSTADDRPOINTER_REG_27_ & ~n39113;
  assign n39195 = ~n39192 & ~n39193;
  assign n39196 = ~n39194 & n39195;
  assign n39197 = ~n39190 & ~n39196;
  assign n39198 = n36752 & n39197;
  assign n39199 = P1_P2_INSTADDRPOINTER_REG_27_ & n39051;
  assign n39200 = ~P1_P2_INSTADDRPOINTER_REG_28_ & ~n39199;
  assign n39201 = n39051 & n39182;
  assign n39202 = ~n39200 & ~n39201;
  assign n39203 = n36754 & n39202;
  assign n39204 = ~n39198 & ~n39203;
  assign n39205 = P1_P2_INSTADDRPOINTER_REG_27_ & n39126;
  assign n39206 = ~P1_P2_INSTADDRPOINTER_REG_28_ & n39205;
  assign n39207 = P1_P2_INSTADDRPOINTER_REG_28_ & ~n39205;
  assign n39208 = ~n39206 & ~n39207;
  assign n39209 = ~n34769 & ~n39208;
  assign n39210 = n34879 & ~n39208;
  assign n39211 = n34722 & ~n39208;
  assign n39212 = ~n39210 & ~n39211;
  assign n39213 = P1_P2_INSTADDRPOINTER_REG_27_ & n39134;
  assign n39214 = ~P1_P2_INSTADDRPOINTER_REG_28_ & n39213;
  assign n39215 = P1_P2_INSTADDRPOINTER_REG_28_ & ~n39213;
  assign n39216 = ~n39214 & ~n39215;
  assign n39217 = n34840 & ~n39216;
  assign n39218 = n34841 & ~n39216;
  assign n39219 = n36655 & ~n39208;
  assign n39220 = n34656 & ~n39216;
  assign n39221 = n36658 & ~n39208;
  assign n39222 = ~n39220 & ~n39221;
  assign n39223 = ~n39217 & ~n39218;
  assign n39224 = ~n39219 & n39223;
  assign n39225 = n39222 & n39224;
  assign n39226 = P1_P2_INSTADDRPOINTER_REG_27_ & n39147;
  assign n39227 = ~P1_P2_INSTADDRPOINTER_REG_28_ & n39226;
  assign n39228 = P1_P2_INSTADDRPOINTER_REG_28_ & ~n39226;
  assign n39229 = ~n39227 & ~n39228;
  assign n39230 = n34680 & ~n39229;
  assign n39231 = n34672 & ~n39229;
  assign n39232 = ~n39230 & ~n39231;
  assign n39233 = n34582 & ~n39216;
  assign n39234 = n34660 & ~n39216;
  assign n39235 = n34664 & ~n39216;
  assign n39236 = ~n39233 & ~n39234;
  assign n39237 = ~n39235 & n39236;
  assign n39238 = P1_P2_INSTADDRPOINTER_REG_27_ & n39089;
  assign n39239 = ~P1_P2_INSTADDRPOINTER_REG_28_ & ~n39238;
  assign n39240 = n39089 & n39182;
  assign n39241 = ~n39239 & ~n39240;
  assign n39242 = n34683 & n39241;
  assign n39243 = n36771 & ~n39208;
  assign n39244 = ~n39242 & ~n39243;
  assign n39245 = n36760 & ~n39208;
  assign n39246 = n36764 & ~n39208;
  assign n39247 = n34726 & ~n39208;
  assign n39248 = ~n39245 & ~n39246;
  assign n39249 = ~n39247 & n39248;
  assign n39250 = n39232 & n39237;
  assign n39251 = n39244 & n39250;
  assign n39252 = n39249 & n39251;
  assign n39253 = n39204 & ~n39209;
  assign n39254 = n39212 & n39253;
  assign n39255 = n39225 & n39254;
  assign n39256 = n39252 & n39255;
  assign n39257 = n36647 & ~n39256;
  assign n39258 = ~n39180 & ~n39181;
  assign n6691 = n39257 | ~n39258;
  assign n39260 = P1_P2_INSTADDRPOINTER_REG_29_ & n36646;
  assign n39261 = P1_P2_REIP_REG_29_ & n36791;
  assign n39262 = ~n37582 & ~n39188;
  assign n39263 = ~n39185 & ~n39262;
  assign n39264 = ~n39183 & n39263;
  assign n39265 = ~P1_P2_INSTADDRPOINTER_REG_29_ & ~n37582;
  assign n39266 = P1_P2_INSTADDRPOINTER_REG_29_ & n37582;
  assign n39267 = ~n39265 & ~n39266;
  assign n39268 = n39264 & ~n39267;
  assign n39269 = ~n39264 & n39267;
  assign n39270 = ~n39268 & ~n39269;
  assign n39271 = n36752 & ~n39270;
  assign n39272 = ~P1_P2_INSTADDRPOINTER_REG_29_ & ~n39201;
  assign n39273 = P1_P2_INSTADDRPOINTER_REG_29_ & n39201;
  assign n39274 = ~n39272 & ~n39273;
  assign n39275 = n36754 & n39274;
  assign n39276 = ~n39271 & ~n39275;
  assign n39277 = P1_P2_INSTADDRPOINTER_REG_28_ & n39205;
  assign n39278 = ~P1_P2_INSTADDRPOINTER_REG_29_ & n39277;
  assign n39279 = P1_P2_INSTADDRPOINTER_REG_29_ & ~n39277;
  assign n39280 = ~n39278 & ~n39279;
  assign n39281 = ~n34769 & ~n39280;
  assign n39282 = n34879 & ~n39280;
  assign n39283 = n34722 & ~n39280;
  assign n39284 = ~n39282 & ~n39283;
  assign n39285 = P1_P2_INSTADDRPOINTER_REG_28_ & n39213;
  assign n39286 = ~P1_P2_INSTADDRPOINTER_REG_29_ & n39285;
  assign n39287 = P1_P2_INSTADDRPOINTER_REG_29_ & ~n39285;
  assign n39288 = ~n39286 & ~n39287;
  assign n39289 = n34840 & ~n39288;
  assign n39290 = n34841 & ~n39288;
  assign n39291 = n36655 & ~n39280;
  assign n39292 = n34656 & ~n39288;
  assign n39293 = n36658 & ~n39280;
  assign n39294 = ~n39292 & ~n39293;
  assign n39295 = ~n39289 & ~n39290;
  assign n39296 = ~n39291 & n39295;
  assign n39297 = n39294 & n39296;
  assign n39298 = P1_P2_INSTADDRPOINTER_REG_28_ & n39226;
  assign n39299 = ~P1_P2_INSTADDRPOINTER_REG_29_ & n39298;
  assign n39300 = P1_P2_INSTADDRPOINTER_REG_29_ & ~n39298;
  assign n39301 = ~n39299 & ~n39300;
  assign n39302 = n34680 & ~n39301;
  assign n39303 = n34672 & ~n39301;
  assign n39304 = ~n39302 & ~n39303;
  assign n39305 = n34582 & ~n39288;
  assign n39306 = n34660 & ~n39288;
  assign n39307 = n34664 & ~n39288;
  assign n39308 = ~n39305 & ~n39306;
  assign n39309 = ~n39307 & n39308;
  assign n39310 = ~P1_P2_INSTADDRPOINTER_REG_29_ & ~n39240;
  assign n39311 = P1_P2_INSTADDRPOINTER_REG_29_ & n39240;
  assign n39312 = ~n39310 & ~n39311;
  assign n39313 = n34683 & n39312;
  assign n39314 = n36771 & ~n39280;
  assign n39315 = ~n39313 & ~n39314;
  assign n39316 = n36760 & ~n39280;
  assign n39317 = n36764 & ~n39280;
  assign n39318 = n34726 & ~n39280;
  assign n39319 = ~n39316 & ~n39317;
  assign n39320 = ~n39318 & n39319;
  assign n39321 = n39304 & n39309;
  assign n39322 = n39315 & n39321;
  assign n39323 = n39320 & n39322;
  assign n39324 = n39276 & ~n39281;
  assign n39325 = n39284 & n39324;
  assign n39326 = n39297 & n39325;
  assign n39327 = n39323 & n39326;
  assign n39328 = n36647 & ~n39327;
  assign n39329 = ~n39260 & ~n39261;
  assign n6696 = n39328 | ~n39329;
  assign n39331 = P1_P2_INSTADDRPOINTER_REG_30_ & n36646;
  assign n39332 = P1_P2_REIP_REG_30_ & n36791;
  assign n39333 = ~P1_P2_INSTADDRPOINTER_REG_30_ & ~n37582;
  assign n39334 = P1_P2_INSTADDRPOINTER_REG_30_ & n37582;
  assign n39335 = ~n39333 & ~n39334;
  assign n39336 = P1_P2_INSTADDRPOINTER_REG_29_ & ~n37582;
  assign n39337 = ~P1_P2_INSTADDRPOINTER_REG_29_ & n37582;
  assign n39338 = ~n39264 & ~n39337;
  assign n39339 = ~n39336 & ~n39338;
  assign n39340 = ~n39335 & n39339;
  assign n39341 = n39335 & ~n39339;
  assign n39342 = ~n39340 & ~n39341;
  assign n39343 = n36752 & ~n39342;
  assign n39344 = ~P1_P2_INSTADDRPOINTER_REG_30_ & n39273;
  assign n39345 = P1_P2_INSTADDRPOINTER_REG_30_ & ~n39273;
  assign n39346 = ~n39344 & ~n39345;
  assign n39347 = n36754 & ~n39346;
  assign n39348 = ~n39343 & ~n39347;
  assign n39349 = P1_P2_INSTADDRPOINTER_REG_29_ & n39277;
  assign n39350 = ~P1_P2_INSTADDRPOINTER_REG_30_ & n39349;
  assign n39351 = P1_P2_INSTADDRPOINTER_REG_30_ & ~n39349;
  assign n39352 = ~n39350 & ~n39351;
  assign n39353 = ~n34769 & ~n39352;
  assign n39354 = n34879 & ~n39352;
  assign n39355 = n34722 & ~n39352;
  assign n39356 = ~n39354 & ~n39355;
  assign n39357 = P1_P2_INSTADDRPOINTER_REG_29_ & n39285;
  assign n39358 = ~P1_P2_INSTADDRPOINTER_REG_30_ & n39357;
  assign n39359 = P1_P2_INSTADDRPOINTER_REG_30_ & ~n39357;
  assign n39360 = ~n39358 & ~n39359;
  assign n39361 = n34840 & ~n39360;
  assign n39362 = n34841 & ~n39360;
  assign n39363 = n36655 & ~n39352;
  assign n39364 = n34656 & ~n39360;
  assign n39365 = n36658 & ~n39352;
  assign n39366 = ~n39364 & ~n39365;
  assign n39367 = ~n39361 & ~n39362;
  assign n39368 = ~n39363 & n39367;
  assign n39369 = n39366 & n39368;
  assign n39370 = P1_P2_INSTADDRPOINTER_REG_29_ & n39298;
  assign n39371 = ~P1_P2_INSTADDRPOINTER_REG_30_ & n39370;
  assign n39372 = P1_P2_INSTADDRPOINTER_REG_30_ & ~n39370;
  assign n39373 = ~n39371 & ~n39372;
  assign n39374 = n34680 & ~n39373;
  assign n39375 = n34672 & ~n39373;
  assign n39376 = ~n39374 & ~n39375;
  assign n39377 = n34582 & ~n39360;
  assign n39378 = n34660 & ~n39360;
  assign n39379 = n34664 & ~n39360;
  assign n39380 = ~n39377 & ~n39378;
  assign n39381 = ~n39379 & n39380;
  assign n39382 = ~P1_P2_INSTADDRPOINTER_REG_30_ & n39311;
  assign n39383 = P1_P2_INSTADDRPOINTER_REG_30_ & ~n39311;
  assign n39384 = ~n39382 & ~n39383;
  assign n39385 = n34683 & ~n39384;
  assign n39386 = n36771 & ~n39352;
  assign n39387 = ~n39385 & ~n39386;
  assign n39388 = n36760 & ~n39352;
  assign n39389 = n36764 & ~n39352;
  assign n39390 = n34726 & ~n39352;
  assign n39391 = ~n39388 & ~n39389;
  assign n39392 = ~n39390 & n39391;
  assign n39393 = n39376 & n39381;
  assign n39394 = n39387 & n39393;
  assign n39395 = n39392 & n39394;
  assign n39396 = n39348 & ~n39353;
  assign n39397 = n39356 & n39396;
  assign n39398 = n39369 & n39397;
  assign n39399 = n39395 & n39398;
  assign n39400 = n36647 & ~n39399;
  assign n39401 = ~n39331 & ~n39332;
  assign n6701 = n39400 | ~n39401;
  assign n39403 = P1_P2_INSTADDRPOINTER_REG_31_ & n36646;
  assign n39404 = P1_P2_REIP_REG_31_ & n36791;
  assign n39405 = P1_P2_INSTADDRPOINTER_REG_30_ & n39311;
  assign n39406 = ~P1_P2_INSTADDRPOINTER_REG_31_ & n39405;
  assign n39407 = P1_P2_INSTADDRPOINTER_REG_31_ & ~n39405;
  assign n39408 = ~n39406 & ~n39407;
  assign n39409 = n34683 & ~n39408;
  assign n39410 = P1_P2_INSTADDRPOINTER_REG_30_ & n39349;
  assign n39411 = ~P1_P2_INSTADDRPOINTER_REG_31_ & n39410;
  assign n39412 = P1_P2_INSTADDRPOINTER_REG_31_ & ~n39410;
  assign n39413 = ~n39411 & ~n39412;
  assign n39414 = n36771 & ~n39413;
  assign n39415 = n34726 & ~n39413;
  assign n39416 = ~n39414 & ~n39415;
  assign n39417 = P1_P2_INSTADDRPOINTER_REG_30_ & n39357;
  assign n39418 = ~P1_P2_INSTADDRPOINTER_REG_31_ & n39417;
  assign n39419 = P1_P2_INSTADDRPOINTER_REG_31_ & ~n39417;
  assign n39420 = ~n39418 & ~n39419;
  assign n39421 = n34664 & ~n39420;
  assign n39422 = n34582 & ~n39420;
  assign n39423 = P1_P2_INSTADDRPOINTER_REG_30_ & n39370;
  assign n39424 = ~P1_P2_INSTADDRPOINTER_REG_31_ & n39423;
  assign n39425 = P1_P2_INSTADDRPOINTER_REG_31_ & ~n39423;
  assign n39426 = ~n39424 & ~n39425;
  assign n39427 = n34672 & ~n39426;
  assign n39428 = ~n39421 & ~n39422;
  assign n39429 = ~n39427 & n39428;
  assign n39430 = n36760 & ~n39413;
  assign n39431 = n36764 & ~n39413;
  assign n39432 = n34680 & ~n39426;
  assign n39433 = ~n39431 & ~n39432;
  assign n39434 = n39429 & ~n39430;
  assign n39435 = n39433 & n39434;
  assign n39436 = ~n39403 & ~n39404;
  assign n39437 = ~n39409 & n39436;
  assign n39438 = n39416 & n39437;
  assign n39439 = n39435 & n39438;
  assign n39440 = P1_P2_INSTADDRPOINTER_REG_30_ & P1_P2_INSTADDRPOINTER_REG_31_;
  assign n39441 = ~n39339 & n39440;
  assign n39442 = n37582 & ~n39441;
  assign n39443 = P1_P2_INSTADDRPOINTER_REG_31_ & ~n37582;
  assign n39444 = ~P1_P2_INSTADDRPOINTER_REG_30_ & n39339;
  assign n39445 = ~n39442 & ~n39443;
  assign n39446 = ~n39444 & n39445;
  assign n39447 = ~P1_P2_INSTADDRPOINTER_REG_30_ & P1_P2_INSTADDRPOINTER_REG_31_;
  assign n39448 = ~n39336 & n39447;
  assign n39449 = ~n39338 & n39448;
  assign n39450 = ~n37582 & ~n39449;
  assign n39451 = P1_P2_INSTADDRPOINTER_REG_31_ & n37582;
  assign n39452 = P1_P2_INSTADDRPOINTER_REG_30_ & ~n39339;
  assign n39453 = ~n39450 & ~n39451;
  assign n39454 = ~n39452 & n39453;
  assign n39455 = ~n39446 & ~n39454;
  assign n39456 = n36752 & n39455;
  assign n39457 = P1_P2_INSTADDRPOINTER_REG_30_ & n39273;
  assign n39458 = ~P1_P2_INSTADDRPOINTER_REG_31_ & n39457;
  assign n39459 = P1_P2_INSTADDRPOINTER_REG_31_ & ~n39457;
  assign n39460 = ~n39458 & ~n39459;
  assign n39461 = n36754 & ~n39460;
  assign n39462 = ~n39456 & ~n39461;
  assign n39463 = ~n34769 & ~n39413;
  assign n39464 = n34879 & ~n39413;
  assign n39465 = n34722 & ~n39413;
  assign n39466 = ~n39464 & ~n39465;
  assign n39467 = n34841 & ~n39420;
  assign n39468 = n39466 & ~n39467;
  assign n39469 = n36655 & ~n39413;
  assign n39470 = n34840 & ~n39420;
  assign n39471 = n34660 & ~n39420;
  assign n39472 = n34656 & ~n39420;
  assign n39473 = n36658 & ~n39413;
  assign n39474 = ~n39471 & ~n39472;
  assign n39475 = ~n39473 & n39474;
  assign n39476 = ~n39469 & ~n39470;
  assign n39477 = n39475 & n39476;
  assign n39478 = n39462 & ~n39463;
  assign n39479 = n39468 & n39478;
  assign n39480 = n39477 & n39479;
  assign n39481 = n39439 & n39480;
  assign n39482 = ~n36647 & ~n39403;
  assign n39483 = ~n39404 & n39482;
  assign n6706 = ~n39481 & ~n39483;
  assign n39485 = P1_P2_STATE2_REG_0_ & ~n34549;
  assign n39486 = ~P1_P2_STATE2_REG_0_ & ~n36614;
  assign n39487 = n34683 & n34686;
  assign n39488 = n34688 & n34692;
  assign n39489 = ~n39487 & ~n39488;
  assign n39490 = n34935 & ~n39489;
  assign n39491 = ~n39486 & ~n39490;
  assign n39492 = n39485 & ~n39491;
  assign n39493 = ~n36751 & n39492;
  assign n39494 = ~n36720 & n39493;
  assign n39495 = n36751 & n39492;
  assign n39496 = ~n36720 & n39495;
  assign n39497 = P1_P2_STATE2_REG_1_ & ~n39491;
  assign n39498 = P1_P2_STATEBS16_REG & n39497;
  assign n39499 = P1_P2_PHYADDRPOINTER_REG_0_ & n39498;
  assign n39500 = ~P1_P2_STATEBS16_REG & n39497;
  assign n39501 = P1_P2_PHYADDRPOINTER_REG_0_ & n39500;
  assign n39502 = P1_P2_PHYADDRPOINTER_REG_0_ & n39491;
  assign n39503 = P1_P2_STATE2_REG_0_ & n34549;
  assign n39504 = ~n39491 & n39503;
  assign n39505 = ~n36768 & n39504;
  assign n39506 = P1_P2_STATE2_REG_2_ & ~P1_P2_STATE2_REG_0_;
  assign n39507 = ~n39491 & n39506;
  assign n39508 = P1_P2_PHYADDRPOINTER_REG_0_ & n39507;
  assign n39509 = n34951 & ~n39491;
  assign n39510 = P1_P2_REIP_REG_0_ & n39509;
  assign n39511 = ~n39502 & ~n39505;
  assign n39512 = ~n39508 & n39511;
  assign n39513 = ~n39510 & n39512;
  assign n39514 = ~n39494 & ~n39496;
  assign n39515 = ~n39499 & n39514;
  assign n39516 = ~n39501 & n39515;
  assign n6711 = ~n39513 | ~n39516;
  assign n39518 = ~n36892 & n39493;
  assign n39519 = ~n36842 & n39495;
  assign n39520 = P1_P2_PHYADDRPOINTER_REG_1_ & n39498;
  assign n39521 = ~P1_P2_PHYADDRPOINTER_REG_1_ & n39500;
  assign n39522 = P1_P2_PHYADDRPOINTER_REG_1_ & n39491;
  assign n39523 = ~n36872 & n39504;
  assign n39524 = ~P1_P2_PHYADDRPOINTER_REG_1_ & n39507;
  assign n39525 = P1_P2_REIP_REG_1_ & n39509;
  assign n39526 = ~n39522 & ~n39523;
  assign n39527 = ~n39524 & n39526;
  assign n39528 = ~n39525 & n39527;
  assign n39529 = ~n39518 & ~n39519;
  assign n39530 = ~n39520 & n39529;
  assign n39531 = ~n39521 & n39530;
  assign n6716 = ~n39528 | ~n39531;
  assign n39533 = ~n36977 & n39493;
  assign n39534 = ~n36964 & n39495;
  assign n39535 = ~P1_P2_PHYADDRPOINTER_REG_2_ & n39498;
  assign n39536 = P1_P2_PHYADDRPOINTER_REG_1_ & ~P1_P2_PHYADDRPOINTER_REG_2_;
  assign n39537 = ~P1_P2_PHYADDRPOINTER_REG_1_ & P1_P2_PHYADDRPOINTER_REG_2_;
  assign n39538 = ~n39536 & ~n39537;
  assign n39539 = n39500 & ~n39538;
  assign n39540 = n39507 & ~n39538;
  assign n39541 = P1_P2_REIP_REG_2_ & n39509;
  assign n39542 = P1_P2_PHYADDRPOINTER_REG_2_ & n39491;
  assign n39543 = ~n37014 & n39504;
  assign n39544 = ~n39540 & ~n39541;
  assign n39545 = ~n39542 & n39544;
  assign n39546 = ~n39543 & n39545;
  assign n39547 = ~n39533 & ~n39534;
  assign n39548 = ~n39535 & n39547;
  assign n39549 = ~n39539 & n39548;
  assign n6721 = ~n39546 | ~n39549;
  assign n39551 = ~n37092 & n39493;
  assign n39552 = n37107 & n39495;
  assign n39553 = P1_P2_PHYADDRPOINTER_REG_2_ & ~P1_P2_PHYADDRPOINTER_REG_3_;
  assign n39554 = ~P1_P2_PHYADDRPOINTER_REG_2_ & P1_P2_PHYADDRPOINTER_REG_3_;
  assign n39555 = ~n39553 & ~n39554;
  assign n39556 = n39498 & ~n39555;
  assign n39557 = P1_P2_PHYADDRPOINTER_REG_1_ & P1_P2_PHYADDRPOINTER_REG_2_;
  assign n39558 = ~P1_P2_PHYADDRPOINTER_REG_3_ & n39557;
  assign n39559 = P1_P2_PHYADDRPOINTER_REG_3_ & ~n39557;
  assign n39560 = ~n39558 & ~n39559;
  assign n39561 = n39500 & ~n39560;
  assign n39562 = n39507 & ~n39560;
  assign n39563 = P1_P2_REIP_REG_3_ & n39509;
  assign n39564 = P1_P2_PHYADDRPOINTER_REG_3_ & n39491;
  assign n39565 = n37145 & n39504;
  assign n39566 = ~n39562 & ~n39563;
  assign n39567 = ~n39564 & n39566;
  assign n39568 = ~n39565 & n39567;
  assign n39569 = ~n39551 & ~n39552;
  assign n39570 = ~n39556 & n39569;
  assign n39571 = ~n39561 & n39570;
  assign n6726 = ~n39568 | ~n39571;
  assign n39573 = P1_P2_PHYADDRPOINTER_REG_2_ & P1_P2_PHYADDRPOINTER_REG_3_;
  assign n39574 = ~P1_P2_PHYADDRPOINTER_REG_4_ & n39573;
  assign n39575 = P1_P2_PHYADDRPOINTER_REG_4_ & ~n39573;
  assign n39576 = ~n39574 & ~n39575;
  assign n39577 = n39498 & ~n39576;
  assign n39578 = P1_P2_PHYADDRPOINTER_REG_3_ & n39557;
  assign n39579 = ~P1_P2_PHYADDRPOINTER_REG_4_ & n39578;
  assign n39580 = P1_P2_PHYADDRPOINTER_REG_4_ & ~n39578;
  assign n39581 = ~n39579 & ~n39580;
  assign n39582 = n39500 & ~n39581;
  assign n39583 = n37220 & n39495;
  assign n39584 = ~n37242 & n39493;
  assign n39585 = n39507 & ~n39581;
  assign n39586 = P1_P2_REIP_REG_4_ & n39509;
  assign n39587 = P1_P2_PHYADDRPOINTER_REG_4_ & n39491;
  assign n39588 = ~n37281 & n39504;
  assign n39589 = ~n39585 & ~n39586;
  assign n39590 = ~n39587 & n39589;
  assign n39591 = ~n39588 & n39590;
  assign n39592 = ~n39577 & ~n39582;
  assign n39593 = ~n39583 & n39592;
  assign n39594 = ~n39584 & n39593;
  assign n6731 = ~n39591 | ~n39594;
  assign n39596 = P1_P2_PHYADDRPOINTER_REG_4_ & n39573;
  assign n39597 = ~P1_P2_PHYADDRPOINTER_REG_5_ & n39596;
  assign n39598 = P1_P2_PHYADDRPOINTER_REG_5_ & ~n39596;
  assign n39599 = ~n39597 & ~n39598;
  assign n39600 = n39498 & ~n39599;
  assign n39601 = P1_P2_PHYADDRPOINTER_REG_4_ & n39578;
  assign n39602 = ~P1_P2_PHYADDRPOINTER_REG_5_ & n39601;
  assign n39603 = P1_P2_PHYADDRPOINTER_REG_5_ & ~n39601;
  assign n39604 = ~n39602 & ~n39603;
  assign n39605 = n39500 & ~n39604;
  assign n39606 = ~n37357 & n39493;
  assign n39607 = ~n37375 & n39495;
  assign n39608 = n39507 & ~n39604;
  assign n39609 = P1_P2_REIP_REG_5_ & n39509;
  assign n39610 = P1_P2_PHYADDRPOINTER_REG_5_ & n39491;
  assign n39611 = n37414 & n39504;
  assign n39612 = ~n39608 & ~n39609;
  assign n39613 = ~n39610 & n39612;
  assign n39614 = ~n39611 & n39613;
  assign n39615 = ~n39600 & ~n39605;
  assign n39616 = ~n39606 & n39615;
  assign n39617 = ~n39607 & n39616;
  assign n6736 = ~n39614 | ~n39617;
  assign n39619 = P1_P2_PHYADDRPOINTER_REG_5_ & n39596;
  assign n39620 = ~P1_P2_PHYADDRPOINTER_REG_6_ & n39619;
  assign n39621 = P1_P2_PHYADDRPOINTER_REG_6_ & ~n39619;
  assign n39622 = ~n39620 & ~n39621;
  assign n39623 = n39498 & ~n39622;
  assign n39624 = P1_P2_PHYADDRPOINTER_REG_5_ & n39601;
  assign n39625 = ~P1_P2_PHYADDRPOINTER_REG_6_ & n39624;
  assign n39626 = P1_P2_PHYADDRPOINTER_REG_6_ & ~n39624;
  assign n39627 = ~n39625 & ~n39626;
  assign n39628 = n39500 & ~n39627;
  assign n39629 = ~n37488 & n39493;
  assign n39630 = ~n37507 & n39495;
  assign n39631 = n39507 & ~n39627;
  assign n39632 = P1_P2_REIP_REG_6_ & n39509;
  assign n39633 = P1_P2_PHYADDRPOINTER_REG_6_ & n39491;
  assign n39634 = ~n37545 & n39504;
  assign n39635 = ~n39631 & ~n39632;
  assign n39636 = ~n39633 & n39635;
  assign n39637 = ~n39634 & n39636;
  assign n39638 = ~n39623 & ~n39628;
  assign n39639 = ~n39629 & n39638;
  assign n39640 = ~n39630 & n39639;
  assign n6741 = ~n39637 | ~n39640;
  assign n39642 = P1_P2_PHYADDRPOINTER_REG_6_ & n39619;
  assign n39643 = ~P1_P2_PHYADDRPOINTER_REG_7_ & n39642;
  assign n39644 = P1_P2_PHYADDRPOINTER_REG_7_ & ~n39642;
  assign n39645 = ~n39643 & ~n39644;
  assign n39646 = n39498 & ~n39645;
  assign n39647 = P1_P2_PHYADDRPOINTER_REG_6_ & n39624;
  assign n39648 = ~P1_P2_PHYADDRPOINTER_REG_7_ & n39647;
  assign n39649 = P1_P2_PHYADDRPOINTER_REG_7_ & ~n39647;
  assign n39650 = ~n39648 & ~n39649;
  assign n39651 = n39500 & ~n39650;
  assign n39652 = ~n37589 & n39493;
  assign n39653 = ~n37607 & n39495;
  assign n39654 = n39507 & ~n39650;
  assign n39655 = P1_P2_REIP_REG_7_ & n39509;
  assign n39656 = P1_P2_PHYADDRPOINTER_REG_7_ & n39491;
  assign n39657 = ~n37643 & n39504;
  assign n39658 = ~n39654 & ~n39655;
  assign n39659 = ~n39656 & n39658;
  assign n39660 = ~n39657 & n39659;
  assign n39661 = ~n39646 & ~n39651;
  assign n39662 = ~n39652 & n39661;
  assign n39663 = ~n39653 & n39662;
  assign n6746 = ~n39660 | ~n39663;
  assign n39665 = P1_P2_PHYADDRPOINTER_REG_7_ & n39642;
  assign n39666 = ~P1_P2_PHYADDRPOINTER_REG_8_ & n39665;
  assign n39667 = P1_P2_PHYADDRPOINTER_REG_8_ & ~n39665;
  assign n39668 = ~n39666 & ~n39667;
  assign n39669 = n39498 & ~n39668;
  assign n39670 = P1_P2_PHYADDRPOINTER_REG_7_ & n39647;
  assign n39671 = ~P1_P2_PHYADDRPOINTER_REG_8_ & n39670;
  assign n39672 = P1_P2_PHYADDRPOINTER_REG_8_ & ~n39670;
  assign n39673 = ~n39671 & ~n39672;
  assign n39674 = n39500 & ~n39673;
  assign n39675 = ~n37683 & n39493;
  assign n39676 = ~n37699 & n39495;
  assign n39677 = n39507 & ~n39673;
  assign n39678 = P1_P2_REIP_REG_8_ & n39509;
  assign n39679 = P1_P2_PHYADDRPOINTER_REG_8_ & n39491;
  assign n39680 = ~n37733 & n39504;
  assign n39681 = ~n39677 & ~n39678;
  assign n39682 = ~n39679 & n39681;
  assign n39683 = ~n39680 & n39682;
  assign n39684 = ~n39669 & ~n39674;
  assign n39685 = ~n39675 & n39684;
  assign n39686 = ~n39676 & n39685;
  assign n6751 = ~n39683 | ~n39686;
  assign n39688 = P1_P2_PHYADDRPOINTER_REG_8_ & n39665;
  assign n39689 = ~P1_P2_PHYADDRPOINTER_REG_9_ & n39688;
  assign n39690 = P1_P2_PHYADDRPOINTER_REG_9_ & ~n39688;
  assign n39691 = ~n39689 & ~n39690;
  assign n39692 = n39498 & ~n39691;
  assign n39693 = P1_P2_PHYADDRPOINTER_REG_8_ & n39670;
  assign n39694 = ~P1_P2_PHYADDRPOINTER_REG_9_ & n39693;
  assign n39695 = P1_P2_PHYADDRPOINTER_REG_9_ & ~n39693;
  assign n39696 = ~n39694 & ~n39695;
  assign n39697 = n39500 & ~n39696;
  assign n39698 = ~n37776 & n39493;
  assign n39699 = n37787 & n39495;
  assign n39700 = n39507 & ~n39696;
  assign n39701 = P1_P2_REIP_REG_9_ & n39509;
  assign n39702 = P1_P2_PHYADDRPOINTER_REG_9_ & n39491;
  assign n39703 = n37816 & n39504;
  assign n39704 = ~n39700 & ~n39701;
  assign n39705 = ~n39702 & n39704;
  assign n39706 = ~n39703 & n39705;
  assign n39707 = ~n39692 & ~n39697;
  assign n39708 = ~n39698 & n39707;
  assign n39709 = ~n39699 & n39708;
  assign n6756 = ~n39706 | ~n39709;
  assign n39711 = P1_P2_PHYADDRPOINTER_REG_9_ & n39688;
  assign n39712 = ~P1_P2_PHYADDRPOINTER_REG_10_ & n39711;
  assign n39713 = P1_P2_PHYADDRPOINTER_REG_10_ & ~n39711;
  assign n39714 = ~n39712 & ~n39713;
  assign n39715 = n39498 & ~n39714;
  assign n39716 = P1_P2_PHYADDRPOINTER_REG_9_ & n39693;
  assign n39717 = ~P1_P2_PHYADDRPOINTER_REG_10_ & n39716;
  assign n39718 = P1_P2_PHYADDRPOINTER_REG_10_ & ~n39716;
  assign n39719 = ~n39717 & ~n39718;
  assign n39720 = n39500 & ~n39719;
  assign n39721 = ~n37859 & n39493;
  assign n39722 = n37867 & n39495;
  assign n39723 = n39507 & ~n39719;
  assign n39724 = P1_P2_REIP_REG_10_ & n39509;
  assign n39725 = P1_P2_PHYADDRPOINTER_REG_10_ & n39491;
  assign n39726 = n37892 & n39504;
  assign n39727 = ~n39723 & ~n39724;
  assign n39728 = ~n39725 & n39727;
  assign n39729 = ~n39726 & n39728;
  assign n39730 = ~n39715 & ~n39720;
  assign n39731 = ~n39721 & n39730;
  assign n39732 = ~n39722 & n39731;
  assign n6761 = ~n39729 | ~n39732;
  assign n39734 = P1_P2_PHYADDRPOINTER_REG_10_ & n39711;
  assign n39735 = ~P1_P2_PHYADDRPOINTER_REG_11_ & n39734;
  assign n39736 = P1_P2_PHYADDRPOINTER_REG_11_ & ~n39734;
  assign n39737 = ~n39735 & ~n39736;
  assign n39738 = n39498 & ~n39737;
  assign n39739 = P1_P2_PHYADDRPOINTER_REG_10_ & n39716;
  assign n39740 = ~P1_P2_PHYADDRPOINTER_REG_11_ & n39739;
  assign n39741 = P1_P2_PHYADDRPOINTER_REG_11_ & ~n39739;
  assign n39742 = ~n39740 & ~n39741;
  assign n39743 = n39500 & ~n39742;
  assign n39744 = ~n37953 & n39493;
  assign n39745 = ~n37966 & n39495;
  assign n39746 = n39507 & ~n39742;
  assign n39747 = P1_P2_REIP_REG_11_ & n39509;
  assign n39748 = P1_P2_PHYADDRPOINTER_REG_11_ & n39491;
  assign n39749 = ~n37936 & n39504;
  assign n39750 = ~n39746 & ~n39747;
  assign n39751 = ~n39748 & n39750;
  assign n39752 = ~n39749 & n39751;
  assign n39753 = ~n39738 & ~n39743;
  assign n39754 = ~n39744 & n39753;
  assign n39755 = ~n39745 & n39754;
  assign n6766 = ~n39752 | ~n39755;
  assign n39757 = P1_P2_PHYADDRPOINTER_REG_11_ & n39734;
  assign n39758 = ~P1_P2_PHYADDRPOINTER_REG_12_ & n39757;
  assign n39759 = P1_P2_PHYADDRPOINTER_REG_12_ & ~n39757;
  assign n39760 = ~n39758 & ~n39759;
  assign n39761 = n39498 & ~n39760;
  assign n39762 = P1_P2_PHYADDRPOINTER_REG_11_ & n39739;
  assign n39763 = ~P1_P2_PHYADDRPOINTER_REG_12_ & n39762;
  assign n39764 = P1_P2_PHYADDRPOINTER_REG_12_ & ~n39762;
  assign n39765 = ~n39763 & ~n39764;
  assign n39766 = n39500 & ~n39765;
  assign n39767 = ~n38007 & n39493;
  assign n39768 = n38016 & n39495;
  assign n39769 = P1_P2_PHYADDRPOINTER_REG_12_ & n39491;
  assign n39770 = P1_P2_REIP_REG_12_ & n39509;
  assign n39771 = n39507 & ~n39765;
  assign n39772 = n38042 & n39504;
  assign n39773 = ~n39769 & ~n39770;
  assign n39774 = ~n39771 & n39773;
  assign n39775 = ~n39772 & n39774;
  assign n39776 = ~n39761 & ~n39766;
  assign n39777 = ~n39767 & n39776;
  assign n39778 = ~n39768 & n39777;
  assign n6771 = ~n39775 | ~n39778;
  assign n39780 = P1_P2_PHYADDRPOINTER_REG_12_ & n39757;
  assign n39781 = ~P1_P2_PHYADDRPOINTER_REG_13_ & n39780;
  assign n39782 = P1_P2_PHYADDRPOINTER_REG_13_ & ~n39780;
  assign n39783 = ~n39781 & ~n39782;
  assign n39784 = n39498 & ~n39783;
  assign n39785 = P1_P2_PHYADDRPOINTER_REG_12_ & n39762;
  assign n39786 = ~P1_P2_PHYADDRPOINTER_REG_13_ & n39785;
  assign n39787 = P1_P2_PHYADDRPOINTER_REG_13_ & ~n39785;
  assign n39788 = ~n39786 & ~n39787;
  assign n39789 = n39500 & ~n39788;
  assign n39790 = n38085 & n39493;
  assign n39791 = n38092 & n39495;
  assign n39792 = P1_P2_PHYADDRPOINTER_REG_13_ & n39491;
  assign n39793 = P1_P2_REIP_REG_13_ & n39509;
  assign n39794 = n39507 & ~n39788;
  assign n39795 = n38117 & n39504;
  assign n39796 = ~n39792 & ~n39793;
  assign n39797 = ~n39794 & n39796;
  assign n39798 = ~n39795 & n39797;
  assign n39799 = ~n39784 & ~n39789;
  assign n39800 = ~n39790 & n39799;
  assign n39801 = ~n39791 & n39800;
  assign n6776 = ~n39798 | ~n39801;
  assign n39803 = P1_P2_PHYADDRPOINTER_REG_13_ & n39780;
  assign n39804 = ~P1_P2_PHYADDRPOINTER_REG_14_ & n39803;
  assign n39805 = P1_P2_PHYADDRPOINTER_REG_14_ & ~n39803;
  assign n39806 = ~n39804 & ~n39805;
  assign n39807 = n39498 & ~n39806;
  assign n39808 = P1_P2_PHYADDRPOINTER_REG_13_ & n39785;
  assign n39809 = ~P1_P2_PHYADDRPOINTER_REG_14_ & n39808;
  assign n39810 = P1_P2_PHYADDRPOINTER_REG_14_ & ~n39808;
  assign n39811 = ~n39809 & ~n39810;
  assign n39812 = n39500 & ~n39811;
  assign n39813 = ~n38188 & n39493;
  assign n39814 = ~n38192 & n39495;
  assign n39815 = P1_P2_PHYADDRPOINTER_REG_14_ & n39491;
  assign n39816 = P1_P2_REIP_REG_14_ & n39509;
  assign n39817 = n39507 & ~n39811;
  assign n39818 = ~n38161 & n39504;
  assign n39819 = ~n39815 & ~n39816;
  assign n39820 = ~n39817 & n39819;
  assign n39821 = ~n39818 & n39820;
  assign n39822 = ~n39807 & ~n39812;
  assign n39823 = ~n39813 & n39822;
  assign n39824 = ~n39814 & n39823;
  assign n6781 = ~n39821 | ~n39824;
  assign n39826 = P1_P2_PHYADDRPOINTER_REG_14_ & n39803;
  assign n39827 = ~P1_P2_PHYADDRPOINTER_REG_15_ & n39826;
  assign n39828 = P1_P2_PHYADDRPOINTER_REG_15_ & ~n39826;
  assign n39829 = ~n39827 & ~n39828;
  assign n39830 = n39498 & ~n39829;
  assign n39831 = P1_P2_PHYADDRPOINTER_REG_14_ & n39808;
  assign n39832 = ~P1_P2_PHYADDRPOINTER_REG_15_ & n39831;
  assign n39833 = P1_P2_PHYADDRPOINTER_REG_15_ & ~n39831;
  assign n39834 = ~n39832 & ~n39833;
  assign n39835 = n39500 & ~n39834;
  assign n39836 = ~n38265 & n39493;
  assign n39837 = n38270 & n39495;
  assign n39838 = P1_P2_PHYADDRPOINTER_REG_15_ & n39491;
  assign n39839 = P1_P2_REIP_REG_15_ & n39509;
  assign n39840 = n39507 & ~n39834;
  assign n39841 = n38237 & n39504;
  assign n39842 = ~n39838 & ~n39839;
  assign n39843 = ~n39840 & n39842;
  assign n39844 = ~n39841 & n39843;
  assign n39845 = ~n39830 & ~n39835;
  assign n39846 = ~n39836 & n39845;
  assign n39847 = ~n39837 & n39846;
  assign n6786 = ~n39844 | ~n39847;
  assign n39849 = P1_P2_PHYADDRPOINTER_REG_15_ & n39826;
  assign n39850 = ~P1_P2_PHYADDRPOINTER_REG_16_ & n39849;
  assign n39851 = P1_P2_PHYADDRPOINTER_REG_16_ & ~n39849;
  assign n39852 = ~n39850 & ~n39851;
  assign n39853 = n39498 & ~n39852;
  assign n39854 = P1_P2_PHYADDRPOINTER_REG_15_ & n39831;
  assign n39855 = ~P1_P2_PHYADDRPOINTER_REG_16_ & n39854;
  assign n39856 = P1_P2_PHYADDRPOINTER_REG_16_ & ~n39854;
  assign n39857 = ~n39855 & ~n39856;
  assign n39858 = n39500 & ~n39857;
  assign n39859 = ~n38329 & n39493;
  assign n39860 = ~n38342 & n39495;
  assign n39861 = P1_P2_PHYADDRPOINTER_REG_16_ & n39491;
  assign n39862 = P1_P2_REIP_REG_16_ & n39509;
  assign n39863 = n39507 & ~n39857;
  assign n39864 = ~n38312 & n39504;
  assign n39865 = ~n39861 & ~n39862;
  assign n39866 = ~n39863 & n39865;
  assign n39867 = ~n39864 & n39866;
  assign n39868 = ~n39853 & ~n39858;
  assign n39869 = ~n39859 & n39868;
  assign n39870 = ~n39860 & n39869;
  assign n6791 = ~n39867 | ~n39870;
  assign n39872 = P1_P2_PHYADDRPOINTER_REG_16_ & n39849;
  assign n39873 = ~P1_P2_PHYADDRPOINTER_REG_17_ & n39872;
  assign n39874 = P1_P2_PHYADDRPOINTER_REG_17_ & ~n39872;
  assign n39875 = ~n39873 & ~n39874;
  assign n39876 = n39498 & ~n39875;
  assign n39877 = P1_P2_PHYADDRPOINTER_REG_16_ & n39854;
  assign n39878 = ~P1_P2_PHYADDRPOINTER_REG_17_ & n39877;
  assign n39879 = P1_P2_PHYADDRPOINTER_REG_17_ & ~n39877;
  assign n39880 = ~n39878 & ~n39879;
  assign n39881 = n39500 & ~n39880;
  assign n39882 = n38385 & n39493;
  assign n39883 = n38393 & n39495;
  assign n39884 = P1_P2_PHYADDRPOINTER_REG_17_ & n39491;
  assign n39885 = P1_P2_REIP_REG_17_ & n39509;
  assign n39886 = n39507 & ~n39880;
  assign n39887 = n38419 & n39504;
  assign n39888 = ~n39884 & ~n39885;
  assign n39889 = ~n39886 & n39888;
  assign n39890 = ~n39887 & n39889;
  assign n39891 = ~n39876 & ~n39881;
  assign n39892 = ~n39882 & n39891;
  assign n39893 = ~n39883 & n39892;
  assign n6796 = ~n39890 | ~n39893;
  assign n39895 = P1_P2_PHYADDRPOINTER_REG_17_ & n39872;
  assign n39896 = ~P1_P2_PHYADDRPOINTER_REG_18_ & n39895;
  assign n39897 = P1_P2_PHYADDRPOINTER_REG_18_ & ~n39895;
  assign n39898 = ~n39896 & ~n39897;
  assign n39899 = n39498 & ~n39898;
  assign n39900 = P1_P2_PHYADDRPOINTER_REG_17_ & n39877;
  assign n39901 = ~P1_P2_PHYADDRPOINTER_REG_18_ & n39900;
  assign n39902 = P1_P2_PHYADDRPOINTER_REG_18_ & ~n39900;
  assign n39903 = ~n39901 & ~n39902;
  assign n39904 = n39500 & ~n39903;
  assign n39905 = ~n38479 & n39493;
  assign n39906 = ~n38492 & n39495;
  assign n39907 = P1_P2_PHYADDRPOINTER_REG_18_ & n39491;
  assign n39908 = P1_P2_REIP_REG_18_ & n39509;
  assign n39909 = n39507 & ~n39903;
  assign n39910 = ~n38463 & n39504;
  assign n39911 = ~n39907 & ~n39908;
  assign n39912 = ~n39909 & n39911;
  assign n39913 = ~n39910 & n39912;
  assign n39914 = ~n39899 & ~n39904;
  assign n39915 = ~n39905 & n39914;
  assign n39916 = ~n39906 & n39915;
  assign n6801 = ~n39913 | ~n39916;
  assign n39918 = P1_P2_PHYADDRPOINTER_REG_18_ & n39895;
  assign n39919 = ~P1_P2_PHYADDRPOINTER_REG_19_ & n39918;
  assign n39920 = P1_P2_PHYADDRPOINTER_REG_19_ & ~n39918;
  assign n39921 = ~n39919 & ~n39920;
  assign n39922 = n39498 & ~n39921;
  assign n39923 = P1_P2_PHYADDRPOINTER_REG_18_ & n39900;
  assign n39924 = ~P1_P2_PHYADDRPOINTER_REG_19_ & n39923;
  assign n39925 = P1_P2_PHYADDRPOINTER_REG_19_ & ~n39923;
  assign n39926 = ~n39924 & ~n39925;
  assign n39927 = n39500 & ~n39926;
  assign n39928 = ~n38533 & n39493;
  assign n39929 = n38542 & n39495;
  assign n39930 = P1_P2_PHYADDRPOINTER_REG_19_ & n39491;
  assign n39931 = P1_P2_REIP_REG_19_ & n39509;
  assign n39932 = n39507 & ~n39926;
  assign n39933 = n38568 & n39504;
  assign n39934 = ~n39930 & ~n39931;
  assign n39935 = ~n39932 & n39934;
  assign n39936 = ~n39933 & n39935;
  assign n39937 = ~n39922 & ~n39927;
  assign n39938 = ~n39928 & n39937;
  assign n39939 = ~n39929 & n39938;
  assign n6806 = ~n39936 | ~n39939;
  assign n39941 = P1_P2_PHYADDRPOINTER_REG_19_ & n39918;
  assign n39942 = ~P1_P2_PHYADDRPOINTER_REG_20_ & n39941;
  assign n39943 = P1_P2_PHYADDRPOINTER_REG_20_ & ~n39941;
  assign n39944 = ~n39942 & ~n39943;
  assign n39945 = n39498 & ~n39944;
  assign n39946 = P1_P2_PHYADDRPOINTER_REG_19_ & n39923;
  assign n39947 = ~P1_P2_PHYADDRPOINTER_REG_20_ & n39946;
  assign n39948 = P1_P2_PHYADDRPOINTER_REG_20_ & ~n39946;
  assign n39949 = ~n39947 & ~n39948;
  assign n39950 = n39500 & ~n39949;
  assign n39951 = n38620 & n39495;
  assign n39952 = P1_P2_PHYADDRPOINTER_REG_20_ & n39491;
  assign n39953 = P1_P2_REIP_REG_20_ & n39509;
  assign n39954 = n39507 & ~n39949;
  assign n39955 = n38644 & n39504;
  assign n39956 = ~n39952 & ~n39953;
  assign n39957 = ~n39954 & n39956;
  assign n39958 = ~n39955 & n39957;
  assign n39959 = n38595 & n39493;
  assign n39960 = ~n39945 & ~n39950;
  assign n39961 = ~n39951 & n39960;
  assign n39962 = n39958 & n39961;
  assign n6811 = n39959 | ~n39962;
  assign n39964 = P1_P2_PHYADDRPOINTER_REG_20_ & n39941;
  assign n39965 = ~P1_P2_PHYADDRPOINTER_REG_21_ & n39964;
  assign n39966 = P1_P2_PHYADDRPOINTER_REG_21_ & ~n39964;
  assign n39967 = ~n39965 & ~n39966;
  assign n39968 = n39498 & ~n39967;
  assign n39969 = P1_P2_PHYADDRPOINTER_REG_20_ & n39946;
  assign n39970 = ~P1_P2_PHYADDRPOINTER_REG_21_ & n39969;
  assign n39971 = P1_P2_PHYADDRPOINTER_REG_21_ & ~n39969;
  assign n39972 = ~n39970 & ~n39971;
  assign n39973 = n39500 & ~n39972;
  assign n39974 = n38677 & n39495;
  assign n39975 = P1_P2_PHYADDRPOINTER_REG_21_ & n39491;
  assign n39976 = P1_P2_REIP_REG_21_ & n39509;
  assign n39977 = n39507 & ~n39972;
  assign n39978 = n38702 & n39504;
  assign n39979 = ~n39975 & ~n39976;
  assign n39980 = ~n39977 & n39979;
  assign n39981 = ~n39978 & n39980;
  assign n39982 = ~n38718 & n39493;
  assign n39983 = ~n39968 & ~n39973;
  assign n39984 = ~n39974 & n39983;
  assign n39985 = n39981 & n39984;
  assign n6816 = n39982 | ~n39985;
  assign n39987 = P1_P2_PHYADDRPOINTER_REG_21_ & n39964;
  assign n39988 = ~P1_P2_PHYADDRPOINTER_REG_22_ & n39987;
  assign n39989 = P1_P2_PHYADDRPOINTER_REG_22_ & ~n39987;
  assign n39990 = ~n39988 & ~n39989;
  assign n39991 = n39498 & ~n39990;
  assign n39992 = ~n38779 & n39493;
  assign n39993 = P1_P2_PHYADDRPOINTER_REG_21_ & n39969;
  assign n39994 = ~P1_P2_PHYADDRPOINTER_REG_22_ & n39993;
  assign n39995 = P1_P2_PHYADDRPOINTER_REG_22_ & ~n39993;
  assign n39996 = ~n39994 & ~n39995;
  assign n39997 = n39500 & ~n39996;
  assign n39998 = ~n38796 & n39495;
  assign n39999 = P1_P2_PHYADDRPOINTER_REG_22_ & n39491;
  assign n40000 = P1_P2_REIP_REG_22_ & n39509;
  assign n40001 = n39507 & ~n39996;
  assign n40002 = ~n38758 & n39504;
  assign n40003 = ~n39999 & ~n40000;
  assign n40004 = ~n40001 & n40003;
  assign n40005 = ~n40002 & n40004;
  assign n40006 = ~n39991 & ~n39992;
  assign n40007 = ~n39997 & n40006;
  assign n40008 = ~n39998 & n40007;
  assign n6821 = ~n40005 | ~n40008;
  assign n40010 = P1_P2_PHYADDRPOINTER_REG_22_ & n39987;
  assign n40011 = ~P1_P2_PHYADDRPOINTER_REG_23_ & n40010;
  assign n40012 = P1_P2_PHYADDRPOINTER_REG_23_ & ~n40010;
  assign n40013 = ~n40011 & ~n40012;
  assign n40014 = n39498 & ~n40013;
  assign n40015 = ~n38855 & n39493;
  assign n40016 = P1_P2_PHYADDRPOINTER_REG_22_ & n39993;
  assign n40017 = ~P1_P2_PHYADDRPOINTER_REG_23_ & n40016;
  assign n40018 = P1_P2_PHYADDRPOINTER_REG_23_ & ~n40016;
  assign n40019 = ~n40017 & ~n40018;
  assign n40020 = n39500 & ~n40019;
  assign n40021 = n38873 & n39495;
  assign n40022 = P1_P2_PHYADDRPOINTER_REG_23_ & n39491;
  assign n40023 = P1_P2_REIP_REG_23_ & n39509;
  assign n40024 = n39507 & ~n40019;
  assign n40025 = n38837 & n39504;
  assign n40026 = ~n40022 & ~n40023;
  assign n40027 = ~n40024 & n40026;
  assign n40028 = ~n40025 & n40027;
  assign n40029 = ~n40014 & ~n40015;
  assign n40030 = ~n40020 & n40029;
  assign n40031 = ~n40021 & n40030;
  assign n6826 = ~n40028 | ~n40031;
  assign n40033 = P1_P2_PHYADDRPOINTER_REG_23_ & n40010;
  assign n40034 = ~P1_P2_PHYADDRPOINTER_REG_24_ & n40033;
  assign n40035 = P1_P2_PHYADDRPOINTER_REG_24_ & ~n40033;
  assign n40036 = ~n40034 & ~n40035;
  assign n40037 = n39498 & ~n40036;
  assign n40038 = ~n38930 & n39493;
  assign n40039 = P1_P2_PHYADDRPOINTER_REG_23_ & n40016;
  assign n40040 = ~P1_P2_PHYADDRPOINTER_REG_24_ & n40039;
  assign n40041 = P1_P2_PHYADDRPOINTER_REG_24_ & ~n40039;
  assign n40042 = ~n40040 & ~n40041;
  assign n40043 = n39500 & ~n40042;
  assign n40044 = ~n38938 & n39495;
  assign n40045 = P1_P2_PHYADDRPOINTER_REG_24_ & n39491;
  assign n40046 = P1_P2_REIP_REG_24_ & n39509;
  assign n40047 = n39507 & ~n40042;
  assign n40048 = ~n38903 & n39504;
  assign n40049 = ~n40045 & ~n40046;
  assign n40050 = ~n40047 & n40049;
  assign n40051 = ~n40048 & n40050;
  assign n40052 = ~n40037 & ~n40038;
  assign n40053 = ~n40043 & n40052;
  assign n40054 = ~n40044 & n40053;
  assign n6831 = ~n40051 | ~n40054;
  assign n40056 = P1_P2_PHYADDRPOINTER_REG_24_ & n40033;
  assign n40057 = ~P1_P2_PHYADDRPOINTER_REG_25_ & n40056;
  assign n40058 = P1_P2_PHYADDRPOINTER_REG_25_ & ~n40056;
  assign n40059 = ~n40057 & ~n40058;
  assign n40060 = n39498 & ~n40059;
  assign n40061 = ~n39007 & n39493;
  assign n40062 = P1_P2_PHYADDRPOINTER_REG_24_ & n40039;
  assign n40063 = ~P1_P2_PHYADDRPOINTER_REG_25_ & n40062;
  assign n40064 = P1_P2_PHYADDRPOINTER_REG_25_ & ~n40062;
  assign n40065 = ~n40063 & ~n40064;
  assign n40066 = n39500 & ~n40065;
  assign n40067 = n39013 & n39495;
  assign n40068 = P1_P2_PHYADDRPOINTER_REG_25_ & n39491;
  assign n40069 = P1_P2_REIP_REG_25_ & n39509;
  assign n40070 = n39507 & ~n40065;
  assign n40071 = n38979 & n39504;
  assign n40072 = ~n40068 & ~n40069;
  assign n40073 = ~n40070 & n40072;
  assign n40074 = ~n40071 & n40073;
  assign n40075 = ~n40060 & ~n40061;
  assign n40076 = ~n40066 & n40075;
  assign n40077 = ~n40067 & n40076;
  assign n6836 = ~n40074 | ~n40077;
  assign n40079 = P1_P2_PHYADDRPOINTER_REG_25_ & n40056;
  assign n40080 = ~P1_P2_PHYADDRPOINTER_REG_26_ & n40079;
  assign n40081 = P1_P2_PHYADDRPOINTER_REG_26_ & ~n40079;
  assign n40082 = ~n40080 & ~n40081;
  assign n40083 = n39498 & ~n40082;
  assign n40084 = n39048 & n39493;
  assign n40085 = P1_P2_PHYADDRPOINTER_REG_25_ & n40062;
  assign n40086 = ~P1_P2_PHYADDRPOINTER_REG_26_ & n40085;
  assign n40087 = P1_P2_PHYADDRPOINTER_REG_26_ & ~n40085;
  assign n40088 = ~n40086 & ~n40087;
  assign n40089 = n39500 & ~n40088;
  assign n40090 = n39052 & n39495;
  assign n40091 = P1_P2_PHYADDRPOINTER_REG_26_ & n39491;
  assign n40092 = n39090 & n39504;
  assign n40093 = n39507 & ~n40088;
  assign n40094 = P1_P2_REIP_REG_26_ & n39509;
  assign n40095 = ~n40091 & ~n40092;
  assign n40096 = ~n40093 & n40095;
  assign n40097 = ~n40094 & n40096;
  assign n40098 = ~n40083 & ~n40084;
  assign n40099 = ~n40089 & n40098;
  assign n40100 = ~n40090 & n40099;
  assign n6841 = ~n40097 | ~n40100;
  assign n40102 = P1_P2_PHYADDRPOINTER_REG_26_ & n40079;
  assign n40103 = ~P1_P2_PHYADDRPOINTER_REG_27_ & n40102;
  assign n40104 = P1_P2_PHYADDRPOINTER_REG_27_ & ~n40102;
  assign n40105 = ~n40103 & ~n40104;
  assign n40106 = n39498 & ~n40105;
  assign n40107 = ~n39119 & n39493;
  assign n40108 = P1_P2_PHYADDRPOINTER_REG_26_ & n40085;
  assign n40109 = ~P1_P2_PHYADDRPOINTER_REG_27_ & n40108;
  assign n40110 = P1_P2_PHYADDRPOINTER_REG_27_ & ~n40108;
  assign n40111 = ~n40109 & ~n40110;
  assign n40112 = n39500 & ~n40111;
  assign n40113 = ~n39123 & n39495;
  assign n40114 = P1_P2_PHYADDRPOINTER_REG_27_ & n39491;
  assign n40115 = ~n39161 & n39504;
  assign n40116 = n39507 & ~n40111;
  assign n40117 = P1_P2_REIP_REG_27_ & n39509;
  assign n40118 = ~n40114 & ~n40115;
  assign n40119 = ~n40116 & n40118;
  assign n40120 = ~n40117 & n40119;
  assign n40121 = ~n40106 & ~n40107;
  assign n40122 = ~n40112 & n40121;
  assign n40123 = ~n40113 & n40122;
  assign n6846 = ~n40120 | ~n40123;
  assign n40125 = n39197 & n39493;
  assign n40126 = n39202 & n39495;
  assign n40127 = P1_P2_PHYADDRPOINTER_REG_27_ & n40102;
  assign n40128 = ~P1_P2_PHYADDRPOINTER_REG_28_ & n40127;
  assign n40129 = P1_P2_PHYADDRPOINTER_REG_28_ & ~n40127;
  assign n40130 = ~n40128 & ~n40129;
  assign n40131 = n39498 & ~n40130;
  assign n40132 = P1_P2_PHYADDRPOINTER_REG_27_ & n40108;
  assign n40133 = ~P1_P2_PHYADDRPOINTER_REG_28_ & n40132;
  assign n40134 = P1_P2_PHYADDRPOINTER_REG_28_ & ~n40132;
  assign n40135 = ~n40133 & ~n40134;
  assign n40136 = n39500 & ~n40135;
  assign n40137 = P1_P2_PHYADDRPOINTER_REG_28_ & n39491;
  assign n40138 = n39241 & n39504;
  assign n40139 = n39507 & ~n40135;
  assign n40140 = P1_P2_REIP_REG_28_ & n39509;
  assign n40141 = ~n40137 & ~n40138;
  assign n40142 = ~n40139 & n40141;
  assign n40143 = ~n40140 & n40142;
  assign n40144 = ~n40125 & ~n40126;
  assign n40145 = ~n40131 & n40144;
  assign n40146 = ~n40136 & n40145;
  assign n6851 = ~n40143 | ~n40146;
  assign n40148 = ~n39270 & n39493;
  assign n40149 = n39274 & n39495;
  assign n40150 = P1_P2_PHYADDRPOINTER_REG_28_ & n40127;
  assign n40151 = ~P1_P2_PHYADDRPOINTER_REG_29_ & n40150;
  assign n40152 = P1_P2_PHYADDRPOINTER_REG_29_ & ~n40150;
  assign n40153 = ~n40151 & ~n40152;
  assign n40154 = n39498 & ~n40153;
  assign n40155 = P1_P2_PHYADDRPOINTER_REG_28_ & n40132;
  assign n40156 = ~P1_P2_PHYADDRPOINTER_REG_29_ & n40155;
  assign n40157 = P1_P2_PHYADDRPOINTER_REG_29_ & ~n40155;
  assign n40158 = ~n40156 & ~n40157;
  assign n40159 = n39500 & ~n40158;
  assign n40160 = P1_P2_PHYADDRPOINTER_REG_29_ & n39491;
  assign n40161 = P1_P2_REIP_REG_29_ & n39509;
  assign n40162 = n39312 & n39504;
  assign n40163 = n39507 & ~n40158;
  assign n40164 = ~n40160 & ~n40161;
  assign n40165 = ~n40162 & n40164;
  assign n40166 = ~n40163 & n40165;
  assign n40167 = ~n40148 & ~n40149;
  assign n40168 = ~n40154 & n40167;
  assign n40169 = ~n40159 & n40168;
  assign n6856 = ~n40166 | ~n40169;
  assign n40171 = ~n39342 & n39493;
  assign n40172 = ~n39346 & n39495;
  assign n40173 = P1_P2_PHYADDRPOINTER_REG_29_ & n40150;
  assign n40174 = ~P1_P2_PHYADDRPOINTER_REG_30_ & n40173;
  assign n40175 = P1_P2_PHYADDRPOINTER_REG_30_ & ~n40173;
  assign n40176 = ~n40174 & ~n40175;
  assign n40177 = n39498 & ~n40176;
  assign n40178 = P1_P2_PHYADDRPOINTER_REG_29_ & n40155;
  assign n40179 = ~P1_P2_PHYADDRPOINTER_REG_30_ & n40178;
  assign n40180 = P1_P2_PHYADDRPOINTER_REG_30_ & ~n40178;
  assign n40181 = ~n40179 & ~n40180;
  assign n40182 = n39500 & ~n40181;
  assign n40183 = P1_P2_PHYADDRPOINTER_REG_30_ & n39491;
  assign n40184 = P1_P2_REIP_REG_30_ & n39509;
  assign n40185 = ~n39384 & n39504;
  assign n40186 = n39507 & ~n40181;
  assign n40187 = ~n40183 & ~n40184;
  assign n40188 = ~n40185 & n40187;
  assign n40189 = ~n40186 & n40188;
  assign n40190 = ~n40171 & ~n40172;
  assign n40191 = ~n40177 & n40190;
  assign n40192 = ~n40182 & n40191;
  assign n6861 = ~n40189 | ~n40192;
  assign n40194 = n39455 & n39493;
  assign n40195 = P1_P2_PHYADDRPOINTER_REG_30_ & n40173;
  assign n40196 = ~P1_P2_PHYADDRPOINTER_REG_31_ & n40195;
  assign n40197 = P1_P2_PHYADDRPOINTER_REG_31_ & ~n40195;
  assign n40198 = ~n40196 & ~n40197;
  assign n40199 = n39498 & ~n40198;
  assign n40200 = ~n39460 & n39495;
  assign n40201 = P1_P2_PHYADDRPOINTER_REG_30_ & n40178;
  assign n40202 = ~P1_P2_PHYADDRPOINTER_REG_31_ & n40201;
  assign n40203 = P1_P2_PHYADDRPOINTER_REG_31_ & ~n40201;
  assign n40204 = ~n40202 & ~n40203;
  assign n40205 = n39500 & ~n40204;
  assign n40206 = P1_P2_PHYADDRPOINTER_REG_31_ & n39491;
  assign n40207 = P1_P2_REIP_REG_31_ & n39509;
  assign n40208 = ~n39408 & n39504;
  assign n40209 = n39507 & ~n40204;
  assign n40210 = ~n40206 & ~n40207;
  assign n40211 = ~n40208 & n40210;
  assign n40212 = ~n40209 & n40211;
  assign n40213 = ~n40194 & ~n40199;
  assign n40214 = ~n40200 & n40213;
  assign n40215 = ~n40205 & n40214;
  assign n6866 = ~n40212 | ~n40215;
  assign n40217 = P1_BUF1_REG_15_ & n12494;
  assign n40218 = P1_BUF2_REG_15_ & ~n12494;
  assign n40219 = ~n40217 & ~n40218;
  assign n40220 = ~n34208 & n34664;
  assign n40221 = n34633 & n40220;
  assign n40222 = ~n34820 & ~n40221;
  assign n40223 = n34935 & ~n40222;
  assign n40224 = ~n34549 & n40223;
  assign n40225 = ~n40219 & n40224;
  assign n40226 = n34549 & n40223;
  assign n40227 = P1_P2_EAX_REG_15_ & n40226;
  assign n40228 = P1_P2_LWORD_REG_15_ & ~n40223;
  assign n40229 = ~n40225 & ~n40227;
  assign n6871 = n40228 | ~n40229;
  assign n40231 = P1_BUF1_REG_14_ & n12494;
  assign n40232 = P1_BUF2_REG_14_ & ~n12494;
  assign n40233 = ~n40231 & ~n40232;
  assign n40234 = n40224 & ~n40233;
  assign n40235 = P1_P2_EAX_REG_14_ & n40226;
  assign n40236 = P1_P2_LWORD_REG_14_ & ~n40223;
  assign n40237 = ~n40234 & ~n40235;
  assign n6876 = n40236 | ~n40237;
  assign n40239 = P1_BUF1_REG_13_ & n12494;
  assign n40240 = P1_BUF2_REG_13_ & ~n12494;
  assign n40241 = ~n40239 & ~n40240;
  assign n40242 = n40224 & ~n40241;
  assign n40243 = P1_P2_EAX_REG_13_ & n40226;
  assign n40244 = P1_P2_LWORD_REG_13_ & ~n40223;
  assign n40245 = ~n40242 & ~n40243;
  assign n6881 = n40244 | ~n40245;
  assign n40247 = P1_BUF1_REG_12_ & n12494;
  assign n40248 = P1_BUF2_REG_12_ & ~n12494;
  assign n40249 = ~n40247 & ~n40248;
  assign n40250 = n40224 & ~n40249;
  assign n40251 = P1_P2_EAX_REG_12_ & n40226;
  assign n40252 = P1_P2_LWORD_REG_12_ & ~n40223;
  assign n40253 = ~n40250 & ~n40251;
  assign n6886 = n40252 | ~n40253;
  assign n40255 = P1_BUF1_REG_11_ & n12494;
  assign n40256 = P1_BUF2_REG_11_ & ~n12494;
  assign n40257 = ~n40255 & ~n40256;
  assign n40258 = n40224 & ~n40257;
  assign n40259 = P1_P2_EAX_REG_11_ & n40226;
  assign n40260 = P1_P2_LWORD_REG_11_ & ~n40223;
  assign n40261 = ~n40258 & ~n40259;
  assign n6891 = n40260 | ~n40261;
  assign n40263 = P1_BUF1_REG_10_ & n12494;
  assign n40264 = P1_BUF2_REG_10_ & ~n12494;
  assign n40265 = ~n40263 & ~n40264;
  assign n40266 = n40224 & ~n40265;
  assign n40267 = P1_P2_EAX_REG_10_ & n40226;
  assign n40268 = P1_P2_LWORD_REG_10_ & ~n40223;
  assign n40269 = ~n40266 & ~n40267;
  assign n6896 = n40268 | ~n40269;
  assign n40271 = P1_BUF1_REG_9_ & n12494;
  assign n40272 = P1_BUF2_REG_9_ & ~n12494;
  assign n40273 = ~n40271 & ~n40272;
  assign n40274 = n40224 & ~n40273;
  assign n40275 = P1_P2_EAX_REG_9_ & n40226;
  assign n40276 = P1_P2_LWORD_REG_9_ & ~n40223;
  assign n40277 = ~n40274 & ~n40275;
  assign n6901 = n40276 | ~n40277;
  assign n40279 = P1_BUF1_REG_8_ & n12494;
  assign n40280 = P1_BUF2_REG_8_ & ~n12494;
  assign n40281 = ~n40279 & ~n40280;
  assign n40282 = n40224 & ~n40281;
  assign n40283 = P1_P2_EAX_REG_8_ & n40226;
  assign n40284 = P1_P2_LWORD_REG_8_ & ~n40223;
  assign n40285 = ~n40282 & ~n40283;
  assign n6906 = n40284 | ~n40285;
  assign n40287 = ~n35072 & n40224;
  assign n40288 = P1_P2_EAX_REG_7_ & n40226;
  assign n40289 = P1_P2_LWORD_REG_7_ & ~n40223;
  assign n40290 = ~n40287 & ~n40288;
  assign n6911 = n40289 | ~n40290;
  assign n40292 = ~n35094 & n40224;
  assign n40293 = P1_P2_EAX_REG_6_ & n40226;
  assign n40294 = P1_P2_LWORD_REG_6_ & ~n40223;
  assign n40295 = ~n40292 & ~n40293;
  assign n6916 = n40294 | ~n40295;
  assign n40297 = ~n35116 & n40224;
  assign n40298 = P1_P2_EAX_REG_5_ & n40226;
  assign n40299 = P1_P2_LWORD_REG_5_ & ~n40223;
  assign n40300 = ~n40297 & ~n40298;
  assign n6921 = n40299 | ~n40300;
  assign n40302 = ~n35138 & n40224;
  assign n40303 = P1_P2_EAX_REG_4_ & n40226;
  assign n40304 = P1_P2_LWORD_REG_4_ & ~n40223;
  assign n40305 = ~n40302 & ~n40303;
  assign n6926 = n40304 | ~n40305;
  assign n40307 = ~n35160 & n40224;
  assign n40308 = P1_P2_EAX_REG_3_ & n40226;
  assign n40309 = P1_P2_LWORD_REG_3_ & ~n40223;
  assign n40310 = ~n40307 & ~n40308;
  assign n6931 = n40309 | ~n40310;
  assign n40312 = ~n35182 & n40224;
  assign n40313 = P1_P2_EAX_REG_2_ & n40226;
  assign n40314 = P1_P2_LWORD_REG_2_ & ~n40223;
  assign n40315 = ~n40312 & ~n40313;
  assign n6936 = n40314 | ~n40315;
  assign n40317 = ~n35204 & n40224;
  assign n40318 = P1_P2_EAX_REG_1_ & n40226;
  assign n40319 = P1_P2_LWORD_REG_1_ & ~n40223;
  assign n40320 = ~n40317 & ~n40318;
  assign n6941 = n40319 | ~n40320;
  assign n40322 = ~n35226 & n40224;
  assign n40323 = P1_P2_EAX_REG_0_ & n40226;
  assign n40324 = P1_P2_LWORD_REG_0_ & ~n40223;
  assign n40325 = ~n40322 & ~n40323;
  assign n6946 = n40324 | ~n40325;
  assign n40327 = P1_P2_EAX_REG_30_ & n40226;
  assign n40328 = P1_P2_UWORD_REG_14_ & ~n40223;
  assign n40329 = ~n40234 & ~n40327;
  assign n6951 = n40328 | ~n40329;
  assign n40331 = P1_P2_EAX_REG_29_ & n40226;
  assign n40332 = P1_P2_UWORD_REG_13_ & ~n40223;
  assign n40333 = ~n40242 & ~n40331;
  assign n6956 = n40332 | ~n40333;
  assign n40335 = P1_P2_EAX_REG_28_ & n40226;
  assign n40336 = P1_P2_UWORD_REG_12_ & ~n40223;
  assign n40337 = ~n40250 & ~n40335;
  assign n6961 = n40336 | ~n40337;
  assign n40339 = P1_P2_EAX_REG_27_ & n40226;
  assign n40340 = P1_P2_UWORD_REG_11_ & ~n40223;
  assign n40341 = ~n40258 & ~n40339;
  assign n6966 = n40340 | ~n40341;
  assign n40343 = P1_P2_EAX_REG_26_ & n40226;
  assign n40344 = P1_P2_UWORD_REG_10_ & ~n40223;
  assign n40345 = ~n40266 & ~n40343;
  assign n6971 = n40344 | ~n40345;
  assign n40347 = P1_P2_EAX_REG_25_ & n40226;
  assign n40348 = P1_P2_UWORD_REG_9_ & ~n40223;
  assign n40349 = ~n40274 & ~n40347;
  assign n6976 = n40348 | ~n40349;
  assign n40351 = P1_P2_EAX_REG_24_ & n40226;
  assign n40352 = P1_P2_UWORD_REG_8_ & ~n40223;
  assign n40353 = ~n40282 & ~n40351;
  assign n6981 = n40352 | ~n40353;
  assign n40355 = P1_P2_EAX_REG_23_ & n40226;
  assign n40356 = P1_P2_UWORD_REG_7_ & ~n40223;
  assign n40357 = ~n40287 & ~n40355;
  assign n6986 = n40356 | ~n40357;
  assign n40359 = P1_P2_EAX_REG_22_ & n40226;
  assign n40360 = P1_P2_UWORD_REG_6_ & ~n40223;
  assign n40361 = ~n40292 & ~n40359;
  assign n6991 = n40360 | ~n40361;
  assign n40363 = P1_P2_EAX_REG_21_ & n40226;
  assign n40364 = P1_P2_UWORD_REG_5_ & ~n40223;
  assign n40365 = ~n40297 & ~n40363;
  assign n6996 = n40364 | ~n40365;
  assign n40367 = P1_P2_EAX_REG_20_ & n40226;
  assign n40368 = P1_P2_UWORD_REG_4_ & ~n40223;
  assign n40369 = ~n40302 & ~n40367;
  assign n7001 = n40368 | ~n40369;
  assign n40371 = P1_P2_EAX_REG_19_ & n40226;
  assign n40372 = P1_P2_UWORD_REG_3_ & ~n40223;
  assign n40373 = ~n40307 & ~n40371;
  assign n7006 = n40372 | ~n40373;
  assign n40375 = P1_P2_EAX_REG_18_ & n40226;
  assign n40376 = P1_P2_UWORD_REG_2_ & ~n40223;
  assign n40377 = ~n40312 & ~n40375;
  assign n7011 = n40376 | ~n40377;
  assign n40379 = P1_P2_EAX_REG_17_ & n40226;
  assign n40380 = P1_P2_UWORD_REG_1_ & ~n40223;
  assign n40381 = ~n40317 & ~n40379;
  assign n7016 = n40380 | ~n40381;
  assign n40383 = P1_P2_EAX_REG_16_ & n40226;
  assign n40384 = P1_P2_UWORD_REG_0_ & ~n40223;
  assign n40385 = ~n40322 & ~n40383;
  assign n7021 = n40384 | ~n40385;
  assign n40387 = ~P1_P2_STATE2_REG_0_ & n34293;
  assign n40388 = n34299 & n34935;
  assign n40389 = ~n34821 & n40388;
  assign n40390 = ~n40387 & ~n40389;
  assign n40391 = P1_P2_STATE2_REG_0_ & ~n40390;
  assign n40392 = P1_P2_EAX_REG_0_ & n40391;
  assign n40393 = ~P1_P2_STATE2_REG_0_ & ~n40390;
  assign n40394 = P1_P2_LWORD_REG_0_ & n40393;
  assign n40395 = P1_P2_DATAO_REG_0_ & n40390;
  assign n40396 = ~n40392 & ~n40394;
  assign n7026 = n40395 | ~n40396;
  assign n40398 = P1_P2_EAX_REG_1_ & n40391;
  assign n40399 = P1_P2_LWORD_REG_1_ & n40393;
  assign n40400 = P1_P2_DATAO_REG_1_ & n40390;
  assign n40401 = ~n40398 & ~n40399;
  assign n7031 = n40400 | ~n40401;
  assign n40403 = P1_P2_EAX_REG_2_ & n40391;
  assign n40404 = P1_P2_LWORD_REG_2_ & n40393;
  assign n40405 = P1_P2_DATAO_REG_2_ & n40390;
  assign n40406 = ~n40403 & ~n40404;
  assign n7036 = n40405 | ~n40406;
  assign n40408 = P1_P2_EAX_REG_3_ & n40391;
  assign n40409 = P1_P2_LWORD_REG_3_ & n40393;
  assign n40410 = P1_P2_DATAO_REG_3_ & n40390;
  assign n40411 = ~n40408 & ~n40409;
  assign n7041 = n40410 | ~n40411;
  assign n40413 = P1_P2_EAX_REG_4_ & n40391;
  assign n40414 = P1_P2_LWORD_REG_4_ & n40393;
  assign n40415 = P1_P2_DATAO_REG_4_ & n40390;
  assign n40416 = ~n40413 & ~n40414;
  assign n7046 = n40415 | ~n40416;
  assign n40418 = P1_P2_EAX_REG_5_ & n40391;
  assign n40419 = P1_P2_LWORD_REG_5_ & n40393;
  assign n40420 = P1_P2_DATAO_REG_5_ & n40390;
  assign n40421 = ~n40418 & ~n40419;
  assign n7051 = n40420 | ~n40421;
  assign n40423 = P1_P2_EAX_REG_6_ & n40391;
  assign n40424 = P1_P2_LWORD_REG_6_ & n40393;
  assign n40425 = P1_P2_DATAO_REG_6_ & n40390;
  assign n40426 = ~n40423 & ~n40424;
  assign n7056 = n40425 | ~n40426;
  assign n40428 = P1_P2_EAX_REG_7_ & n40391;
  assign n40429 = P1_P2_LWORD_REG_7_ & n40393;
  assign n40430 = P1_P2_DATAO_REG_7_ & n40390;
  assign n40431 = ~n40428 & ~n40429;
  assign n7061 = n40430 | ~n40431;
  assign n40433 = P1_P2_EAX_REG_8_ & n40391;
  assign n40434 = P1_P2_LWORD_REG_8_ & n40393;
  assign n40435 = P1_P2_DATAO_REG_8_ & n40390;
  assign n40436 = ~n40433 & ~n40434;
  assign n7066 = n40435 | ~n40436;
  assign n40438 = P1_P2_EAX_REG_9_ & n40391;
  assign n40439 = P1_P2_LWORD_REG_9_ & n40393;
  assign n40440 = P1_P2_DATAO_REG_9_ & n40390;
  assign n40441 = ~n40438 & ~n40439;
  assign n7071 = n40440 | ~n40441;
  assign n40443 = P1_P2_EAX_REG_10_ & n40391;
  assign n40444 = P1_P2_LWORD_REG_10_ & n40393;
  assign n40445 = P1_P2_DATAO_REG_10_ & n40390;
  assign n40446 = ~n40443 & ~n40444;
  assign n7076 = n40445 | ~n40446;
  assign n40448 = P1_P2_EAX_REG_11_ & n40391;
  assign n40449 = P1_P2_LWORD_REG_11_ & n40393;
  assign n40450 = P1_P2_DATAO_REG_11_ & n40390;
  assign n40451 = ~n40448 & ~n40449;
  assign n7081 = n40450 | ~n40451;
  assign n40453 = P1_P2_EAX_REG_12_ & n40391;
  assign n40454 = P1_P2_LWORD_REG_12_ & n40393;
  assign n40455 = P1_P2_DATAO_REG_12_ & n40390;
  assign n40456 = ~n40453 & ~n40454;
  assign n7086 = n40455 | ~n40456;
  assign n40458 = P1_P2_EAX_REG_13_ & n40391;
  assign n40459 = P1_P2_LWORD_REG_13_ & n40393;
  assign n40460 = P1_P2_DATAO_REG_13_ & n40390;
  assign n40461 = ~n40458 & ~n40459;
  assign n7091 = n40460 | ~n40461;
  assign n40463 = P1_P2_EAX_REG_14_ & n40391;
  assign n40464 = P1_P2_LWORD_REG_14_ & n40393;
  assign n40465 = P1_P2_DATAO_REG_14_ & n40390;
  assign n40466 = ~n40463 & ~n40464;
  assign n7096 = n40465 | ~n40466;
  assign n40468 = P1_P2_EAX_REG_15_ & n40391;
  assign n40469 = P1_P2_LWORD_REG_15_ & n40393;
  assign n40470 = P1_P2_DATAO_REG_15_ & n40390;
  assign n40471 = ~n40468 & ~n40469;
  assign n7101 = n40470 | ~n40471;
  assign n40473 = P1_P2_UWORD_REG_0_ & n40393;
  assign n40474 = P1_P2_DATAO_REG_16_ & n40390;
  assign n40475 = ~n40473 & ~n40474;
  assign n40476 = ~n34580 & n40391;
  assign n40477 = P1_P2_EAX_REG_16_ & n40476;
  assign n7106 = ~n40475 | n40477;
  assign n40479 = P1_P2_UWORD_REG_1_ & n40393;
  assign n40480 = P1_P2_DATAO_REG_17_ & n40390;
  assign n40481 = ~n40479 & ~n40480;
  assign n40482 = P1_P2_EAX_REG_17_ & n40476;
  assign n7111 = ~n40481 | n40482;
  assign n40484 = P1_P2_UWORD_REG_2_ & n40393;
  assign n40485 = P1_P2_DATAO_REG_18_ & n40390;
  assign n40486 = ~n40484 & ~n40485;
  assign n40487 = P1_P2_EAX_REG_18_ & n40476;
  assign n7116 = ~n40486 | n40487;
  assign n40489 = P1_P2_UWORD_REG_3_ & n40393;
  assign n40490 = P1_P2_DATAO_REG_19_ & n40390;
  assign n40491 = ~n40489 & ~n40490;
  assign n40492 = P1_P2_EAX_REG_19_ & n40476;
  assign n7121 = ~n40491 | n40492;
  assign n40494 = P1_P2_UWORD_REG_4_ & n40393;
  assign n40495 = P1_P2_DATAO_REG_20_ & n40390;
  assign n40496 = ~n40494 & ~n40495;
  assign n40497 = P1_P2_EAX_REG_20_ & n40476;
  assign n7126 = ~n40496 | n40497;
  assign n40499 = P1_P2_UWORD_REG_5_ & n40393;
  assign n40500 = P1_P2_DATAO_REG_21_ & n40390;
  assign n40501 = ~n40499 & ~n40500;
  assign n40502 = P1_P2_EAX_REG_21_ & n40476;
  assign n7131 = ~n40501 | n40502;
  assign n40504 = P1_P2_UWORD_REG_6_ & n40393;
  assign n40505 = P1_P2_DATAO_REG_22_ & n40390;
  assign n40506 = ~n40504 & ~n40505;
  assign n40507 = P1_P2_EAX_REG_22_ & n40476;
  assign n7136 = ~n40506 | n40507;
  assign n40509 = P1_P2_UWORD_REG_7_ & n40393;
  assign n40510 = P1_P2_DATAO_REG_23_ & n40390;
  assign n40511 = ~n40509 & ~n40510;
  assign n40512 = P1_P2_EAX_REG_23_ & n40476;
  assign n7141 = ~n40511 | n40512;
  assign n40514 = P1_P2_UWORD_REG_8_ & n40393;
  assign n40515 = P1_P2_DATAO_REG_24_ & n40390;
  assign n40516 = ~n40514 & ~n40515;
  assign n40517 = P1_P2_EAX_REG_24_ & n40476;
  assign n7146 = ~n40516 | n40517;
  assign n40519 = P1_P2_UWORD_REG_9_ & n40393;
  assign n40520 = P1_P2_DATAO_REG_25_ & n40390;
  assign n40521 = ~n40519 & ~n40520;
  assign n40522 = P1_P2_EAX_REG_25_ & n40476;
  assign n7151 = ~n40521 | n40522;
  assign n40524 = P1_P2_UWORD_REG_10_ & n40393;
  assign n40525 = P1_P2_DATAO_REG_26_ & n40390;
  assign n40526 = ~n40524 & ~n40525;
  assign n40527 = P1_P2_EAX_REG_26_ & n40476;
  assign n7156 = ~n40526 | n40527;
  assign n40529 = P1_P2_UWORD_REG_11_ & n40393;
  assign n40530 = P1_P2_DATAO_REG_27_ & n40390;
  assign n40531 = ~n40529 & ~n40530;
  assign n40532 = P1_P2_EAX_REG_27_ & n40476;
  assign n7161 = ~n40531 | n40532;
  assign n40534 = P1_P2_UWORD_REG_12_ & n40393;
  assign n40535 = P1_P2_DATAO_REG_28_ & n40390;
  assign n40536 = ~n40534 & ~n40535;
  assign n40537 = P1_P2_EAX_REG_28_ & n40476;
  assign n7166 = ~n40536 | n40537;
  assign n40539 = P1_P2_UWORD_REG_13_ & n40393;
  assign n40540 = P1_P2_DATAO_REG_29_ & n40390;
  assign n40541 = ~n40539 & ~n40540;
  assign n40542 = P1_P2_EAX_REG_29_ & n40476;
  assign n7171 = ~n40541 | n40542;
  assign n40544 = P1_P2_UWORD_REG_14_ & n40393;
  assign n40545 = P1_P2_DATAO_REG_30_ & n40390;
  assign n40546 = ~n40544 & ~n40545;
  assign n40547 = P1_P2_EAX_REG_30_ & n40476;
  assign n7176 = ~n40546 | n40547;
  assign n7181 = P1_P2_DATAO_REG_31_ & n40390;
  assign n40550 = n34815 & ~n34879;
  assign n40551 = n34935 & ~n40550;
  assign n40552 = n34669 & n40551;
  assign n40553 = ~n36717 & n40552;
  assign n40554 = ~n34452 & n40551;
  assign n40555 = ~n34669 & n40554;
  assign n40556 = ~n35226 & n40555;
  assign n40557 = P1_P2_EAX_REG_0_ & ~n40551;
  assign n40558 = n34452 & n40551;
  assign n40559 = ~P1_P2_EAX_REG_0_ & n40558;
  assign n40560 = ~n40557 & ~n40559;
  assign n40561 = ~n40553 & ~n40556;
  assign n7186 = ~n40560 | ~n40561;
  assign n40563 = ~n36835 & n40552;
  assign n40564 = ~n35204 & n40555;
  assign n40565 = P1_P2_EAX_REG_1_ & ~n40551;
  assign n40566 = ~P1_P2_EAX_REG_0_ & P1_P2_EAX_REG_1_;
  assign n40567 = P1_P2_EAX_REG_0_ & ~P1_P2_EAX_REG_1_;
  assign n40568 = ~n40566 & ~n40567;
  assign n40569 = n40558 & ~n40568;
  assign n40570 = ~n40565 & ~n40569;
  assign n40571 = ~n40563 & ~n40564;
  assign n7191 = ~n40570 | ~n40571;
  assign n40573 = ~n36955 & n40552;
  assign n40574 = ~n35182 & n40555;
  assign n40575 = P1_P2_EAX_REG_2_ & ~n40551;
  assign n40576 = P1_P2_EAX_REG_0_ & P1_P2_EAX_REG_1_;
  assign n40577 = ~P1_P2_EAX_REG_2_ & n40576;
  assign n40578 = P1_P2_EAX_REG_2_ & ~n40576;
  assign n40579 = ~n40577 & ~n40578;
  assign n40580 = n40558 & ~n40579;
  assign n40581 = ~n40575 & ~n40580;
  assign n40582 = ~n40573 & ~n40574;
  assign n7196 = ~n40581 | ~n40582;
  assign n40584 = ~n37079 & n40552;
  assign n40585 = ~n35160 & n40555;
  assign n40586 = P1_P2_EAX_REG_3_ & ~n40551;
  assign n40587 = P1_P2_EAX_REG_0_ & P1_P2_EAX_REG_2_;
  assign n40588 = P1_P2_EAX_REG_1_ & n40587;
  assign n40589 = P1_P2_EAX_REG_3_ & ~n40588;
  assign n40590 = ~P1_P2_EAX_REG_3_ & n40588;
  assign n40591 = ~n40589 & ~n40590;
  assign n40592 = n40558 & ~n40591;
  assign n40593 = ~n40586 & ~n40592;
  assign n40594 = ~n40584 & ~n40585;
  assign n7201 = ~n40593 | ~n40594;
  assign n40596 = ~n37206 & n40552;
  assign n40597 = ~n35138 & n40555;
  assign n40598 = P1_P2_EAX_REG_4_ & ~n40551;
  assign n40599 = P1_P2_EAX_REG_3_ & n40588;
  assign n40600 = ~P1_P2_EAX_REG_4_ & n40599;
  assign n40601 = P1_P2_EAX_REG_4_ & ~n40599;
  assign n40602 = ~n40600 & ~n40601;
  assign n40603 = n40558 & ~n40602;
  assign n40604 = ~n40598 & ~n40603;
  assign n40605 = ~n40596 & ~n40597;
  assign n7206 = ~n40604 | ~n40605;
  assign n40607 = ~n37347 & n40552;
  assign n40608 = ~n35116 & n40555;
  assign n40609 = P1_P2_EAX_REG_5_ & ~n40551;
  assign n40610 = P1_P2_EAX_REG_3_ & P1_P2_EAX_REG_4_;
  assign n40611 = n40588 & n40610;
  assign n40612 = P1_P2_EAX_REG_5_ & ~n40611;
  assign n40613 = ~P1_P2_EAX_REG_5_ & n40611;
  assign n40614 = ~n40612 & ~n40613;
  assign n40615 = n40558 & ~n40614;
  assign n40616 = ~n40609 & ~n40615;
  assign n40617 = ~n40607 & ~n40608;
  assign n7211 = ~n40616 | ~n40617;
  assign n40619 = ~n37479 & n40552;
  assign n40620 = ~n35094 & n40555;
  assign n40621 = P1_P2_EAX_REG_6_ & ~n40551;
  assign n40622 = P1_P2_EAX_REG_5_ & n40611;
  assign n40623 = ~P1_P2_EAX_REG_6_ & n40622;
  assign n40624 = P1_P2_EAX_REG_6_ & ~n40622;
  assign n40625 = ~n40623 & ~n40624;
  assign n40626 = n40558 & ~n40625;
  assign n40627 = ~n40621 & ~n40626;
  assign n40628 = ~n40619 & ~n40620;
  assign n7216 = ~n40627 | ~n40628;
  assign n40630 = ~n36751 & n40552;
  assign n40631 = ~n35072 & n40555;
  assign n40632 = P1_P2_EAX_REG_7_ & ~n40551;
  assign n40633 = P1_P2_EAX_REG_5_ & P1_P2_EAX_REG_6_;
  assign n40634 = n40611 & n40633;
  assign n40635 = P1_P2_EAX_REG_7_ & ~n40634;
  assign n40636 = ~P1_P2_EAX_REG_7_ & n40634;
  assign n40637 = ~n40635 & ~n40636;
  assign n40638 = n40558 & ~n40637;
  assign n40639 = ~n40632 & ~n40638;
  assign n40640 = ~n40630 & ~n40631;
  assign n7221 = ~n40639 | ~n40640;
  assign n40642 = ~n34829 & ~n34836;
  assign n40643 = ~n34780 & ~n40642;
  assign n40644 = n34310 & n40643;
  assign n40645 = P1_P2_INSTQUEUE_REG_15__0_ & n40644;
  assign n40646 = n34314 & n40643;
  assign n40647 = P1_P2_INSTQUEUE_REG_14__0_ & n40646;
  assign n40648 = n34301 & n40643;
  assign n40649 = P1_P2_INSTQUEUE_REG_13__0_ & n40648;
  assign n40650 = n34305 & n40643;
  assign n40651 = P1_P2_INSTQUEUE_REG_12__0_ & n40650;
  assign n40652 = ~n40645 & ~n40647;
  assign n40653 = ~n40649 & n40652;
  assign n40654 = ~n40651 & n40653;
  assign n40655 = n34780 & ~n40642;
  assign n40656 = n34310 & n40655;
  assign n40657 = P1_P2_INSTQUEUE_REG_11__0_ & n40656;
  assign n40658 = n34314 & n40655;
  assign n40659 = P1_P2_INSTQUEUE_REG_10__0_ & n40658;
  assign n40660 = n34301 & n40655;
  assign n40661 = P1_P2_INSTQUEUE_REG_9__0_ & n40660;
  assign n40662 = n34305 & n40655;
  assign n40663 = P1_P2_INSTQUEUE_REG_8__0_ & n40662;
  assign n40664 = ~n40657 & ~n40659;
  assign n40665 = ~n40661 & n40664;
  assign n40666 = ~n40663 & n40665;
  assign n40667 = ~n34780 & n40642;
  assign n40668 = n34310 & n40667;
  assign n40669 = P1_P2_INSTQUEUE_REG_7__0_ & n40668;
  assign n40670 = n34314 & n40667;
  assign n40671 = P1_P2_INSTQUEUE_REG_6__0_ & n40670;
  assign n40672 = n34301 & n40667;
  assign n40673 = P1_P2_INSTQUEUE_REG_5__0_ & n40672;
  assign n40674 = n34305 & n40667;
  assign n40675 = P1_P2_INSTQUEUE_REG_4__0_ & n40674;
  assign n40676 = ~n40669 & ~n40671;
  assign n40677 = ~n40673 & n40676;
  assign n40678 = ~n40675 & n40677;
  assign n40679 = n34780 & n40642;
  assign n40680 = n34310 & n40679;
  assign n40681 = P1_P2_INSTQUEUE_REG_3__0_ & n40680;
  assign n40682 = n34314 & n40679;
  assign n40683 = P1_P2_INSTQUEUE_REG_2__0_ & n40682;
  assign n40684 = n34301 & n40679;
  assign n40685 = P1_P2_INSTQUEUE_REG_1__0_ & n40684;
  assign n40686 = n34305 & n40679;
  assign n40687 = P1_P2_INSTQUEUE_REG_0__0_ & n40686;
  assign n40688 = ~n40681 & ~n40683;
  assign n40689 = ~n40685 & n40688;
  assign n40690 = ~n40687 & n40689;
  assign n40691 = n40654 & n40666;
  assign n40692 = n40678 & n40691;
  assign n40693 = n40690 & n40692;
  assign n40694 = n40552 & ~n40693;
  assign n40695 = ~n40281 & n40555;
  assign n40696 = P1_P2_EAX_REG_8_ & ~n40551;
  assign n40697 = P1_P2_EAX_REG_7_ & n40634;
  assign n40698 = ~P1_P2_EAX_REG_8_ & n40697;
  assign n40699 = P1_P2_EAX_REG_8_ & ~n40697;
  assign n40700 = ~n40698 & ~n40699;
  assign n40701 = n40558 & ~n40700;
  assign n40702 = ~n40696 & ~n40701;
  assign n40703 = ~n40694 & ~n40695;
  assign n7226 = ~n40702 | ~n40703;
  assign n40705 = P1_P2_INSTQUEUE_REG_15__1_ & n40644;
  assign n40706 = P1_P2_INSTQUEUE_REG_14__1_ & n40646;
  assign n40707 = P1_P2_INSTQUEUE_REG_13__1_ & n40648;
  assign n40708 = P1_P2_INSTQUEUE_REG_12__1_ & n40650;
  assign n40709 = ~n40705 & ~n40706;
  assign n40710 = ~n40707 & n40709;
  assign n40711 = ~n40708 & n40710;
  assign n40712 = P1_P2_INSTQUEUE_REG_11__1_ & n40656;
  assign n40713 = P1_P2_INSTQUEUE_REG_10__1_ & n40658;
  assign n40714 = P1_P2_INSTQUEUE_REG_9__1_ & n40660;
  assign n40715 = P1_P2_INSTQUEUE_REG_8__1_ & n40662;
  assign n40716 = ~n40712 & ~n40713;
  assign n40717 = ~n40714 & n40716;
  assign n40718 = ~n40715 & n40717;
  assign n40719 = P1_P2_INSTQUEUE_REG_7__1_ & n40668;
  assign n40720 = P1_P2_INSTQUEUE_REG_6__1_ & n40670;
  assign n40721 = P1_P2_INSTQUEUE_REG_5__1_ & n40672;
  assign n40722 = P1_P2_INSTQUEUE_REG_4__1_ & n40674;
  assign n40723 = ~n40719 & ~n40720;
  assign n40724 = ~n40721 & n40723;
  assign n40725 = ~n40722 & n40724;
  assign n40726 = P1_P2_INSTQUEUE_REG_3__1_ & n40680;
  assign n40727 = P1_P2_INSTQUEUE_REG_2__1_ & n40682;
  assign n40728 = P1_P2_INSTQUEUE_REG_1__1_ & n40684;
  assign n40729 = P1_P2_INSTQUEUE_REG_0__1_ & n40686;
  assign n40730 = ~n40726 & ~n40727;
  assign n40731 = ~n40728 & n40730;
  assign n40732 = ~n40729 & n40731;
  assign n40733 = n40711 & n40718;
  assign n40734 = n40725 & n40733;
  assign n40735 = n40732 & n40734;
  assign n40736 = n40552 & ~n40735;
  assign n40737 = ~n40273 & n40555;
  assign n40738 = P1_P2_EAX_REG_9_ & ~n40551;
  assign n40739 = P1_P2_EAX_REG_7_ & P1_P2_EAX_REG_8_;
  assign n40740 = n40634 & n40739;
  assign n40741 = P1_P2_EAX_REG_9_ & ~n40740;
  assign n40742 = ~P1_P2_EAX_REG_9_ & n40740;
  assign n40743 = ~n40741 & ~n40742;
  assign n40744 = n40558 & ~n40743;
  assign n40745 = ~n40738 & ~n40744;
  assign n40746 = ~n40736 & ~n40737;
  assign n7231 = ~n40745 | ~n40746;
  assign n40748 = P1_P2_INSTQUEUE_REG_15__2_ & n40644;
  assign n40749 = P1_P2_INSTQUEUE_REG_14__2_ & n40646;
  assign n40750 = P1_P2_INSTQUEUE_REG_13__2_ & n40648;
  assign n40751 = P1_P2_INSTQUEUE_REG_12__2_ & n40650;
  assign n40752 = ~n40748 & ~n40749;
  assign n40753 = ~n40750 & n40752;
  assign n40754 = ~n40751 & n40753;
  assign n40755 = P1_P2_INSTQUEUE_REG_11__2_ & n40656;
  assign n40756 = P1_P2_INSTQUEUE_REG_10__2_ & n40658;
  assign n40757 = P1_P2_INSTQUEUE_REG_9__2_ & n40660;
  assign n40758 = P1_P2_INSTQUEUE_REG_8__2_ & n40662;
  assign n40759 = ~n40755 & ~n40756;
  assign n40760 = ~n40757 & n40759;
  assign n40761 = ~n40758 & n40760;
  assign n40762 = P1_P2_INSTQUEUE_REG_7__2_ & n40668;
  assign n40763 = P1_P2_INSTQUEUE_REG_6__2_ & n40670;
  assign n40764 = P1_P2_INSTQUEUE_REG_5__2_ & n40672;
  assign n40765 = P1_P2_INSTQUEUE_REG_4__2_ & n40674;
  assign n40766 = ~n40762 & ~n40763;
  assign n40767 = ~n40764 & n40766;
  assign n40768 = ~n40765 & n40767;
  assign n40769 = P1_P2_INSTQUEUE_REG_3__2_ & n40680;
  assign n40770 = P1_P2_INSTQUEUE_REG_2__2_ & n40682;
  assign n40771 = P1_P2_INSTQUEUE_REG_1__2_ & n40684;
  assign n40772 = P1_P2_INSTQUEUE_REG_0__2_ & n40686;
  assign n40773 = ~n40769 & ~n40770;
  assign n40774 = ~n40771 & n40773;
  assign n40775 = ~n40772 & n40774;
  assign n40776 = n40754 & n40761;
  assign n40777 = n40768 & n40776;
  assign n40778 = n40775 & n40777;
  assign n40779 = n40552 & ~n40778;
  assign n40780 = ~n40265 & n40555;
  assign n40781 = P1_P2_EAX_REG_10_ & ~n40551;
  assign n40782 = P1_P2_EAX_REG_9_ & n40740;
  assign n40783 = ~P1_P2_EAX_REG_10_ & n40782;
  assign n40784 = P1_P2_EAX_REG_10_ & ~n40782;
  assign n40785 = ~n40783 & ~n40784;
  assign n40786 = n40558 & ~n40785;
  assign n40787 = ~n40781 & ~n40786;
  assign n40788 = ~n40779 & ~n40780;
  assign n7236 = ~n40787 | ~n40788;
  assign n40790 = P1_P2_INSTQUEUE_REG_15__3_ & n40644;
  assign n40791 = P1_P2_INSTQUEUE_REG_14__3_ & n40646;
  assign n40792 = P1_P2_INSTQUEUE_REG_13__3_ & n40648;
  assign n40793 = P1_P2_INSTQUEUE_REG_12__3_ & n40650;
  assign n40794 = ~n40790 & ~n40791;
  assign n40795 = ~n40792 & n40794;
  assign n40796 = ~n40793 & n40795;
  assign n40797 = P1_P2_INSTQUEUE_REG_11__3_ & n40656;
  assign n40798 = P1_P2_INSTQUEUE_REG_10__3_ & n40658;
  assign n40799 = P1_P2_INSTQUEUE_REG_9__3_ & n40660;
  assign n40800 = P1_P2_INSTQUEUE_REG_8__3_ & n40662;
  assign n40801 = ~n40797 & ~n40798;
  assign n40802 = ~n40799 & n40801;
  assign n40803 = ~n40800 & n40802;
  assign n40804 = P1_P2_INSTQUEUE_REG_7__3_ & n40668;
  assign n40805 = P1_P2_INSTQUEUE_REG_6__3_ & n40670;
  assign n40806 = P1_P2_INSTQUEUE_REG_5__3_ & n40672;
  assign n40807 = P1_P2_INSTQUEUE_REG_4__3_ & n40674;
  assign n40808 = ~n40804 & ~n40805;
  assign n40809 = ~n40806 & n40808;
  assign n40810 = ~n40807 & n40809;
  assign n40811 = P1_P2_INSTQUEUE_REG_3__3_ & n40680;
  assign n40812 = P1_P2_INSTQUEUE_REG_2__3_ & n40682;
  assign n40813 = P1_P2_INSTQUEUE_REG_1__3_ & n40684;
  assign n40814 = P1_P2_INSTQUEUE_REG_0__3_ & n40686;
  assign n40815 = ~n40811 & ~n40812;
  assign n40816 = ~n40813 & n40815;
  assign n40817 = ~n40814 & n40816;
  assign n40818 = n40796 & n40803;
  assign n40819 = n40810 & n40818;
  assign n40820 = n40817 & n40819;
  assign n40821 = n40552 & ~n40820;
  assign n40822 = ~n40257 & n40555;
  assign n40823 = P1_P2_EAX_REG_11_ & ~n40551;
  assign n40824 = P1_P2_EAX_REG_9_ & P1_P2_EAX_REG_10_;
  assign n40825 = n40740 & n40824;
  assign n40826 = P1_P2_EAX_REG_11_ & ~n40825;
  assign n40827 = ~P1_P2_EAX_REG_11_ & n40825;
  assign n40828 = ~n40826 & ~n40827;
  assign n40829 = n40558 & ~n40828;
  assign n40830 = ~n40823 & ~n40829;
  assign n40831 = ~n40821 & ~n40822;
  assign n7241 = ~n40830 | ~n40831;
  assign n40833 = P1_P2_INSTQUEUE_REG_15__4_ & n40644;
  assign n40834 = P1_P2_INSTQUEUE_REG_14__4_ & n40646;
  assign n40835 = P1_P2_INSTQUEUE_REG_13__4_ & n40648;
  assign n40836 = P1_P2_INSTQUEUE_REG_12__4_ & n40650;
  assign n40837 = ~n40833 & ~n40834;
  assign n40838 = ~n40835 & n40837;
  assign n40839 = ~n40836 & n40838;
  assign n40840 = P1_P2_INSTQUEUE_REG_11__4_ & n40656;
  assign n40841 = P1_P2_INSTQUEUE_REG_10__4_ & n40658;
  assign n40842 = P1_P2_INSTQUEUE_REG_9__4_ & n40660;
  assign n40843 = P1_P2_INSTQUEUE_REG_8__4_ & n40662;
  assign n40844 = ~n40840 & ~n40841;
  assign n40845 = ~n40842 & n40844;
  assign n40846 = ~n40843 & n40845;
  assign n40847 = P1_P2_INSTQUEUE_REG_7__4_ & n40668;
  assign n40848 = P1_P2_INSTQUEUE_REG_6__4_ & n40670;
  assign n40849 = P1_P2_INSTQUEUE_REG_5__4_ & n40672;
  assign n40850 = P1_P2_INSTQUEUE_REG_4__4_ & n40674;
  assign n40851 = ~n40847 & ~n40848;
  assign n40852 = ~n40849 & n40851;
  assign n40853 = ~n40850 & n40852;
  assign n40854 = P1_P2_INSTQUEUE_REG_3__4_ & n40680;
  assign n40855 = P1_P2_INSTQUEUE_REG_2__4_ & n40682;
  assign n40856 = P1_P2_INSTQUEUE_REG_1__4_ & n40684;
  assign n40857 = P1_P2_INSTQUEUE_REG_0__4_ & n40686;
  assign n40858 = ~n40854 & ~n40855;
  assign n40859 = ~n40856 & n40858;
  assign n40860 = ~n40857 & n40859;
  assign n40861 = n40839 & n40846;
  assign n40862 = n40853 & n40861;
  assign n40863 = n40860 & n40862;
  assign n40864 = n40552 & ~n40863;
  assign n40865 = ~n40249 & n40555;
  assign n40866 = P1_P2_EAX_REG_12_ & ~n40551;
  assign n40867 = P1_P2_EAX_REG_11_ & n40825;
  assign n40868 = ~P1_P2_EAX_REG_12_ & n40867;
  assign n40869 = P1_P2_EAX_REG_12_ & ~n40867;
  assign n40870 = ~n40868 & ~n40869;
  assign n40871 = n40558 & ~n40870;
  assign n40872 = ~n40866 & ~n40871;
  assign n40873 = ~n40864 & ~n40865;
  assign n7246 = ~n40872 | ~n40873;
  assign n40875 = ~n40241 & n40555;
  assign n40876 = P1_P2_INSTQUEUE_REG_15__5_ & n40644;
  assign n40877 = P1_P2_INSTQUEUE_REG_14__5_ & n40646;
  assign n40878 = P1_P2_INSTQUEUE_REG_13__5_ & n40648;
  assign n40879 = P1_P2_INSTQUEUE_REG_12__5_ & n40650;
  assign n40880 = ~n40876 & ~n40877;
  assign n40881 = ~n40878 & n40880;
  assign n40882 = ~n40879 & n40881;
  assign n40883 = P1_P2_INSTQUEUE_REG_11__5_ & n40656;
  assign n40884 = P1_P2_INSTQUEUE_REG_10__5_ & n40658;
  assign n40885 = P1_P2_INSTQUEUE_REG_9__5_ & n40660;
  assign n40886 = P1_P2_INSTQUEUE_REG_8__5_ & n40662;
  assign n40887 = ~n40883 & ~n40884;
  assign n40888 = ~n40885 & n40887;
  assign n40889 = ~n40886 & n40888;
  assign n40890 = P1_P2_INSTQUEUE_REG_7__5_ & n40668;
  assign n40891 = P1_P2_INSTQUEUE_REG_6__5_ & n40670;
  assign n40892 = P1_P2_INSTQUEUE_REG_5__5_ & n40672;
  assign n40893 = P1_P2_INSTQUEUE_REG_4__5_ & n40674;
  assign n40894 = ~n40890 & ~n40891;
  assign n40895 = ~n40892 & n40894;
  assign n40896 = ~n40893 & n40895;
  assign n40897 = P1_P2_INSTQUEUE_REG_3__5_ & n40680;
  assign n40898 = P1_P2_INSTQUEUE_REG_2__5_ & n40682;
  assign n40899 = P1_P2_INSTQUEUE_REG_1__5_ & n40684;
  assign n40900 = P1_P2_INSTQUEUE_REG_0__5_ & n40686;
  assign n40901 = ~n40897 & ~n40898;
  assign n40902 = ~n40899 & n40901;
  assign n40903 = ~n40900 & n40902;
  assign n40904 = n40882 & n40889;
  assign n40905 = n40896 & n40904;
  assign n40906 = n40903 & n40905;
  assign n40907 = n40552 & ~n40906;
  assign n40908 = P1_P2_EAX_REG_13_ & ~n40551;
  assign n40909 = ~n40907 & ~n40908;
  assign n40910 = P1_P2_EAX_REG_11_ & P1_P2_EAX_REG_12_;
  assign n40911 = n40825 & n40910;
  assign n40912 = P1_P2_EAX_REG_13_ & ~n40911;
  assign n40913 = ~P1_P2_EAX_REG_13_ & n40911;
  assign n40914 = ~n40912 & ~n40913;
  assign n40915 = n40558 & ~n40914;
  assign n40916 = ~n40875 & n40909;
  assign n7251 = n40915 | ~n40916;
  assign n40918 = ~n40233 & n40555;
  assign n40919 = P1_P2_INSTQUEUE_REG_15__6_ & n40644;
  assign n40920 = P1_P2_INSTQUEUE_REG_14__6_ & n40646;
  assign n40921 = P1_P2_INSTQUEUE_REG_13__6_ & n40648;
  assign n40922 = P1_P2_INSTQUEUE_REG_12__6_ & n40650;
  assign n40923 = ~n40919 & ~n40920;
  assign n40924 = ~n40921 & n40923;
  assign n40925 = ~n40922 & n40924;
  assign n40926 = P1_P2_INSTQUEUE_REG_11__6_ & n40656;
  assign n40927 = P1_P2_INSTQUEUE_REG_10__6_ & n40658;
  assign n40928 = P1_P2_INSTQUEUE_REG_9__6_ & n40660;
  assign n40929 = P1_P2_INSTQUEUE_REG_8__6_ & n40662;
  assign n40930 = ~n40926 & ~n40927;
  assign n40931 = ~n40928 & n40930;
  assign n40932 = ~n40929 & n40931;
  assign n40933 = P1_P2_INSTQUEUE_REG_7__6_ & n40668;
  assign n40934 = P1_P2_INSTQUEUE_REG_6__6_ & n40670;
  assign n40935 = P1_P2_INSTQUEUE_REG_5__6_ & n40672;
  assign n40936 = P1_P2_INSTQUEUE_REG_4__6_ & n40674;
  assign n40937 = ~n40933 & ~n40934;
  assign n40938 = ~n40935 & n40937;
  assign n40939 = ~n40936 & n40938;
  assign n40940 = P1_P2_INSTQUEUE_REG_3__6_ & n40680;
  assign n40941 = P1_P2_INSTQUEUE_REG_2__6_ & n40682;
  assign n40942 = P1_P2_INSTQUEUE_REG_1__6_ & n40684;
  assign n40943 = P1_P2_INSTQUEUE_REG_0__6_ & n40686;
  assign n40944 = ~n40940 & ~n40941;
  assign n40945 = ~n40942 & n40944;
  assign n40946 = ~n40943 & n40945;
  assign n40947 = n40925 & n40932;
  assign n40948 = n40939 & n40947;
  assign n40949 = n40946 & n40948;
  assign n40950 = n40552 & ~n40949;
  assign n40951 = P1_P2_EAX_REG_14_ & ~n40551;
  assign n40952 = ~n40950 & ~n40951;
  assign n40953 = P1_P2_EAX_REG_13_ & n40911;
  assign n40954 = ~P1_P2_EAX_REG_14_ & n40953;
  assign n40955 = P1_P2_EAX_REG_14_ & ~n40953;
  assign n40956 = ~n40954 & ~n40955;
  assign n40957 = n40558 & ~n40956;
  assign n40958 = ~n40918 & n40952;
  assign n7256 = n40957 | ~n40958;
  assign n40960 = ~n40219 & n40555;
  assign n40961 = P1_P2_INSTQUEUE_REG_15__7_ & n40644;
  assign n40962 = P1_P2_INSTQUEUE_REG_14__7_ & n40646;
  assign n40963 = P1_P2_INSTQUEUE_REG_13__7_ & n40648;
  assign n40964 = P1_P2_INSTQUEUE_REG_12__7_ & n40650;
  assign n40965 = ~n40961 & ~n40962;
  assign n40966 = ~n40963 & n40965;
  assign n40967 = ~n40964 & n40966;
  assign n40968 = P1_P2_INSTQUEUE_REG_11__7_ & n40656;
  assign n40969 = P1_P2_INSTQUEUE_REG_10__7_ & n40658;
  assign n40970 = P1_P2_INSTQUEUE_REG_9__7_ & n40660;
  assign n40971 = P1_P2_INSTQUEUE_REG_8__7_ & n40662;
  assign n40972 = ~n40968 & ~n40969;
  assign n40973 = ~n40970 & n40972;
  assign n40974 = ~n40971 & n40973;
  assign n40975 = P1_P2_INSTQUEUE_REG_7__7_ & n40668;
  assign n40976 = P1_P2_INSTQUEUE_REG_6__7_ & n40670;
  assign n40977 = P1_P2_INSTQUEUE_REG_5__7_ & n40672;
  assign n40978 = P1_P2_INSTQUEUE_REG_4__7_ & n40674;
  assign n40979 = ~n40975 & ~n40976;
  assign n40980 = ~n40977 & n40979;
  assign n40981 = ~n40978 & n40980;
  assign n40982 = P1_P2_INSTQUEUE_REG_3__7_ & n40680;
  assign n40983 = P1_P2_INSTQUEUE_REG_2__7_ & n40682;
  assign n40984 = P1_P2_INSTQUEUE_REG_1__7_ & n40684;
  assign n40985 = P1_P2_INSTQUEUE_REG_0__7_ & n40686;
  assign n40986 = ~n40982 & ~n40983;
  assign n40987 = ~n40984 & n40986;
  assign n40988 = ~n40985 & n40987;
  assign n40989 = n40967 & n40974;
  assign n40990 = n40981 & n40989;
  assign n40991 = n40988 & n40990;
  assign n40992 = n40552 & ~n40991;
  assign n40993 = P1_P2_EAX_REG_15_ & ~n40551;
  assign n40994 = ~n40992 & ~n40993;
  assign n40995 = P1_P2_EAX_REG_13_ & P1_P2_EAX_REG_14_;
  assign n40996 = n40911 & n40995;
  assign n40997 = P1_P2_EAX_REG_15_ & ~n40996;
  assign n40998 = ~P1_P2_EAX_REG_15_ & n40996;
  assign n40999 = ~n40997 & ~n40998;
  assign n41000 = n40558 & ~n40999;
  assign n41001 = ~n40960 & n40994;
  assign n7261 = n41000 | ~n41001;
  assign n41003 = ~n34389 & n40554;
  assign n41004 = ~n35212 & n41003;
  assign n41005 = n34358 & n40554;
  assign n41006 = ~n35226 & n41005;
  assign n41007 = P1_P2_EAX_REG_16_ & ~n40551;
  assign n41008 = P1_P2_INSTQUEUERD_ADDR_REG_2_ & ~n34314;
  assign n41009 = ~P1_P2_INSTQUEUERD_ADDR_REG_3_ & n41008;
  assign n41010 = P1_P2_INSTQUEUERD_ADDR_REG_3_ & ~n41008;
  assign n41011 = ~n41009 & ~n41010;
  assign n41012 = ~n34315 & ~n41008;
  assign n41013 = n41011 & n41012;
  assign n41014 = n36667 & n41013;
  assign n41015 = P1_P2_INSTQUEUE_REG_7__0_ & n41014;
  assign n41016 = n36664 & n41013;
  assign n41017 = P1_P2_INSTQUEUE_REG_6__0_ & n41016;
  assign n41018 = n36673 & n41013;
  assign n41019 = P1_P2_INSTQUEUE_REG_5__0_ & n41018;
  assign n41020 = n36670 & n41013;
  assign n41021 = P1_P2_INSTQUEUE_REG_4__0_ & n41020;
  assign n41022 = ~n41015 & ~n41017;
  assign n41023 = ~n41019 & n41022;
  assign n41024 = ~n41021 & n41023;
  assign n41025 = n41011 & ~n41012;
  assign n41026 = n36667 & n41025;
  assign n41027 = P1_P2_INSTQUEUE_REG_3__0_ & n41026;
  assign n41028 = n36664 & n41025;
  assign n41029 = P1_P2_INSTQUEUE_REG_2__0_ & n41028;
  assign n41030 = n36673 & n41025;
  assign n41031 = P1_P2_INSTQUEUE_REG_1__0_ & n41030;
  assign n41032 = n36670 & n41025;
  assign n41033 = P1_P2_INSTQUEUE_REG_0__0_ & n41032;
  assign n41034 = ~n41027 & ~n41029;
  assign n41035 = ~n41031 & n41034;
  assign n41036 = ~n41033 & n41035;
  assign n41037 = ~n41011 & n41012;
  assign n41038 = n36667 & n41037;
  assign n41039 = P1_P2_INSTQUEUE_REG_15__0_ & n41038;
  assign n41040 = n36664 & n41037;
  assign n41041 = P1_P2_INSTQUEUE_REG_14__0_ & n41040;
  assign n41042 = n36673 & n41037;
  assign n41043 = P1_P2_INSTQUEUE_REG_13__0_ & n41042;
  assign n41044 = n36670 & n41037;
  assign n41045 = P1_P2_INSTQUEUE_REG_12__0_ & n41044;
  assign n41046 = ~n41039 & ~n41041;
  assign n41047 = ~n41043 & n41046;
  assign n41048 = ~n41045 & n41047;
  assign n41049 = ~n41011 & ~n41012;
  assign n41050 = n36667 & n41049;
  assign n41051 = P1_P2_INSTQUEUE_REG_11__0_ & n41050;
  assign n41052 = n36664 & n41049;
  assign n41053 = P1_P2_INSTQUEUE_REG_10__0_ & n41052;
  assign n41054 = n36673 & n41049;
  assign n41055 = P1_P2_INSTQUEUE_REG_9__0_ & n41054;
  assign n41056 = n36670 & n41049;
  assign n41057 = P1_P2_INSTQUEUE_REG_8__0_ & n41056;
  assign n41058 = ~n41051 & ~n41053;
  assign n41059 = ~n41055 & n41058;
  assign n41060 = ~n41057 & n41059;
  assign n41061 = n41024 & n41036;
  assign n41062 = n41048 & n41061;
  assign n41063 = n41060 & n41062;
  assign n41064 = n40552 & ~n41063;
  assign n41065 = ~n41007 & ~n41064;
  assign n41066 = P1_P2_EAX_REG_15_ & n40996;
  assign n41067 = ~P1_P2_EAX_REG_16_ & n41066;
  assign n41068 = P1_P2_EAX_REG_16_ & ~n41066;
  assign n41069 = ~n41067 & ~n41068;
  assign n41070 = n40558 & ~n41069;
  assign n41071 = ~n41004 & ~n41006;
  assign n41072 = n41065 & n41071;
  assign n7266 = n41070 | ~n41072;
  assign n41074 = ~n35190 & n41003;
  assign n41075 = ~n35204 & n41005;
  assign n41076 = P1_P2_EAX_REG_17_ & ~n40551;
  assign n41077 = P1_P2_INSTQUEUE_REG_7__1_ & n41014;
  assign n41078 = P1_P2_INSTQUEUE_REG_6__1_ & n41016;
  assign n41079 = P1_P2_INSTQUEUE_REG_5__1_ & n41018;
  assign n41080 = P1_P2_INSTQUEUE_REG_4__1_ & n41020;
  assign n41081 = ~n41077 & ~n41078;
  assign n41082 = ~n41079 & n41081;
  assign n41083 = ~n41080 & n41082;
  assign n41084 = P1_P2_INSTQUEUE_REG_3__1_ & n41026;
  assign n41085 = P1_P2_INSTQUEUE_REG_2__1_ & n41028;
  assign n41086 = P1_P2_INSTQUEUE_REG_1__1_ & n41030;
  assign n41087 = P1_P2_INSTQUEUE_REG_0__1_ & n41032;
  assign n41088 = ~n41084 & ~n41085;
  assign n41089 = ~n41086 & n41088;
  assign n41090 = ~n41087 & n41089;
  assign n41091 = P1_P2_INSTQUEUE_REG_15__1_ & n41038;
  assign n41092 = P1_P2_INSTQUEUE_REG_14__1_ & n41040;
  assign n41093 = P1_P2_INSTQUEUE_REG_13__1_ & n41042;
  assign n41094 = P1_P2_INSTQUEUE_REG_12__1_ & n41044;
  assign n41095 = ~n41091 & ~n41092;
  assign n41096 = ~n41093 & n41095;
  assign n41097 = ~n41094 & n41096;
  assign n41098 = P1_P2_INSTQUEUE_REG_11__1_ & n41050;
  assign n41099 = P1_P2_INSTQUEUE_REG_10__1_ & n41052;
  assign n41100 = P1_P2_INSTQUEUE_REG_9__1_ & n41054;
  assign n41101 = P1_P2_INSTQUEUE_REG_8__1_ & n41056;
  assign n41102 = ~n41098 & ~n41099;
  assign n41103 = ~n41100 & n41102;
  assign n41104 = ~n41101 & n41103;
  assign n41105 = n41083 & n41090;
  assign n41106 = n41097 & n41105;
  assign n41107 = n41104 & n41106;
  assign n41108 = n40552 & ~n41107;
  assign n41109 = ~n41076 & ~n41108;
  assign n41110 = P1_P2_EAX_REG_15_ & P1_P2_EAX_REG_16_;
  assign n41111 = n40996 & n41110;
  assign n41112 = P1_P2_EAX_REG_17_ & ~n41111;
  assign n41113 = ~P1_P2_EAX_REG_17_ & n41111;
  assign n41114 = ~n41112 & ~n41113;
  assign n41115 = n40558 & ~n41114;
  assign n41116 = ~n41074 & ~n41075;
  assign n41117 = n41109 & n41116;
  assign n7271 = n41115 | ~n41117;
  assign n41119 = ~n35168 & n41003;
  assign n41120 = ~n35182 & n41005;
  assign n41121 = P1_P2_EAX_REG_18_ & ~n40551;
  assign n41122 = P1_P2_INSTQUEUE_REG_7__2_ & n41014;
  assign n41123 = P1_P2_INSTQUEUE_REG_6__2_ & n41016;
  assign n41124 = P1_P2_INSTQUEUE_REG_5__2_ & n41018;
  assign n41125 = P1_P2_INSTQUEUE_REG_4__2_ & n41020;
  assign n41126 = ~n41122 & ~n41123;
  assign n41127 = ~n41124 & n41126;
  assign n41128 = ~n41125 & n41127;
  assign n41129 = P1_P2_INSTQUEUE_REG_3__2_ & n41026;
  assign n41130 = P1_P2_INSTQUEUE_REG_2__2_ & n41028;
  assign n41131 = P1_P2_INSTQUEUE_REG_1__2_ & n41030;
  assign n41132 = P1_P2_INSTQUEUE_REG_0__2_ & n41032;
  assign n41133 = ~n41129 & ~n41130;
  assign n41134 = ~n41131 & n41133;
  assign n41135 = ~n41132 & n41134;
  assign n41136 = P1_P2_INSTQUEUE_REG_15__2_ & n41038;
  assign n41137 = P1_P2_INSTQUEUE_REG_14__2_ & n41040;
  assign n41138 = P1_P2_INSTQUEUE_REG_13__2_ & n41042;
  assign n41139 = P1_P2_INSTQUEUE_REG_12__2_ & n41044;
  assign n41140 = ~n41136 & ~n41137;
  assign n41141 = ~n41138 & n41140;
  assign n41142 = ~n41139 & n41141;
  assign n41143 = P1_P2_INSTQUEUE_REG_11__2_ & n41050;
  assign n41144 = P1_P2_INSTQUEUE_REG_10__2_ & n41052;
  assign n41145 = P1_P2_INSTQUEUE_REG_9__2_ & n41054;
  assign n41146 = P1_P2_INSTQUEUE_REG_8__2_ & n41056;
  assign n41147 = ~n41143 & ~n41144;
  assign n41148 = ~n41145 & n41147;
  assign n41149 = ~n41146 & n41148;
  assign n41150 = n41128 & n41135;
  assign n41151 = n41142 & n41150;
  assign n41152 = n41149 & n41151;
  assign n41153 = n40552 & ~n41152;
  assign n41154 = ~n41121 & ~n41153;
  assign n41155 = P1_P2_EAX_REG_17_ & n41111;
  assign n41156 = ~P1_P2_EAX_REG_18_ & n41155;
  assign n41157 = P1_P2_EAX_REG_18_ & ~n41155;
  assign n41158 = ~n41156 & ~n41157;
  assign n41159 = n40558 & ~n41158;
  assign n41160 = ~n41119 & ~n41120;
  assign n41161 = n41154 & n41160;
  assign n7276 = n41159 | ~n41161;
  assign n41163 = ~n35146 & n41003;
  assign n41164 = ~n35160 & n41005;
  assign n41165 = P1_P2_EAX_REG_19_ & ~n40551;
  assign n41166 = P1_P2_INSTQUEUE_REG_7__3_ & n41014;
  assign n41167 = P1_P2_INSTQUEUE_REG_6__3_ & n41016;
  assign n41168 = P1_P2_INSTQUEUE_REG_5__3_ & n41018;
  assign n41169 = P1_P2_INSTQUEUE_REG_4__3_ & n41020;
  assign n41170 = ~n41166 & ~n41167;
  assign n41171 = ~n41168 & n41170;
  assign n41172 = ~n41169 & n41171;
  assign n41173 = P1_P2_INSTQUEUE_REG_3__3_ & n41026;
  assign n41174 = P1_P2_INSTQUEUE_REG_2__3_ & n41028;
  assign n41175 = P1_P2_INSTQUEUE_REG_1__3_ & n41030;
  assign n41176 = P1_P2_INSTQUEUE_REG_0__3_ & n41032;
  assign n41177 = ~n41173 & ~n41174;
  assign n41178 = ~n41175 & n41177;
  assign n41179 = ~n41176 & n41178;
  assign n41180 = P1_P2_INSTQUEUE_REG_15__3_ & n41038;
  assign n41181 = P1_P2_INSTQUEUE_REG_14__3_ & n41040;
  assign n41182 = P1_P2_INSTQUEUE_REG_13__3_ & n41042;
  assign n41183 = P1_P2_INSTQUEUE_REG_12__3_ & n41044;
  assign n41184 = ~n41180 & ~n41181;
  assign n41185 = ~n41182 & n41184;
  assign n41186 = ~n41183 & n41185;
  assign n41187 = P1_P2_INSTQUEUE_REG_11__3_ & n41050;
  assign n41188 = P1_P2_INSTQUEUE_REG_10__3_ & n41052;
  assign n41189 = P1_P2_INSTQUEUE_REG_9__3_ & n41054;
  assign n41190 = P1_P2_INSTQUEUE_REG_8__3_ & n41056;
  assign n41191 = ~n41187 & ~n41188;
  assign n41192 = ~n41189 & n41191;
  assign n41193 = ~n41190 & n41192;
  assign n41194 = n41172 & n41179;
  assign n41195 = n41186 & n41194;
  assign n41196 = n41193 & n41195;
  assign n41197 = n40552 & ~n41196;
  assign n41198 = ~n41165 & ~n41197;
  assign n41199 = P1_P2_EAX_REG_17_ & P1_P2_EAX_REG_18_;
  assign n41200 = n41111 & n41199;
  assign n41201 = P1_P2_EAX_REG_19_ & ~n41200;
  assign n41202 = ~P1_P2_EAX_REG_19_ & n41200;
  assign n41203 = ~n41201 & ~n41202;
  assign n41204 = n40558 & ~n41203;
  assign n41205 = ~n41163 & ~n41164;
  assign n41206 = n41198 & n41205;
  assign n7281 = n41204 | ~n41206;
  assign n41208 = ~n35124 & n41003;
  assign n41209 = ~n35138 & n41005;
  assign n41210 = P1_P2_EAX_REG_20_ & ~n40551;
  assign n41211 = P1_P2_INSTQUEUE_REG_7__4_ & n41014;
  assign n41212 = P1_P2_INSTQUEUE_REG_6__4_ & n41016;
  assign n41213 = P1_P2_INSTQUEUE_REG_5__4_ & n41018;
  assign n41214 = P1_P2_INSTQUEUE_REG_4__4_ & n41020;
  assign n41215 = ~n41211 & ~n41212;
  assign n41216 = ~n41213 & n41215;
  assign n41217 = ~n41214 & n41216;
  assign n41218 = P1_P2_INSTQUEUE_REG_3__4_ & n41026;
  assign n41219 = P1_P2_INSTQUEUE_REG_2__4_ & n41028;
  assign n41220 = P1_P2_INSTQUEUE_REG_1__4_ & n41030;
  assign n41221 = P1_P2_INSTQUEUE_REG_0__4_ & n41032;
  assign n41222 = ~n41218 & ~n41219;
  assign n41223 = ~n41220 & n41222;
  assign n41224 = ~n41221 & n41223;
  assign n41225 = P1_P2_INSTQUEUE_REG_15__4_ & n41038;
  assign n41226 = P1_P2_INSTQUEUE_REG_14__4_ & n41040;
  assign n41227 = P1_P2_INSTQUEUE_REG_13__4_ & n41042;
  assign n41228 = P1_P2_INSTQUEUE_REG_12__4_ & n41044;
  assign n41229 = ~n41225 & ~n41226;
  assign n41230 = ~n41227 & n41229;
  assign n41231 = ~n41228 & n41230;
  assign n41232 = P1_P2_INSTQUEUE_REG_11__4_ & n41050;
  assign n41233 = P1_P2_INSTQUEUE_REG_10__4_ & n41052;
  assign n41234 = P1_P2_INSTQUEUE_REG_9__4_ & n41054;
  assign n41235 = P1_P2_INSTQUEUE_REG_8__4_ & n41056;
  assign n41236 = ~n41232 & ~n41233;
  assign n41237 = ~n41234 & n41236;
  assign n41238 = ~n41235 & n41237;
  assign n41239 = n41217 & n41224;
  assign n41240 = n41231 & n41239;
  assign n41241 = n41238 & n41240;
  assign n41242 = n40552 & ~n41241;
  assign n41243 = ~n41210 & ~n41242;
  assign n41244 = P1_P2_EAX_REG_19_ & n41200;
  assign n41245 = ~P1_P2_EAX_REG_20_ & n41244;
  assign n41246 = P1_P2_EAX_REG_20_ & ~n41244;
  assign n41247 = ~n41245 & ~n41246;
  assign n41248 = n40558 & ~n41247;
  assign n41249 = ~n41208 & ~n41209;
  assign n41250 = n41243 & n41249;
  assign n7286 = n41248 | ~n41250;
  assign n41252 = ~n35102 & n41003;
  assign n41253 = ~n35116 & n41005;
  assign n41254 = P1_P2_EAX_REG_21_ & ~n40551;
  assign n41255 = P1_P2_INSTQUEUE_REG_7__5_ & n41014;
  assign n41256 = P1_P2_INSTQUEUE_REG_6__5_ & n41016;
  assign n41257 = P1_P2_INSTQUEUE_REG_5__5_ & n41018;
  assign n41258 = P1_P2_INSTQUEUE_REG_4__5_ & n41020;
  assign n41259 = ~n41255 & ~n41256;
  assign n41260 = ~n41257 & n41259;
  assign n41261 = ~n41258 & n41260;
  assign n41262 = P1_P2_INSTQUEUE_REG_3__5_ & n41026;
  assign n41263 = P1_P2_INSTQUEUE_REG_2__5_ & n41028;
  assign n41264 = P1_P2_INSTQUEUE_REG_1__5_ & n41030;
  assign n41265 = P1_P2_INSTQUEUE_REG_0__5_ & n41032;
  assign n41266 = ~n41262 & ~n41263;
  assign n41267 = ~n41264 & n41266;
  assign n41268 = ~n41265 & n41267;
  assign n41269 = P1_P2_INSTQUEUE_REG_15__5_ & n41038;
  assign n41270 = P1_P2_INSTQUEUE_REG_14__5_ & n41040;
  assign n41271 = P1_P2_INSTQUEUE_REG_13__5_ & n41042;
  assign n41272 = P1_P2_INSTQUEUE_REG_12__5_ & n41044;
  assign n41273 = ~n41269 & ~n41270;
  assign n41274 = ~n41271 & n41273;
  assign n41275 = ~n41272 & n41274;
  assign n41276 = P1_P2_INSTQUEUE_REG_11__5_ & n41050;
  assign n41277 = P1_P2_INSTQUEUE_REG_10__5_ & n41052;
  assign n41278 = P1_P2_INSTQUEUE_REG_9__5_ & n41054;
  assign n41279 = P1_P2_INSTQUEUE_REG_8__5_ & n41056;
  assign n41280 = ~n41276 & ~n41277;
  assign n41281 = ~n41278 & n41280;
  assign n41282 = ~n41279 & n41281;
  assign n41283 = n41261 & n41268;
  assign n41284 = n41275 & n41283;
  assign n41285 = n41282 & n41284;
  assign n41286 = n40552 & ~n41285;
  assign n41287 = ~n41254 & ~n41286;
  assign n41288 = P1_P2_EAX_REG_19_ & P1_P2_EAX_REG_20_;
  assign n41289 = n41200 & n41288;
  assign n41290 = P1_P2_EAX_REG_21_ & ~n41289;
  assign n41291 = ~P1_P2_EAX_REG_21_ & n41289;
  assign n41292 = ~n41290 & ~n41291;
  assign n41293 = n40558 & ~n41292;
  assign n41294 = ~n41252 & ~n41253;
  assign n41295 = n41287 & n41294;
  assign n7291 = n41293 | ~n41295;
  assign n41297 = ~n35080 & n41003;
  assign n41298 = ~n35094 & n41005;
  assign n41299 = P1_P2_EAX_REG_22_ & ~n40551;
  assign n41300 = P1_P2_INSTQUEUE_REG_7__6_ & n41014;
  assign n41301 = P1_P2_INSTQUEUE_REG_6__6_ & n41016;
  assign n41302 = P1_P2_INSTQUEUE_REG_5__6_ & n41018;
  assign n41303 = P1_P2_INSTQUEUE_REG_4__6_ & n41020;
  assign n41304 = ~n41300 & ~n41301;
  assign n41305 = ~n41302 & n41304;
  assign n41306 = ~n41303 & n41305;
  assign n41307 = P1_P2_INSTQUEUE_REG_3__6_ & n41026;
  assign n41308 = P1_P2_INSTQUEUE_REG_2__6_ & n41028;
  assign n41309 = P1_P2_INSTQUEUE_REG_1__6_ & n41030;
  assign n41310 = P1_P2_INSTQUEUE_REG_0__6_ & n41032;
  assign n41311 = ~n41307 & ~n41308;
  assign n41312 = ~n41309 & n41311;
  assign n41313 = ~n41310 & n41312;
  assign n41314 = P1_P2_INSTQUEUE_REG_15__6_ & n41038;
  assign n41315 = P1_P2_INSTQUEUE_REG_14__6_ & n41040;
  assign n41316 = P1_P2_INSTQUEUE_REG_13__6_ & n41042;
  assign n41317 = P1_P2_INSTQUEUE_REG_12__6_ & n41044;
  assign n41318 = ~n41314 & ~n41315;
  assign n41319 = ~n41316 & n41318;
  assign n41320 = ~n41317 & n41319;
  assign n41321 = P1_P2_INSTQUEUE_REG_11__6_ & n41050;
  assign n41322 = P1_P2_INSTQUEUE_REG_10__6_ & n41052;
  assign n41323 = P1_P2_INSTQUEUE_REG_9__6_ & n41054;
  assign n41324 = P1_P2_INSTQUEUE_REG_8__6_ & n41056;
  assign n41325 = ~n41321 & ~n41322;
  assign n41326 = ~n41323 & n41325;
  assign n41327 = ~n41324 & n41326;
  assign n41328 = n41306 & n41313;
  assign n41329 = n41320 & n41328;
  assign n41330 = n41327 & n41329;
  assign n41331 = n40552 & ~n41330;
  assign n41332 = ~n41299 & ~n41331;
  assign n41333 = P1_P2_EAX_REG_21_ & n41289;
  assign n41334 = ~P1_P2_EAX_REG_22_ & n41333;
  assign n41335 = P1_P2_EAX_REG_22_ & ~n41333;
  assign n41336 = ~n41334 & ~n41335;
  assign n41337 = n40558 & ~n41336;
  assign n41338 = ~n41297 & ~n41298;
  assign n41339 = n41332 & n41338;
  assign n7296 = n41337 | ~n41339;
  assign n41341 = ~n35052 & n41003;
  assign n41342 = ~n35072 & n41005;
  assign n41343 = P1_P2_EAX_REG_23_ & ~n40551;
  assign n41344 = P1_P2_INSTQUEUERD_ADDR_REG_3_ & ~P1_P2_INSTQUEUERD_ADDR_REG_2_;
  assign n41345 = ~n34331 & ~n41344;
  assign n41346 = n34302 & n41345;
  assign n41347 = P1_P2_INSTQUEUE_REG_7__0_ & n41346;
  assign n41348 = n34306 & n41345;
  assign n41349 = P1_P2_INSTQUEUE_REG_6__0_ & n41348;
  assign n41350 = n34311 & n41345;
  assign n41351 = P1_P2_INSTQUEUE_REG_5__0_ & n41350;
  assign n41352 = n34315 & n41345;
  assign n41353 = P1_P2_INSTQUEUE_REG_4__0_ & n41352;
  assign n41354 = ~n41347 & ~n41349;
  assign n41355 = ~n41351 & n41354;
  assign n41356 = ~n41353 & n41355;
  assign n41357 = P1_P2_INSTQUEUERD_ADDR_REG_2_ & n41345;
  assign n41358 = n34301 & n41357;
  assign n41359 = P1_P2_INSTQUEUE_REG_3__0_ & n41358;
  assign n41360 = n34305 & n41357;
  assign n41361 = P1_P2_INSTQUEUE_REG_2__0_ & n41360;
  assign n41362 = n34310 & n41357;
  assign n41363 = P1_P2_INSTQUEUE_REG_1__0_ & n41362;
  assign n41364 = n34314 & n41357;
  assign n41365 = P1_P2_INSTQUEUE_REG_0__0_ & n41364;
  assign n41366 = ~n41359 & ~n41361;
  assign n41367 = ~n41363 & n41366;
  assign n41368 = ~n41365 & n41367;
  assign n41369 = n34302 & ~n41345;
  assign n41370 = P1_P2_INSTQUEUE_REG_15__0_ & n41369;
  assign n41371 = n34306 & ~n41345;
  assign n41372 = P1_P2_INSTQUEUE_REG_14__0_ & n41371;
  assign n41373 = n34311 & ~n41345;
  assign n41374 = P1_P2_INSTQUEUE_REG_13__0_ & n41373;
  assign n41375 = n34315 & ~n41345;
  assign n41376 = P1_P2_INSTQUEUE_REG_12__0_ & n41375;
  assign n41377 = ~n41370 & ~n41372;
  assign n41378 = ~n41374 & n41377;
  assign n41379 = ~n41376 & n41378;
  assign n41380 = P1_P2_INSTQUEUERD_ADDR_REG_2_ & ~n41345;
  assign n41381 = n34301 & n41380;
  assign n41382 = P1_P2_INSTQUEUE_REG_11__0_ & n41381;
  assign n41383 = n34305 & n41380;
  assign n41384 = P1_P2_INSTQUEUE_REG_10__0_ & n41383;
  assign n41385 = n34310 & n41380;
  assign n41386 = P1_P2_INSTQUEUE_REG_9__0_ & n41385;
  assign n41387 = n34314 & n41380;
  assign n41388 = P1_P2_INSTQUEUE_REG_8__0_ & n41387;
  assign n41389 = ~n41382 & ~n41384;
  assign n41390 = ~n41386 & n41389;
  assign n41391 = ~n41388 & n41390;
  assign n41392 = n41356 & n41368;
  assign n41393 = n41379 & n41392;
  assign n41394 = n41391 & n41393;
  assign n41395 = P1_P2_INSTQUEUE_REG_7__7_ & n41014;
  assign n41396 = P1_P2_INSTQUEUE_REG_6__7_ & n41016;
  assign n41397 = P1_P2_INSTQUEUE_REG_5__7_ & n41018;
  assign n41398 = P1_P2_INSTQUEUE_REG_4__7_ & n41020;
  assign n41399 = ~n41395 & ~n41396;
  assign n41400 = ~n41397 & n41399;
  assign n41401 = ~n41398 & n41400;
  assign n41402 = P1_P2_INSTQUEUE_REG_3__7_ & n41026;
  assign n41403 = P1_P2_INSTQUEUE_REG_2__7_ & n41028;
  assign n41404 = P1_P2_INSTQUEUE_REG_1__7_ & n41030;
  assign n41405 = P1_P2_INSTQUEUE_REG_0__7_ & n41032;
  assign n41406 = ~n41402 & ~n41403;
  assign n41407 = ~n41404 & n41406;
  assign n41408 = ~n41405 & n41407;
  assign n41409 = P1_P2_INSTQUEUE_REG_15__7_ & n41038;
  assign n41410 = P1_P2_INSTQUEUE_REG_14__7_ & n41040;
  assign n41411 = P1_P2_INSTQUEUE_REG_13__7_ & n41042;
  assign n41412 = P1_P2_INSTQUEUE_REG_12__7_ & n41044;
  assign n41413 = ~n41409 & ~n41410;
  assign n41414 = ~n41411 & n41413;
  assign n41415 = ~n41412 & n41414;
  assign n41416 = P1_P2_INSTQUEUE_REG_11__7_ & n41050;
  assign n41417 = P1_P2_INSTQUEUE_REG_10__7_ & n41052;
  assign n41418 = P1_P2_INSTQUEUE_REG_9__7_ & n41054;
  assign n41419 = P1_P2_INSTQUEUE_REG_8__7_ & n41056;
  assign n41420 = ~n41416 & ~n41417;
  assign n41421 = ~n41418 & n41420;
  assign n41422 = ~n41419 & n41421;
  assign n41423 = n41401 & n41408;
  assign n41424 = n41415 & n41423;
  assign n41425 = n41422 & n41424;
  assign n41426 = ~n41394 & n41425;
  assign n41427 = n41394 & ~n41425;
  assign n41428 = ~n41426 & ~n41427;
  assign n41429 = n40552 & ~n41428;
  assign n41430 = ~n41343 & ~n41429;
  assign n41431 = P1_P2_EAX_REG_21_ & P1_P2_EAX_REG_22_;
  assign n41432 = n41289 & n41431;
  assign n41433 = P1_P2_EAX_REG_23_ & ~n41432;
  assign n41434 = ~P1_P2_EAX_REG_23_ & n41432;
  assign n41435 = ~n41433 & ~n41434;
  assign n41436 = n40558 & ~n41435;
  assign n41437 = ~n41341 & ~n41342;
  assign n41438 = n41430 & n41437;
  assign n7301 = n41436 | ~n41438;
  assign n41440 = ~n35220 & n41003;
  assign n41441 = ~n40281 & n41005;
  assign n41442 = P1_P2_EAX_REG_24_ & ~n40551;
  assign n41443 = ~n41394 & ~n41425;
  assign n41444 = P1_P2_INSTQUEUE_REG_7__1_ & n41346;
  assign n41445 = P1_P2_INSTQUEUE_REG_6__1_ & n41348;
  assign n41446 = P1_P2_INSTQUEUE_REG_5__1_ & n41350;
  assign n41447 = P1_P2_INSTQUEUE_REG_4__1_ & n41352;
  assign n41448 = ~n41444 & ~n41445;
  assign n41449 = ~n41446 & n41448;
  assign n41450 = ~n41447 & n41449;
  assign n41451 = P1_P2_INSTQUEUE_REG_3__1_ & n41358;
  assign n41452 = P1_P2_INSTQUEUE_REG_2__1_ & n41360;
  assign n41453 = P1_P2_INSTQUEUE_REG_1__1_ & n41362;
  assign n41454 = P1_P2_INSTQUEUE_REG_0__1_ & n41364;
  assign n41455 = ~n41451 & ~n41452;
  assign n41456 = ~n41453 & n41455;
  assign n41457 = ~n41454 & n41456;
  assign n41458 = P1_P2_INSTQUEUE_REG_15__1_ & n41369;
  assign n41459 = P1_P2_INSTQUEUE_REG_14__1_ & n41371;
  assign n41460 = P1_P2_INSTQUEUE_REG_13__1_ & n41373;
  assign n41461 = P1_P2_INSTQUEUE_REG_12__1_ & n41375;
  assign n41462 = ~n41458 & ~n41459;
  assign n41463 = ~n41460 & n41462;
  assign n41464 = ~n41461 & n41463;
  assign n41465 = P1_P2_INSTQUEUE_REG_11__1_ & n41381;
  assign n41466 = P1_P2_INSTQUEUE_REG_10__1_ & n41383;
  assign n41467 = P1_P2_INSTQUEUE_REG_9__1_ & n41385;
  assign n41468 = P1_P2_INSTQUEUE_REG_8__1_ & n41387;
  assign n41469 = ~n41465 & ~n41466;
  assign n41470 = ~n41467 & n41469;
  assign n41471 = ~n41468 & n41470;
  assign n41472 = n41450 & n41457;
  assign n41473 = n41464 & n41472;
  assign n41474 = n41471 & n41473;
  assign n41475 = n41443 & n41474;
  assign n41476 = ~n41443 & ~n41474;
  assign n41477 = ~n41475 & ~n41476;
  assign n41478 = n40552 & ~n41477;
  assign n41479 = ~n41442 & ~n41478;
  assign n41480 = P1_P2_EAX_REG_23_ & n41432;
  assign n41481 = ~P1_P2_EAX_REG_24_ & n41480;
  assign n41482 = P1_P2_EAX_REG_24_ & ~n41480;
  assign n41483 = ~n41481 & ~n41482;
  assign n41484 = n40558 & ~n41483;
  assign n41485 = ~n41440 & ~n41441;
  assign n41486 = n41479 & n41485;
  assign n7306 = n41484 | ~n41486;
  assign n41488 = ~n35198 & n41003;
  assign n41489 = ~n40273 & n41005;
  assign n41490 = P1_P2_EAX_REG_25_ & ~n40551;
  assign n41491 = n41443 & ~n41474;
  assign n41492 = P1_P2_INSTQUEUE_REG_7__2_ & n41346;
  assign n41493 = P1_P2_INSTQUEUE_REG_6__2_ & n41348;
  assign n41494 = P1_P2_INSTQUEUE_REG_5__2_ & n41350;
  assign n41495 = P1_P2_INSTQUEUE_REG_4__2_ & n41352;
  assign n41496 = ~n41492 & ~n41493;
  assign n41497 = ~n41494 & n41496;
  assign n41498 = ~n41495 & n41497;
  assign n41499 = P1_P2_INSTQUEUE_REG_3__2_ & n41358;
  assign n41500 = P1_P2_INSTQUEUE_REG_2__2_ & n41360;
  assign n41501 = P1_P2_INSTQUEUE_REG_1__2_ & n41362;
  assign n41502 = P1_P2_INSTQUEUE_REG_0__2_ & n41364;
  assign n41503 = ~n41499 & ~n41500;
  assign n41504 = ~n41501 & n41503;
  assign n41505 = ~n41502 & n41504;
  assign n41506 = P1_P2_INSTQUEUE_REG_15__2_ & n41369;
  assign n41507 = P1_P2_INSTQUEUE_REG_14__2_ & n41371;
  assign n41508 = P1_P2_INSTQUEUE_REG_13__2_ & n41373;
  assign n41509 = P1_P2_INSTQUEUE_REG_12__2_ & n41375;
  assign n41510 = ~n41506 & ~n41507;
  assign n41511 = ~n41508 & n41510;
  assign n41512 = ~n41509 & n41511;
  assign n41513 = P1_P2_INSTQUEUE_REG_11__2_ & n41381;
  assign n41514 = P1_P2_INSTQUEUE_REG_10__2_ & n41383;
  assign n41515 = P1_P2_INSTQUEUE_REG_9__2_ & n41385;
  assign n41516 = P1_P2_INSTQUEUE_REG_8__2_ & n41387;
  assign n41517 = ~n41513 & ~n41514;
  assign n41518 = ~n41515 & n41517;
  assign n41519 = ~n41516 & n41518;
  assign n41520 = n41498 & n41505;
  assign n41521 = n41512 & n41520;
  assign n41522 = n41519 & n41521;
  assign n41523 = n41491 & n41522;
  assign n41524 = ~n41491 & ~n41522;
  assign n41525 = ~n41523 & ~n41524;
  assign n41526 = n40552 & ~n41525;
  assign n41527 = ~n41490 & ~n41526;
  assign n41528 = P1_P2_EAX_REG_23_ & P1_P2_EAX_REG_24_;
  assign n41529 = n41432 & n41528;
  assign n41530 = P1_P2_EAX_REG_25_ & ~n41529;
  assign n41531 = ~P1_P2_EAX_REG_25_ & n41529;
  assign n41532 = ~n41530 & ~n41531;
  assign n41533 = n40558 & ~n41532;
  assign n41534 = ~n41488 & ~n41489;
  assign n41535 = n41527 & n41534;
  assign n7311 = n41533 | ~n41535;
  assign n41537 = ~n35176 & n41003;
  assign n41538 = ~n40265 & n41005;
  assign n41539 = P1_P2_EAX_REG_26_ & ~n40551;
  assign n41540 = n41491 & ~n41522;
  assign n41541 = P1_P2_INSTQUEUE_REG_7__3_ & n41346;
  assign n41542 = P1_P2_INSTQUEUE_REG_6__3_ & n41348;
  assign n41543 = P1_P2_INSTQUEUE_REG_5__3_ & n41350;
  assign n41544 = P1_P2_INSTQUEUE_REG_4__3_ & n41352;
  assign n41545 = ~n41541 & ~n41542;
  assign n41546 = ~n41543 & n41545;
  assign n41547 = ~n41544 & n41546;
  assign n41548 = P1_P2_INSTQUEUE_REG_3__3_ & n41358;
  assign n41549 = P1_P2_INSTQUEUE_REG_2__3_ & n41360;
  assign n41550 = P1_P2_INSTQUEUE_REG_1__3_ & n41362;
  assign n41551 = P1_P2_INSTQUEUE_REG_0__3_ & n41364;
  assign n41552 = ~n41548 & ~n41549;
  assign n41553 = ~n41550 & n41552;
  assign n41554 = ~n41551 & n41553;
  assign n41555 = P1_P2_INSTQUEUE_REG_15__3_ & n41369;
  assign n41556 = P1_P2_INSTQUEUE_REG_14__3_ & n41371;
  assign n41557 = P1_P2_INSTQUEUE_REG_13__3_ & n41373;
  assign n41558 = P1_P2_INSTQUEUE_REG_12__3_ & n41375;
  assign n41559 = ~n41555 & ~n41556;
  assign n41560 = ~n41557 & n41559;
  assign n41561 = ~n41558 & n41560;
  assign n41562 = P1_P2_INSTQUEUE_REG_11__3_ & n41381;
  assign n41563 = P1_P2_INSTQUEUE_REG_10__3_ & n41383;
  assign n41564 = P1_P2_INSTQUEUE_REG_9__3_ & n41385;
  assign n41565 = P1_P2_INSTQUEUE_REG_8__3_ & n41387;
  assign n41566 = ~n41562 & ~n41563;
  assign n41567 = ~n41564 & n41566;
  assign n41568 = ~n41565 & n41567;
  assign n41569 = n41547 & n41554;
  assign n41570 = n41561 & n41569;
  assign n41571 = n41568 & n41570;
  assign n41572 = n41540 & n41571;
  assign n41573 = ~n41540 & ~n41571;
  assign n41574 = ~n41572 & ~n41573;
  assign n41575 = n40552 & ~n41574;
  assign n41576 = ~n41539 & ~n41575;
  assign n41577 = P1_P2_EAX_REG_25_ & n41529;
  assign n41578 = ~P1_P2_EAX_REG_26_ & n41577;
  assign n41579 = P1_P2_EAX_REG_26_ & ~n41577;
  assign n41580 = ~n41578 & ~n41579;
  assign n41581 = n40558 & ~n41580;
  assign n41582 = ~n41537 & ~n41538;
  assign n41583 = n41576 & n41582;
  assign n7316 = n41581 | ~n41583;
  assign n41585 = ~n35154 & n41003;
  assign n41586 = ~n40257 & n41005;
  assign n41587 = P1_P2_EAX_REG_27_ & ~n40551;
  assign n41588 = n41540 & ~n41571;
  assign n41589 = P1_P2_INSTQUEUE_REG_7__4_ & n41346;
  assign n41590 = P1_P2_INSTQUEUE_REG_6__4_ & n41348;
  assign n41591 = P1_P2_INSTQUEUE_REG_5__4_ & n41350;
  assign n41592 = P1_P2_INSTQUEUE_REG_4__4_ & n41352;
  assign n41593 = ~n41589 & ~n41590;
  assign n41594 = ~n41591 & n41593;
  assign n41595 = ~n41592 & n41594;
  assign n41596 = P1_P2_INSTQUEUE_REG_3__4_ & n41358;
  assign n41597 = P1_P2_INSTQUEUE_REG_2__4_ & n41360;
  assign n41598 = P1_P2_INSTQUEUE_REG_1__4_ & n41362;
  assign n41599 = P1_P2_INSTQUEUE_REG_0__4_ & n41364;
  assign n41600 = ~n41596 & ~n41597;
  assign n41601 = ~n41598 & n41600;
  assign n41602 = ~n41599 & n41601;
  assign n41603 = P1_P2_INSTQUEUE_REG_15__4_ & n41369;
  assign n41604 = P1_P2_INSTQUEUE_REG_14__4_ & n41371;
  assign n41605 = P1_P2_INSTQUEUE_REG_13__4_ & n41373;
  assign n41606 = P1_P2_INSTQUEUE_REG_12__4_ & n41375;
  assign n41607 = ~n41603 & ~n41604;
  assign n41608 = ~n41605 & n41607;
  assign n41609 = ~n41606 & n41608;
  assign n41610 = P1_P2_INSTQUEUE_REG_11__4_ & n41381;
  assign n41611 = P1_P2_INSTQUEUE_REG_10__4_ & n41383;
  assign n41612 = P1_P2_INSTQUEUE_REG_9__4_ & n41385;
  assign n41613 = P1_P2_INSTQUEUE_REG_8__4_ & n41387;
  assign n41614 = ~n41610 & ~n41611;
  assign n41615 = ~n41612 & n41614;
  assign n41616 = ~n41613 & n41615;
  assign n41617 = n41595 & n41602;
  assign n41618 = n41609 & n41617;
  assign n41619 = n41616 & n41618;
  assign n41620 = n41588 & n41619;
  assign n41621 = ~n41588 & ~n41619;
  assign n41622 = ~n41620 & ~n41621;
  assign n41623 = n40552 & ~n41622;
  assign n41624 = ~n41587 & ~n41623;
  assign n41625 = P1_P2_EAX_REG_25_ & P1_P2_EAX_REG_26_;
  assign n41626 = n41529 & n41625;
  assign n41627 = P1_P2_EAX_REG_27_ & ~n41626;
  assign n41628 = ~P1_P2_EAX_REG_27_ & n41626;
  assign n41629 = ~n41627 & ~n41628;
  assign n41630 = n40558 & ~n41629;
  assign n41631 = ~n41585 & ~n41586;
  assign n41632 = n41624 & n41631;
  assign n7321 = n41630 | ~n41632;
  assign n41634 = ~n35132 & n41003;
  assign n41635 = ~n40249 & n41005;
  assign n41636 = P1_P2_EAX_REG_28_ & ~n40551;
  assign n41637 = n41588 & ~n41619;
  assign n41638 = P1_P2_INSTQUEUE_REG_7__5_ & n41346;
  assign n41639 = P1_P2_INSTQUEUE_REG_6__5_ & n41348;
  assign n41640 = P1_P2_INSTQUEUE_REG_5__5_ & n41350;
  assign n41641 = P1_P2_INSTQUEUE_REG_4__5_ & n41352;
  assign n41642 = ~n41638 & ~n41639;
  assign n41643 = ~n41640 & n41642;
  assign n41644 = ~n41641 & n41643;
  assign n41645 = P1_P2_INSTQUEUE_REG_3__5_ & n41358;
  assign n41646 = P1_P2_INSTQUEUE_REG_2__5_ & n41360;
  assign n41647 = P1_P2_INSTQUEUE_REG_1__5_ & n41362;
  assign n41648 = P1_P2_INSTQUEUE_REG_0__5_ & n41364;
  assign n41649 = ~n41645 & ~n41646;
  assign n41650 = ~n41647 & n41649;
  assign n41651 = ~n41648 & n41650;
  assign n41652 = P1_P2_INSTQUEUE_REG_15__5_ & n41369;
  assign n41653 = P1_P2_INSTQUEUE_REG_14__5_ & n41371;
  assign n41654 = P1_P2_INSTQUEUE_REG_13__5_ & n41373;
  assign n41655 = P1_P2_INSTQUEUE_REG_12__5_ & n41375;
  assign n41656 = ~n41652 & ~n41653;
  assign n41657 = ~n41654 & n41656;
  assign n41658 = ~n41655 & n41657;
  assign n41659 = P1_P2_INSTQUEUE_REG_11__5_ & n41381;
  assign n41660 = P1_P2_INSTQUEUE_REG_10__5_ & n41383;
  assign n41661 = P1_P2_INSTQUEUE_REG_9__5_ & n41385;
  assign n41662 = P1_P2_INSTQUEUE_REG_8__5_ & n41387;
  assign n41663 = ~n41659 & ~n41660;
  assign n41664 = ~n41661 & n41663;
  assign n41665 = ~n41662 & n41664;
  assign n41666 = n41644 & n41651;
  assign n41667 = n41658 & n41666;
  assign n41668 = n41665 & n41667;
  assign n41669 = n41637 & n41668;
  assign n41670 = ~n41637 & ~n41668;
  assign n41671 = ~n41669 & ~n41670;
  assign n41672 = n40552 & ~n41671;
  assign n41673 = P1_P2_EAX_REG_27_ & n41626;
  assign n41674 = ~P1_P2_EAX_REG_28_ & n41673;
  assign n41675 = P1_P2_EAX_REG_28_ & ~n41673;
  assign n41676 = ~n41674 & ~n41675;
  assign n41677 = n40558 & ~n41676;
  assign n41678 = ~n41634 & ~n41635;
  assign n41679 = ~n41636 & n41678;
  assign n41680 = ~n41672 & n41679;
  assign n7326 = n41677 | ~n41680;
  assign n41682 = ~n35110 & n41003;
  assign n41683 = ~n40241 & n41005;
  assign n41684 = P1_P2_EAX_REG_29_ & ~n40551;
  assign n41685 = n41637 & ~n41668;
  assign n41686 = P1_P2_INSTQUEUE_REG_7__6_ & n41346;
  assign n41687 = P1_P2_INSTQUEUE_REG_6__6_ & n41348;
  assign n41688 = P1_P2_INSTQUEUE_REG_5__6_ & n41350;
  assign n41689 = P1_P2_INSTQUEUE_REG_4__6_ & n41352;
  assign n41690 = ~n41686 & ~n41687;
  assign n41691 = ~n41688 & n41690;
  assign n41692 = ~n41689 & n41691;
  assign n41693 = P1_P2_INSTQUEUE_REG_3__6_ & n41358;
  assign n41694 = P1_P2_INSTQUEUE_REG_2__6_ & n41360;
  assign n41695 = P1_P2_INSTQUEUE_REG_1__6_ & n41362;
  assign n41696 = P1_P2_INSTQUEUE_REG_0__6_ & n41364;
  assign n41697 = ~n41693 & ~n41694;
  assign n41698 = ~n41695 & n41697;
  assign n41699 = ~n41696 & n41698;
  assign n41700 = P1_P2_INSTQUEUE_REG_15__6_ & n41369;
  assign n41701 = P1_P2_INSTQUEUE_REG_14__6_ & n41371;
  assign n41702 = P1_P2_INSTQUEUE_REG_13__6_ & n41373;
  assign n41703 = P1_P2_INSTQUEUE_REG_12__6_ & n41375;
  assign n41704 = ~n41700 & ~n41701;
  assign n41705 = ~n41702 & n41704;
  assign n41706 = ~n41703 & n41705;
  assign n41707 = P1_P2_INSTQUEUE_REG_11__6_ & n41381;
  assign n41708 = P1_P2_INSTQUEUE_REG_10__6_ & n41383;
  assign n41709 = P1_P2_INSTQUEUE_REG_9__6_ & n41385;
  assign n41710 = P1_P2_INSTQUEUE_REG_8__6_ & n41387;
  assign n41711 = ~n41707 & ~n41708;
  assign n41712 = ~n41709 & n41711;
  assign n41713 = ~n41710 & n41712;
  assign n41714 = n41692 & n41699;
  assign n41715 = n41706 & n41714;
  assign n41716 = n41713 & n41715;
  assign n41717 = n41685 & n41716;
  assign n41718 = ~n41685 & ~n41716;
  assign n41719 = ~n41717 & ~n41718;
  assign n41720 = n40552 & ~n41719;
  assign n41721 = P1_P2_EAX_REG_27_ & P1_P2_EAX_REG_28_;
  assign n41722 = n41626 & n41721;
  assign n41723 = P1_P2_EAX_REG_29_ & ~n41722;
  assign n41724 = ~P1_P2_EAX_REG_29_ & n41722;
  assign n41725 = ~n41723 & ~n41724;
  assign n41726 = n40558 & ~n41725;
  assign n41727 = ~n41682 & ~n41683;
  assign n41728 = ~n41684 & n41727;
  assign n41729 = ~n41720 & n41728;
  assign n7331 = n41726 | ~n41729;
  assign n41731 = ~n35088 & n41003;
  assign n41732 = ~n40233 & n41005;
  assign n41733 = P1_P2_EAX_REG_30_ & ~n40551;
  assign n41734 = n41685 & ~n41716;
  assign n41735 = P1_P2_INSTQUEUE_REG_7__7_ & n41346;
  assign n41736 = P1_P2_INSTQUEUE_REG_6__7_ & n41348;
  assign n41737 = P1_P2_INSTQUEUE_REG_5__7_ & n41350;
  assign n41738 = P1_P2_INSTQUEUE_REG_4__7_ & n41352;
  assign n41739 = ~n41735 & ~n41736;
  assign n41740 = ~n41737 & n41739;
  assign n41741 = ~n41738 & n41740;
  assign n41742 = P1_P2_INSTQUEUE_REG_3__7_ & n41358;
  assign n41743 = P1_P2_INSTQUEUE_REG_2__7_ & n41360;
  assign n41744 = P1_P2_INSTQUEUE_REG_1__7_ & n41362;
  assign n41745 = P1_P2_INSTQUEUE_REG_0__7_ & n41364;
  assign n41746 = ~n41742 & ~n41743;
  assign n41747 = ~n41744 & n41746;
  assign n41748 = ~n41745 & n41747;
  assign n41749 = P1_P2_INSTQUEUE_REG_15__7_ & n41369;
  assign n41750 = P1_P2_INSTQUEUE_REG_14__7_ & n41371;
  assign n41751 = P1_P2_INSTQUEUE_REG_13__7_ & n41373;
  assign n41752 = P1_P2_INSTQUEUE_REG_12__7_ & n41375;
  assign n41753 = ~n41749 & ~n41750;
  assign n41754 = ~n41751 & n41753;
  assign n41755 = ~n41752 & n41754;
  assign n41756 = P1_P2_INSTQUEUE_REG_11__7_ & n41381;
  assign n41757 = P1_P2_INSTQUEUE_REG_10__7_ & n41383;
  assign n41758 = P1_P2_INSTQUEUE_REG_9__7_ & n41385;
  assign n41759 = P1_P2_INSTQUEUE_REG_8__7_ & n41387;
  assign n41760 = ~n41756 & ~n41757;
  assign n41761 = ~n41758 & n41760;
  assign n41762 = ~n41759 & n41761;
  assign n41763 = n41741 & n41748;
  assign n41764 = n41755 & n41763;
  assign n41765 = n41762 & n41764;
  assign n41766 = n41734 & n41765;
  assign n41767 = ~n41734 & ~n41765;
  assign n41768 = ~n41766 & ~n41767;
  assign n41769 = n40552 & ~n41768;
  assign n41770 = P1_P2_EAX_REG_29_ & n41722;
  assign n41771 = ~P1_P2_EAX_REG_30_ & n41770;
  assign n41772 = P1_P2_EAX_REG_30_ & ~n41770;
  assign n41773 = ~n41771 & ~n41772;
  assign n41774 = n40558 & ~n41773;
  assign n41775 = ~n41731 & ~n41732;
  assign n41776 = ~n41733 & n41775;
  assign n41777 = ~n41769 & n41776;
  assign n7336 = n41774 | ~n41777;
  assign n41779 = P1_P2_EAX_REG_31_ & ~n40551;
  assign n41780 = ~n35063 & n41003;
  assign n41781 = P1_P2_EAX_REG_30_ & n41770;
  assign n41782 = ~P1_P2_EAX_REG_31_ & n41781;
  assign n41783 = P1_P2_EAX_REG_31_ & ~n41781;
  assign n41784 = ~n41782 & ~n41783;
  assign n41785 = n40558 & ~n41784;
  assign n41786 = ~n41779 & ~n41780;
  assign n7341 = n41785 | ~n41786;
  assign n41788 = ~n34722 & ~n34816;
  assign n41789 = n34935 & ~n41788;
  assign n41790 = n34452 & n41789;
  assign n41791 = ~P1_P2_EBX_REG_0_ & n41790;
  assign n41792 = ~n34452 & n41789;
  assign n41793 = P1_P2_INSTQUEUE_REG_0__0_ & n41792;
  assign n41794 = P1_P2_EBX_REG_0_ & ~n41789;
  assign n41795 = ~n41791 & ~n41793;
  assign n7346 = n41794 | ~n41795;
  assign n41797 = ~P1_P2_EBX_REG_0_ & P1_P2_EBX_REG_1_;
  assign n41798 = P1_P2_EBX_REG_0_ & ~P1_P2_EBX_REG_1_;
  assign n41799 = ~n41797 & ~n41798;
  assign n41800 = n41790 & ~n41799;
  assign n41801 = P1_P2_INSTQUEUE_REG_0__1_ & n41792;
  assign n41802 = P1_P2_EBX_REG_1_ & ~n41789;
  assign n41803 = ~n41800 & ~n41801;
  assign n7351 = n41802 | ~n41803;
  assign n41805 = P1_P2_EBX_REG_0_ & P1_P2_EBX_REG_1_;
  assign n41806 = ~P1_P2_EBX_REG_2_ & n41805;
  assign n41807 = P1_P2_EBX_REG_2_ & ~n41805;
  assign n41808 = ~n41806 & ~n41807;
  assign n41809 = n41790 & ~n41808;
  assign n41810 = P1_P2_INSTQUEUE_REG_0__2_ & n41792;
  assign n41811 = P1_P2_EBX_REG_2_ & ~n41789;
  assign n41812 = ~n41809 & ~n41810;
  assign n7356 = n41811 | ~n41812;
  assign n41814 = P1_P2_EBX_REG_0_ & P1_P2_EBX_REG_2_;
  assign n41815 = P1_P2_EBX_REG_1_ & n41814;
  assign n41816 = P1_P2_EBX_REG_3_ & ~n41815;
  assign n41817 = ~P1_P2_EBX_REG_3_ & n41815;
  assign n41818 = ~n41816 & ~n41817;
  assign n41819 = n41790 & ~n41818;
  assign n41820 = P1_P2_INSTQUEUE_REG_0__3_ & n41792;
  assign n41821 = P1_P2_EBX_REG_3_ & ~n41789;
  assign n41822 = ~n41819 & ~n41820;
  assign n7361 = n41821 | ~n41822;
  assign n41824 = P1_P2_EBX_REG_3_ & n41815;
  assign n41825 = ~P1_P2_EBX_REG_4_ & n41824;
  assign n41826 = P1_P2_EBX_REG_4_ & ~n41824;
  assign n41827 = ~n41825 & ~n41826;
  assign n41828 = n41790 & ~n41827;
  assign n41829 = P1_P2_INSTQUEUE_REG_0__4_ & n41792;
  assign n41830 = P1_P2_EBX_REG_4_ & ~n41789;
  assign n41831 = ~n41828 & ~n41829;
  assign n7366 = n41830 | ~n41831;
  assign n41833 = P1_P2_EBX_REG_3_ & P1_P2_EBX_REG_4_;
  assign n41834 = n41815 & n41833;
  assign n41835 = P1_P2_EBX_REG_5_ & ~n41834;
  assign n41836 = ~P1_P2_EBX_REG_5_ & n41834;
  assign n41837 = ~n41835 & ~n41836;
  assign n41838 = n41790 & ~n41837;
  assign n41839 = P1_P2_INSTQUEUE_REG_0__5_ & n41792;
  assign n41840 = P1_P2_EBX_REG_5_ & ~n41789;
  assign n41841 = ~n41838 & ~n41839;
  assign n7371 = n41840 | ~n41841;
  assign n41843 = P1_P2_EBX_REG_5_ & n41834;
  assign n41844 = ~P1_P2_EBX_REG_6_ & n41843;
  assign n41845 = P1_P2_EBX_REG_6_ & ~n41843;
  assign n41846 = ~n41844 & ~n41845;
  assign n41847 = n41790 & ~n41846;
  assign n41848 = P1_P2_INSTQUEUE_REG_0__6_ & n41792;
  assign n41849 = P1_P2_EBX_REG_6_ & ~n41789;
  assign n41850 = ~n41847 & ~n41848;
  assign n7376 = n41849 | ~n41850;
  assign n41852 = P1_P2_EBX_REG_5_ & P1_P2_EBX_REG_6_;
  assign n41853 = n41834 & n41852;
  assign n41854 = P1_P2_EBX_REG_7_ & ~n41853;
  assign n41855 = ~P1_P2_EBX_REG_7_ & n41853;
  assign n41856 = ~n41854 & ~n41855;
  assign n41857 = n41790 & ~n41856;
  assign n41858 = P1_P2_INSTQUEUE_REG_0__7_ & n41792;
  assign n41859 = P1_P2_EBX_REG_7_ & ~n41789;
  assign n41860 = ~n41857 & ~n41858;
  assign n7381 = n41859 | ~n41860;
  assign n41862 = P1_P2_EBX_REG_7_ & n41853;
  assign n41863 = ~P1_P2_EBX_REG_8_ & n41862;
  assign n41864 = P1_P2_EBX_REG_8_ & ~n41862;
  assign n41865 = ~n41863 & ~n41864;
  assign n41866 = n41790 & ~n41865;
  assign n41867 = ~n40693 & n41792;
  assign n41868 = P1_P2_EBX_REG_8_ & ~n41789;
  assign n41869 = ~n41866 & ~n41867;
  assign n7386 = n41868 | ~n41869;
  assign n41871 = P1_P2_EBX_REG_7_ & P1_P2_EBX_REG_8_;
  assign n41872 = n41853 & n41871;
  assign n41873 = P1_P2_EBX_REG_9_ & ~n41872;
  assign n41874 = ~P1_P2_EBX_REG_9_ & n41872;
  assign n41875 = ~n41873 & ~n41874;
  assign n41876 = n41790 & ~n41875;
  assign n41877 = ~n40735 & n41792;
  assign n41878 = P1_P2_EBX_REG_9_ & ~n41789;
  assign n41879 = ~n41876 & ~n41877;
  assign n7391 = n41878 | ~n41879;
  assign n41881 = P1_P2_EBX_REG_10_ & ~n41789;
  assign n41882 = ~n40778 & n41792;
  assign n41883 = P1_P2_EBX_REG_9_ & n41872;
  assign n41884 = ~P1_P2_EBX_REG_10_ & n41883;
  assign n41885 = P1_P2_EBX_REG_10_ & ~n41883;
  assign n41886 = ~n41884 & ~n41885;
  assign n41887 = n41790 & ~n41886;
  assign n41888 = ~n41881 & ~n41882;
  assign n7396 = n41887 | ~n41888;
  assign n41890 = P1_P2_EBX_REG_11_ & ~n41789;
  assign n41891 = ~n40820 & n41792;
  assign n41892 = P1_P2_EBX_REG_9_ & P1_P2_EBX_REG_10_;
  assign n41893 = n41872 & n41892;
  assign n41894 = P1_P2_EBX_REG_11_ & ~n41893;
  assign n41895 = ~P1_P2_EBX_REG_11_ & n41893;
  assign n41896 = ~n41894 & ~n41895;
  assign n41897 = n41790 & ~n41896;
  assign n41898 = ~n41890 & ~n41891;
  assign n7401 = n41897 | ~n41898;
  assign n41900 = P1_P2_EBX_REG_12_ & ~n41789;
  assign n41901 = ~n40863 & n41792;
  assign n41902 = P1_P2_EBX_REG_11_ & n41893;
  assign n41903 = ~P1_P2_EBX_REG_12_ & n41902;
  assign n41904 = P1_P2_EBX_REG_12_ & ~n41902;
  assign n41905 = ~n41903 & ~n41904;
  assign n41906 = n41790 & ~n41905;
  assign n41907 = ~n41900 & ~n41901;
  assign n7406 = n41906 | ~n41907;
  assign n41909 = P1_P2_EBX_REG_13_ & ~n41789;
  assign n41910 = ~n40906 & n41792;
  assign n41911 = P1_P2_EBX_REG_11_ & P1_P2_EBX_REG_12_;
  assign n41912 = n41893 & n41911;
  assign n41913 = P1_P2_EBX_REG_13_ & ~n41912;
  assign n41914 = ~P1_P2_EBX_REG_13_ & n41912;
  assign n41915 = ~n41913 & ~n41914;
  assign n41916 = n41790 & ~n41915;
  assign n41917 = ~n41909 & ~n41910;
  assign n7411 = n41916 | ~n41917;
  assign n41919 = P1_P2_EBX_REG_14_ & ~n41789;
  assign n41920 = ~n40949 & n41792;
  assign n41921 = P1_P2_EBX_REG_13_ & n41912;
  assign n41922 = ~P1_P2_EBX_REG_14_ & n41921;
  assign n41923 = P1_P2_EBX_REG_14_ & ~n41921;
  assign n41924 = ~n41922 & ~n41923;
  assign n41925 = n41790 & ~n41924;
  assign n41926 = ~n41919 & ~n41920;
  assign n7416 = n41925 | ~n41926;
  assign n41928 = P1_P2_EBX_REG_15_ & ~n41789;
  assign n41929 = ~n40991 & n41792;
  assign n41930 = P1_P2_EBX_REG_13_ & P1_P2_EBX_REG_14_;
  assign n41931 = n41912 & n41930;
  assign n41932 = P1_P2_EBX_REG_15_ & ~n41931;
  assign n41933 = ~P1_P2_EBX_REG_15_ & n41931;
  assign n41934 = ~n41932 & ~n41933;
  assign n41935 = n41790 & ~n41934;
  assign n41936 = ~n41928 & ~n41929;
  assign n7421 = n41935 | ~n41936;
  assign n41938 = P1_P2_EBX_REG_16_ & ~n41789;
  assign n41939 = ~n41063 & n41792;
  assign n41940 = P1_P2_EBX_REG_15_ & n41931;
  assign n41941 = ~P1_P2_EBX_REG_16_ & n41940;
  assign n41942 = P1_P2_EBX_REG_16_ & ~n41940;
  assign n41943 = ~n41941 & ~n41942;
  assign n41944 = n41790 & ~n41943;
  assign n41945 = ~n41938 & ~n41939;
  assign n7426 = n41944 | ~n41945;
  assign n41947 = P1_P2_EBX_REG_17_ & ~n41789;
  assign n41948 = ~n41107 & n41792;
  assign n41949 = P1_P2_EBX_REG_15_ & P1_P2_EBX_REG_16_;
  assign n41950 = n41931 & n41949;
  assign n41951 = P1_P2_EBX_REG_17_ & ~n41950;
  assign n41952 = ~P1_P2_EBX_REG_17_ & n41950;
  assign n41953 = ~n41951 & ~n41952;
  assign n41954 = n41790 & ~n41953;
  assign n41955 = ~n41947 & ~n41948;
  assign n7431 = n41954 | ~n41955;
  assign n41957 = P1_P2_EBX_REG_18_ & ~n41789;
  assign n41958 = ~n41152 & n41792;
  assign n41959 = P1_P2_EBX_REG_17_ & n41950;
  assign n41960 = ~P1_P2_EBX_REG_18_ & n41959;
  assign n41961 = P1_P2_EBX_REG_18_ & ~n41959;
  assign n41962 = ~n41960 & ~n41961;
  assign n41963 = n41790 & ~n41962;
  assign n41964 = ~n41957 & ~n41958;
  assign n7436 = n41963 | ~n41964;
  assign n41966 = P1_P2_EBX_REG_19_ & ~n41789;
  assign n41967 = ~n41196 & n41792;
  assign n41968 = P1_P2_EBX_REG_17_ & P1_P2_EBX_REG_18_;
  assign n41969 = n41950 & n41968;
  assign n41970 = P1_P2_EBX_REG_19_ & ~n41969;
  assign n41971 = ~P1_P2_EBX_REG_19_ & n41969;
  assign n41972 = ~n41970 & ~n41971;
  assign n41973 = n41790 & ~n41972;
  assign n41974 = ~n41966 & ~n41967;
  assign n7441 = n41973 | ~n41974;
  assign n41976 = P1_P2_EBX_REG_20_ & ~n41789;
  assign n41977 = ~n41241 & n41792;
  assign n41978 = P1_P2_EBX_REG_19_ & n41969;
  assign n41979 = ~P1_P2_EBX_REG_20_ & n41978;
  assign n41980 = P1_P2_EBX_REG_20_ & ~n41978;
  assign n41981 = ~n41979 & ~n41980;
  assign n41982 = n41790 & ~n41981;
  assign n41983 = ~n41976 & ~n41977;
  assign n7446 = n41982 | ~n41983;
  assign n41985 = P1_P2_EBX_REG_21_ & ~n41789;
  assign n41986 = ~n41285 & n41792;
  assign n41987 = P1_P2_EBX_REG_19_ & P1_P2_EBX_REG_20_;
  assign n41988 = n41969 & n41987;
  assign n41989 = P1_P2_EBX_REG_21_ & ~n41988;
  assign n41990 = ~P1_P2_EBX_REG_21_ & n41988;
  assign n41991 = ~n41989 & ~n41990;
  assign n41992 = n41790 & ~n41991;
  assign n41993 = ~n41985 & ~n41986;
  assign n7451 = n41992 | ~n41993;
  assign n41995 = P1_P2_EBX_REG_22_ & ~n41789;
  assign n41996 = ~n41330 & n41792;
  assign n41997 = P1_P2_EBX_REG_21_ & n41988;
  assign n41998 = ~P1_P2_EBX_REG_22_ & n41997;
  assign n41999 = P1_P2_EBX_REG_22_ & ~n41997;
  assign n42000 = ~n41998 & ~n41999;
  assign n42001 = n41790 & ~n42000;
  assign n42002 = ~n41995 & ~n41996;
  assign n7456 = n42001 | ~n42002;
  assign n42004 = P1_P2_EBX_REG_23_ & ~n41789;
  assign n42005 = ~n41428 & n41792;
  assign n42006 = P1_P2_EBX_REG_21_ & P1_P2_EBX_REG_22_;
  assign n42007 = n41988 & n42006;
  assign n42008 = P1_P2_EBX_REG_23_ & ~n42007;
  assign n42009 = ~P1_P2_EBX_REG_23_ & n42007;
  assign n42010 = ~n42008 & ~n42009;
  assign n42011 = n41790 & ~n42010;
  assign n42012 = ~n42004 & ~n42005;
  assign n7461 = n42011 | ~n42012;
  assign n42014 = P1_P2_EBX_REG_24_ & ~n41789;
  assign n42015 = ~n41477 & n41792;
  assign n42016 = P1_P2_EBX_REG_23_ & n42007;
  assign n42017 = ~P1_P2_EBX_REG_24_ & n42016;
  assign n42018 = P1_P2_EBX_REG_24_ & ~n42016;
  assign n42019 = ~n42017 & ~n42018;
  assign n42020 = n41790 & ~n42019;
  assign n42021 = ~n42014 & ~n42015;
  assign n7466 = n42020 | ~n42021;
  assign n42023 = P1_P2_EBX_REG_25_ & ~n41789;
  assign n42024 = ~n41525 & n41792;
  assign n42025 = P1_P2_EBX_REG_23_ & P1_P2_EBX_REG_24_;
  assign n42026 = n42007 & n42025;
  assign n42027 = P1_P2_EBX_REG_25_ & ~n42026;
  assign n42028 = ~P1_P2_EBX_REG_25_ & n42026;
  assign n42029 = ~n42027 & ~n42028;
  assign n42030 = n41790 & ~n42029;
  assign n42031 = ~n42023 & ~n42024;
  assign n7471 = n42030 | ~n42031;
  assign n42033 = P1_P2_EBX_REG_26_ & ~n41789;
  assign n42034 = ~n41574 & n41792;
  assign n42035 = P1_P2_EBX_REG_25_ & n42026;
  assign n42036 = ~P1_P2_EBX_REG_26_ & n42035;
  assign n42037 = P1_P2_EBX_REG_26_ & ~n42035;
  assign n42038 = ~n42036 & ~n42037;
  assign n42039 = n41790 & ~n42038;
  assign n42040 = ~n42033 & ~n42034;
  assign n7476 = n42039 | ~n42040;
  assign n42042 = P1_P2_EBX_REG_27_ & ~n41789;
  assign n42043 = ~n41622 & n41792;
  assign n42044 = P1_P2_EBX_REG_25_ & P1_P2_EBX_REG_26_;
  assign n42045 = n42026 & n42044;
  assign n42046 = P1_P2_EBX_REG_27_ & ~n42045;
  assign n42047 = ~P1_P2_EBX_REG_27_ & n42045;
  assign n42048 = ~n42046 & ~n42047;
  assign n42049 = n41790 & ~n42048;
  assign n42050 = ~n42042 & ~n42043;
  assign n7481 = n42049 | ~n42050;
  assign n42052 = P1_P2_EBX_REG_28_ & ~n41789;
  assign n42053 = ~n41671 & n41792;
  assign n42054 = P1_P2_EBX_REG_27_ & n42045;
  assign n42055 = ~P1_P2_EBX_REG_28_ & n42054;
  assign n42056 = P1_P2_EBX_REG_28_ & ~n42054;
  assign n42057 = ~n42055 & ~n42056;
  assign n42058 = n41790 & ~n42057;
  assign n42059 = ~n42052 & ~n42053;
  assign n7486 = n42058 | ~n42059;
  assign n42061 = P1_P2_EBX_REG_29_ & ~n41789;
  assign n42062 = ~n41719 & n41792;
  assign n42063 = P1_P2_EBX_REG_27_ & P1_P2_EBX_REG_28_;
  assign n42064 = n42045 & n42063;
  assign n42065 = P1_P2_EBX_REG_29_ & ~n42064;
  assign n42066 = ~P1_P2_EBX_REG_29_ & n42064;
  assign n42067 = ~n42065 & ~n42066;
  assign n42068 = n41790 & ~n42067;
  assign n42069 = ~n42061 & ~n42062;
  assign n7491 = n42068 | ~n42069;
  assign n42071 = P1_P2_EBX_REG_30_ & ~n41789;
  assign n42072 = ~n41768 & n41792;
  assign n42073 = P1_P2_EBX_REG_29_ & n42064;
  assign n42074 = ~P1_P2_EBX_REG_30_ & n42073;
  assign n42075 = P1_P2_EBX_REG_30_ & ~n42073;
  assign n42076 = ~n42074 & ~n42075;
  assign n42077 = n41790 & ~n42076;
  assign n42078 = ~n42071 & ~n42072;
  assign n7496 = n42077 | ~n42078;
  assign n42080 = P1_P2_EBX_REG_31_ & ~n41789;
  assign n42081 = P1_P2_EBX_REG_30_ & n42073;
  assign n42082 = ~P1_P2_EBX_REG_31_ & n42081;
  assign n42083 = P1_P2_EBX_REG_31_ & ~n42081;
  assign n42084 = ~n42082 & ~n42083;
  assign n42085 = n41790 & ~n42084;
  assign n7501 = n42080 | n42085;
  assign n42087 = ~n34946 & ~n34985;
  assign n42088 = ~n36621 & n42087;
  assign n42089 = n34813 & n34821;
  assign n42090 = n34935 & ~n42089;
  assign n42091 = n42088 & ~n42090;
  assign n42092 = P1_P2_STATE2_REG_2_ & ~n42091;
  assign n42093 = n34663 & n42092;
  assign n42094 = ~n34296 & n42093;
  assign n42095 = ~P1_P2_EBX_REG_31_ & n42094;
  assign n42096 = n34581 & n42092;
  assign n42097 = ~n34299 & n42096;
  assign n42098 = n34299 & n42096;
  assign n42099 = ~n34296 & n42098;
  assign n42100 = ~n42095 & ~n42097;
  assign n42101 = ~n42099 & n42100;
  assign n42102 = P1_P2_EBX_REG_0_ & ~n42101;
  assign n42103 = n34296 & n42098;
  assign n42104 = P1_P2_REIP_REG_0_ & n42103;
  assign n42105 = P1_P2_EBX_REG_31_ & n42094;
  assign n42106 = P1_P2_EBX_REG_0_ & n42105;
  assign n42107 = n34658 & n42092;
  assign n42108 = ~P1_P2_INSTQUEUERD_ADDR_REG_0_ & n42107;
  assign n42109 = n34654 & n42092;
  assign n42110 = ~P1_P2_INSTQUEUERD_ADDR_REG_0_ & n42109;
  assign n42111 = ~n42108 & ~n42110;
  assign n42112 = ~n42104 & ~n42106;
  assign n42113 = n42111 & n42112;
  assign n42114 = n34296 & n42093;
  assign n42115 = P1_P2_REIP_REG_0_ & n42114;
  assign n42116 = P1_P2_STATE2_REG_1_ & ~n42091;
  assign n42117 = n40204 & n42116;
  assign n42118 = P1_P2_PHYADDRPOINTER_REG_0_ & n42117;
  assign n42119 = P1_P2_REIP_REG_0_ & n42091;
  assign n42120 = P1_P2_STATE2_REG_3_ & ~n42091;
  assign n42121 = P1_P2_PHYADDRPOINTER_REG_0_ & n42120;
  assign n42122 = ~n42119 & ~n42121;
  assign n42123 = ~n40204 & n42116;
  assign n42124 = P1_P2_PHYADDRPOINTER_REG_0_ & n42123;
  assign n42125 = n42122 & ~n42124;
  assign n42126 = ~n42102 & n42113;
  assign n42127 = ~n42115 & n42126;
  assign n42128 = ~n42118 & n42127;
  assign n7506 = ~n42125 | ~n42128;
  assign n42130 = P1_P2_EBX_REG_1_ & ~n42101;
  assign n42131 = ~P1_P2_REIP_REG_1_ & n42103;
  assign n42132 = ~n41799 & n42105;
  assign n42133 = ~n34305 & ~n34310;
  assign n42134 = n42107 & ~n42133;
  assign n42135 = n42109 & ~n42133;
  assign n42136 = ~n42134 & ~n42135;
  assign n42137 = ~n42131 & ~n42132;
  assign n42138 = n42136 & n42137;
  assign n42139 = ~P1_P2_REIP_REG_1_ & n42114;
  assign n42140 = ~P1_P2_PHYADDRPOINTER_REG_1_ & n42117;
  assign n42141 = P1_P2_REIP_REG_1_ & n42091;
  assign n42142 = P1_P2_PHYADDRPOINTER_REG_1_ & n42120;
  assign n42143 = ~n42141 & ~n42142;
  assign n42144 = P1_P2_PHYADDRPOINTER_REG_0_ & P1_P2_PHYADDRPOINTER_REG_1_;
  assign n42145 = ~P1_P2_PHYADDRPOINTER_REG_0_ & ~P1_P2_PHYADDRPOINTER_REG_1_;
  assign n42146 = ~n42144 & ~n42145;
  assign n42147 = n42123 & ~n42146;
  assign n42148 = n42143 & ~n42147;
  assign n42149 = ~n42130 & n42138;
  assign n42150 = ~n42139 & n42149;
  assign n42151 = ~n42140 & n42150;
  assign n7511 = ~n42148 | ~n42151;
  assign n42153 = P1_P2_EBX_REG_2_ & ~n42101;
  assign n42154 = P1_P2_REIP_REG_1_ & ~P1_P2_REIP_REG_2_;
  assign n42155 = ~P1_P2_REIP_REG_1_ & P1_P2_REIP_REG_2_;
  assign n42156 = ~n42154 & ~n42155;
  assign n42157 = n42103 & ~n42156;
  assign n42158 = ~P1_P2_EBX_REG_0_ & ~P1_P2_EBX_REG_1_;
  assign n42159 = P1_P2_EBX_REG_2_ & ~n42158;
  assign n42160 = ~P1_P2_EBX_REG_2_ & n42158;
  assign n42161 = ~n42159 & ~n42160;
  assign n42162 = n42105 & n42161;
  assign n42163 = ~n34783 & n42107;
  assign n42164 = ~n34783 & n42109;
  assign n42165 = ~n42163 & ~n42164;
  assign n42166 = ~n42157 & ~n42162;
  assign n42167 = n42165 & n42166;
  assign n42168 = n42114 & ~n42156;
  assign n42169 = ~n39538 & n42117;
  assign n42170 = P1_P2_REIP_REG_2_ & n42091;
  assign n42171 = P1_P2_PHYADDRPOINTER_REG_2_ & n42120;
  assign n42172 = ~n42170 & ~n42171;
  assign n42173 = ~P1_P2_PHYADDRPOINTER_REG_0_ & P1_P2_PHYADDRPOINTER_REG_1_;
  assign n42174 = ~n39538 & ~n42173;
  assign n42175 = n39538 & n42173;
  assign n42176 = ~n42174 & ~n42175;
  assign n42177 = n42123 & n42176;
  assign n42178 = n42172 & ~n42177;
  assign n42179 = ~n42153 & n42167;
  assign n42180 = ~n42168 & n42179;
  assign n42181 = ~n42169 & n42180;
  assign n7516 = ~n42178 | ~n42181;
  assign n42183 = P1_P2_EBX_REG_3_ & ~n42101;
  assign n42184 = P1_P2_REIP_REG_1_ & P1_P2_REIP_REG_2_;
  assign n42185 = ~P1_P2_REIP_REG_3_ & n42184;
  assign n42186 = P1_P2_REIP_REG_3_ & ~n42184;
  assign n42187 = ~n42185 & ~n42186;
  assign n42188 = n42103 & ~n42187;
  assign n42189 = ~P1_P2_EBX_REG_3_ & n42160;
  assign n42190 = P1_P2_EBX_REG_3_ & ~n42160;
  assign n42191 = ~n42189 & ~n42190;
  assign n42192 = n42105 & n42191;
  assign n42193 = ~P1_P2_INSTQUEUERD_ADDR_REG_3_ & n34831;
  assign n42194 = ~n34832 & ~n42193;
  assign n42195 = n42107 & ~n42194;
  assign n42196 = n42109 & ~n42194;
  assign n42197 = ~n42195 & ~n42196;
  assign n42198 = ~n42188 & ~n42192;
  assign n42199 = n42197 & n42198;
  assign n42200 = n42114 & ~n42187;
  assign n42201 = ~n39560 & n42117;
  assign n42202 = P1_P2_REIP_REG_3_ & n42091;
  assign n42203 = P1_P2_PHYADDRPOINTER_REG_3_ & n42120;
  assign n42204 = ~n42202 & ~n42203;
  assign n42205 = n39560 & n42175;
  assign n42206 = ~n39560 & ~n42175;
  assign n42207 = ~n42205 & ~n42206;
  assign n42208 = n42123 & n42207;
  assign n42209 = n42204 & ~n42208;
  assign n42210 = ~n42183 & n42199;
  assign n42211 = ~n42200 & n42210;
  assign n42212 = ~n42201 & n42211;
  assign n7521 = ~n42209 | ~n42212;
  assign n42214 = P1_P2_INSTQUEUERD_ADDR_REG_3_ & n34831;
  assign n42215 = ~P1_P2_INSTQUEUERD_ADDR_REG_4_ & n42214;
  assign n42216 = P1_P2_INSTQUEUERD_ADDR_REG_4_ & ~n42214;
  assign n42217 = ~n42215 & ~n42216;
  assign n42218 = n42109 & ~n42217;
  assign n42219 = n42107 & ~n42217;
  assign n42220 = ~n42218 & ~n42219;
  assign n42221 = P1_P2_EBX_REG_4_ & ~n42101;
  assign n42222 = P1_P2_EBX_REG_4_ & ~n42189;
  assign n42223 = ~P1_P2_EBX_REG_3_ & ~P1_P2_EBX_REG_4_;
  assign n42224 = n42160 & n42223;
  assign n42225 = ~n42222 & ~n42224;
  assign n42226 = n42105 & n42225;
  assign n42227 = n36620 & ~n42091;
  assign n42228 = P1_P2_REIP_REG_3_ & n42184;
  assign n42229 = ~P1_P2_REIP_REG_4_ & n42228;
  assign n42230 = P1_P2_REIP_REG_4_ & ~n42228;
  assign n42231 = ~n42229 & ~n42230;
  assign n42232 = n42103 & ~n42231;
  assign n42233 = ~n42226 & ~n42227;
  assign n42234 = ~n42232 & n42233;
  assign n42235 = n42114 & ~n42231;
  assign n42236 = ~n39581 & n42117;
  assign n42237 = n42220 & ~n42221;
  assign n42238 = n42234 & n42237;
  assign n42239 = ~n42235 & n42238;
  assign n42240 = ~n42236 & n42239;
  assign n42241 = P1_P2_REIP_REG_4_ & n42091;
  assign n42242 = P1_P2_PHYADDRPOINTER_REG_4_ & n42120;
  assign n42243 = ~n42241 & ~n42242;
  assign n42244 = ~n39581 & ~n42205;
  assign n42245 = n39560 & n39581;
  assign n42246 = n42175 & n42245;
  assign n42247 = ~n42244 & ~n42246;
  assign n42248 = n42123 & n42247;
  assign n42249 = n42243 & ~n42248;
  assign n7526 = ~n42240 | ~n42249;
  assign n42251 = P1_P2_INSTQUEUERD_ADDR_REG_4_ & n42214;
  assign n42252 = n42109 & n42251;
  assign n42253 = n42107 & n42251;
  assign n42254 = ~n42252 & ~n42253;
  assign n42255 = P1_P2_EBX_REG_5_ & ~n42101;
  assign n42256 = ~P1_P2_EBX_REG_5_ & n42224;
  assign n42257 = P1_P2_EBX_REG_5_ & ~n42224;
  assign n42258 = ~n42256 & ~n42257;
  assign n42259 = n42105 & n42258;
  assign n42260 = P1_P2_REIP_REG_4_ & n42228;
  assign n42261 = ~P1_P2_REIP_REG_5_ & n42260;
  assign n42262 = P1_P2_REIP_REG_5_ & ~n42260;
  assign n42263 = ~n42261 & ~n42262;
  assign n42264 = n42103 & ~n42263;
  assign n42265 = ~n42227 & ~n42259;
  assign n42266 = ~n42264 & n42265;
  assign n42267 = n42114 & ~n42263;
  assign n42268 = ~n39604 & n42117;
  assign n42269 = n42254 & ~n42255;
  assign n42270 = n42266 & n42269;
  assign n42271 = ~n42267 & n42270;
  assign n42272 = ~n42268 & n42271;
  assign n42273 = P1_P2_REIP_REG_5_ & n42091;
  assign n42274 = P1_P2_PHYADDRPOINTER_REG_5_ & n42120;
  assign n42275 = ~n42273 & ~n42274;
  assign n42276 = n39604 & n42246;
  assign n42277 = ~n39604 & ~n42246;
  assign n42278 = ~n42276 & ~n42277;
  assign n42279 = n42123 & n42278;
  assign n42280 = n42275 & ~n42279;
  assign n7531 = ~n42272 | ~n42280;
  assign n42282 = P1_P2_REIP_REG_5_ & n42260;
  assign n42283 = ~P1_P2_REIP_REG_6_ & n42282;
  assign n42284 = P1_P2_REIP_REG_6_ & ~n42282;
  assign n42285 = ~n42283 & ~n42284;
  assign n42286 = n42114 & ~n42285;
  assign n42287 = P1_P2_EBX_REG_6_ & ~n42101;
  assign n42288 = P1_P2_EBX_REG_6_ & ~n42256;
  assign n42289 = ~P1_P2_EBX_REG_5_ & ~P1_P2_EBX_REG_6_;
  assign n42290 = n42224 & n42289;
  assign n42291 = ~n42288 & ~n42290;
  assign n42292 = n42105 & n42291;
  assign n42293 = n42103 & ~n42285;
  assign n42294 = ~n42227 & ~n42292;
  assign n42295 = ~n42293 & n42294;
  assign n42296 = ~n39627 & ~n42276;
  assign n42297 = n39604 & n39627;
  assign n42298 = n42246 & n42297;
  assign n42299 = ~n42296 & ~n42298;
  assign n42300 = n42123 & n42299;
  assign n42301 = P1_P2_REIP_REG_6_ & n42091;
  assign n42302 = P1_P2_PHYADDRPOINTER_REG_6_ & n42120;
  assign n42303 = ~n42301 & ~n42302;
  assign n42304 = ~n39627 & n42117;
  assign n42305 = n42303 & ~n42304;
  assign n42306 = ~n42286 & ~n42287;
  assign n42307 = n42295 & n42306;
  assign n42308 = ~n42300 & n42307;
  assign n7536 = ~n42305 | ~n42308;
  assign n42310 = P1_P2_REIP_REG_6_ & n42282;
  assign n42311 = ~P1_P2_REIP_REG_7_ & n42310;
  assign n42312 = P1_P2_REIP_REG_7_ & ~n42310;
  assign n42313 = ~n42311 & ~n42312;
  assign n42314 = n42114 & ~n42313;
  assign n42315 = P1_P2_EBX_REG_7_ & ~n42101;
  assign n42316 = ~P1_P2_EBX_REG_7_ & n42290;
  assign n42317 = P1_P2_EBX_REG_7_ & ~n42290;
  assign n42318 = ~n42316 & ~n42317;
  assign n42319 = n42105 & n42318;
  assign n42320 = n42103 & ~n42313;
  assign n42321 = ~n42227 & ~n42319;
  assign n42322 = ~n42320 & n42321;
  assign n42323 = n39650 & n42298;
  assign n42324 = ~n39650 & ~n42298;
  assign n42325 = ~n42323 & ~n42324;
  assign n42326 = n42123 & n42325;
  assign n42327 = P1_P2_REIP_REG_7_ & n42091;
  assign n42328 = P1_P2_PHYADDRPOINTER_REG_7_ & n42120;
  assign n42329 = ~n42327 & ~n42328;
  assign n42330 = ~n39650 & n42117;
  assign n42331 = n42329 & ~n42330;
  assign n42332 = ~n42314 & ~n42315;
  assign n42333 = n42322 & n42332;
  assign n42334 = ~n42326 & n42333;
  assign n7541 = ~n42331 | ~n42334;
  assign n42336 = P1_P2_REIP_REG_7_ & n42310;
  assign n42337 = ~P1_P2_REIP_REG_8_ & n42336;
  assign n42338 = P1_P2_REIP_REG_8_ & ~n42336;
  assign n42339 = ~n42337 & ~n42338;
  assign n42340 = n42114 & ~n42339;
  assign n42341 = P1_P2_EBX_REG_8_ & ~n42101;
  assign n42342 = P1_P2_EBX_REG_8_ & ~n42316;
  assign n42343 = ~P1_P2_EBX_REG_7_ & ~P1_P2_EBX_REG_8_;
  assign n42344 = n42290 & n42343;
  assign n42345 = ~n42342 & ~n42344;
  assign n42346 = n42105 & n42345;
  assign n42347 = n42103 & ~n42339;
  assign n42348 = ~n42227 & ~n42346;
  assign n42349 = ~n42347 & n42348;
  assign n42350 = ~n39673 & ~n42323;
  assign n42351 = n39650 & n39673;
  assign n42352 = n42298 & n42351;
  assign n42353 = ~n42350 & ~n42352;
  assign n42354 = n42123 & n42353;
  assign n42355 = P1_P2_REIP_REG_8_ & n42091;
  assign n42356 = P1_P2_PHYADDRPOINTER_REG_8_ & n42120;
  assign n42357 = ~n42355 & ~n42356;
  assign n42358 = ~n39673 & n42117;
  assign n42359 = n42357 & ~n42358;
  assign n42360 = ~n42340 & ~n42341;
  assign n42361 = n42349 & n42360;
  assign n42362 = ~n42354 & n42361;
  assign n7546 = ~n42359 | ~n42362;
  assign n42364 = P1_P2_REIP_REG_8_ & n42336;
  assign n42365 = ~P1_P2_REIP_REG_9_ & n42364;
  assign n42366 = P1_P2_REIP_REG_9_ & ~n42364;
  assign n42367 = ~n42365 & ~n42366;
  assign n42368 = n42114 & ~n42367;
  assign n42369 = P1_P2_EBX_REG_9_ & ~n42101;
  assign n42370 = ~P1_P2_EBX_REG_9_ & n42344;
  assign n42371 = P1_P2_EBX_REG_9_ & ~n42344;
  assign n42372 = ~n42370 & ~n42371;
  assign n42373 = n42105 & n42372;
  assign n42374 = n42103 & ~n42367;
  assign n42375 = ~n42227 & ~n42373;
  assign n42376 = ~n42374 & n42375;
  assign n42377 = n39696 & n42352;
  assign n42378 = ~n39696 & ~n42352;
  assign n42379 = ~n42377 & ~n42378;
  assign n42380 = n42123 & n42379;
  assign n42381 = P1_P2_REIP_REG_9_ & n42091;
  assign n42382 = P1_P2_PHYADDRPOINTER_REG_9_ & n42120;
  assign n42383 = ~n42381 & ~n42382;
  assign n42384 = ~n39696 & n42117;
  assign n42385 = n42383 & ~n42384;
  assign n42386 = ~n42368 & ~n42369;
  assign n42387 = n42376 & n42386;
  assign n42388 = ~n42380 & n42387;
  assign n7551 = ~n42385 | ~n42388;
  assign n42390 = P1_P2_REIP_REG_9_ & n42364;
  assign n42391 = ~P1_P2_REIP_REG_10_ & n42390;
  assign n42392 = P1_P2_REIP_REG_10_ & ~n42390;
  assign n42393 = ~n42391 & ~n42392;
  assign n42394 = n42114 & ~n42393;
  assign n42395 = P1_P2_EBX_REG_10_ & ~n42101;
  assign n42396 = P1_P2_EBX_REG_10_ & ~n42370;
  assign n42397 = ~P1_P2_EBX_REG_9_ & ~P1_P2_EBX_REG_10_;
  assign n42398 = n42344 & n42397;
  assign n42399 = ~n42396 & ~n42398;
  assign n42400 = n42105 & n42399;
  assign n42401 = n42103 & ~n42393;
  assign n42402 = ~n42227 & ~n42400;
  assign n42403 = ~n42401 & n42402;
  assign n42404 = ~n39719 & ~n42377;
  assign n42405 = n39696 & n39719;
  assign n42406 = n42352 & n42405;
  assign n42407 = ~n42404 & ~n42406;
  assign n42408 = n42123 & n42407;
  assign n42409 = P1_P2_REIP_REG_10_ & n42091;
  assign n42410 = P1_P2_PHYADDRPOINTER_REG_10_ & n42120;
  assign n42411 = ~n42409 & ~n42410;
  assign n42412 = ~n39719 & n42117;
  assign n42413 = n42411 & ~n42412;
  assign n42414 = ~n42394 & ~n42395;
  assign n42415 = n42403 & n42414;
  assign n42416 = ~n42408 & n42415;
  assign n7556 = ~n42413 | ~n42416;
  assign n42418 = P1_P2_REIP_REG_10_ & n42390;
  assign n42419 = ~P1_P2_REIP_REG_11_ & n42418;
  assign n42420 = P1_P2_REIP_REG_11_ & ~n42418;
  assign n42421 = ~n42419 & ~n42420;
  assign n42422 = n42114 & ~n42421;
  assign n42423 = P1_P2_EBX_REG_11_ & ~n42101;
  assign n42424 = ~P1_P2_EBX_REG_11_ & n42398;
  assign n42425 = P1_P2_EBX_REG_11_ & ~n42398;
  assign n42426 = ~n42424 & ~n42425;
  assign n42427 = n42105 & n42426;
  assign n42428 = n42103 & ~n42421;
  assign n42429 = ~n42227 & ~n42427;
  assign n42430 = ~n42428 & n42429;
  assign n42431 = n39742 & n42406;
  assign n42432 = ~n39742 & ~n42406;
  assign n42433 = ~n42431 & ~n42432;
  assign n42434 = n42123 & n42433;
  assign n42435 = P1_P2_REIP_REG_11_ & n42091;
  assign n42436 = P1_P2_PHYADDRPOINTER_REG_11_ & n42120;
  assign n42437 = ~n42435 & ~n42436;
  assign n42438 = ~n39742 & n42117;
  assign n42439 = n42437 & ~n42438;
  assign n42440 = ~n42422 & ~n42423;
  assign n42441 = n42430 & n42440;
  assign n42442 = ~n42434 & n42441;
  assign n7561 = ~n42439 | ~n42442;
  assign n42444 = P1_P2_REIP_REG_11_ & n42418;
  assign n42445 = ~P1_P2_REIP_REG_12_ & n42444;
  assign n42446 = P1_P2_REIP_REG_12_ & ~n42444;
  assign n42447 = ~n42445 & ~n42446;
  assign n42448 = n42114 & ~n42447;
  assign n42449 = P1_P2_EBX_REG_12_ & ~n42101;
  assign n42450 = P1_P2_EBX_REG_12_ & ~n42424;
  assign n42451 = ~P1_P2_EBX_REG_11_ & ~P1_P2_EBX_REG_12_;
  assign n42452 = n42398 & n42451;
  assign n42453 = ~n42450 & ~n42452;
  assign n42454 = n42105 & n42453;
  assign n42455 = n42103 & ~n42447;
  assign n42456 = ~n42227 & ~n42454;
  assign n42457 = ~n42455 & n42456;
  assign n42458 = ~n39765 & ~n42431;
  assign n42459 = n39742 & n39765;
  assign n42460 = n42406 & n42459;
  assign n42461 = ~n42458 & ~n42460;
  assign n42462 = n42123 & n42461;
  assign n42463 = P1_P2_REIP_REG_12_ & n42091;
  assign n42464 = P1_P2_PHYADDRPOINTER_REG_12_ & n42120;
  assign n42465 = ~n42463 & ~n42464;
  assign n42466 = ~n39765 & n42117;
  assign n42467 = n42465 & ~n42466;
  assign n42468 = ~n42448 & ~n42449;
  assign n42469 = n42457 & n42468;
  assign n42470 = ~n42462 & n42469;
  assign n7566 = ~n42467 | ~n42470;
  assign n42472 = P1_P2_REIP_REG_12_ & n42444;
  assign n42473 = ~P1_P2_REIP_REG_13_ & n42472;
  assign n42474 = P1_P2_REIP_REG_13_ & ~n42472;
  assign n42475 = ~n42473 & ~n42474;
  assign n42476 = n42114 & ~n42475;
  assign n42477 = P1_P2_EBX_REG_13_ & ~n42101;
  assign n42478 = ~P1_P2_EBX_REG_13_ & n42452;
  assign n42479 = P1_P2_EBX_REG_13_ & ~n42452;
  assign n42480 = ~n42478 & ~n42479;
  assign n42481 = n42105 & n42480;
  assign n42482 = n42103 & ~n42475;
  assign n42483 = ~n42227 & ~n42481;
  assign n42484 = ~n42482 & n42483;
  assign n42485 = n39788 & n42460;
  assign n42486 = ~n39788 & ~n42460;
  assign n42487 = ~n42485 & ~n42486;
  assign n42488 = n42123 & n42487;
  assign n42489 = P1_P2_REIP_REG_13_ & n42091;
  assign n42490 = P1_P2_PHYADDRPOINTER_REG_13_ & n42120;
  assign n42491 = ~n42489 & ~n42490;
  assign n42492 = ~n39788 & n42117;
  assign n42493 = n42491 & ~n42492;
  assign n42494 = ~n42476 & ~n42477;
  assign n42495 = n42484 & n42494;
  assign n42496 = ~n42488 & n42495;
  assign n7571 = ~n42493 | ~n42496;
  assign n42498 = P1_P2_REIP_REG_13_ & n42472;
  assign n42499 = ~P1_P2_REIP_REG_14_ & n42498;
  assign n42500 = P1_P2_REIP_REG_14_ & ~n42498;
  assign n42501 = ~n42499 & ~n42500;
  assign n42502 = n42114 & ~n42501;
  assign n42503 = P1_P2_EBX_REG_14_ & ~n42101;
  assign n42504 = P1_P2_EBX_REG_14_ & ~n42478;
  assign n42505 = ~P1_P2_EBX_REG_13_ & ~P1_P2_EBX_REG_14_;
  assign n42506 = n42452 & n42505;
  assign n42507 = ~n42504 & ~n42506;
  assign n42508 = n42105 & n42507;
  assign n42509 = n42103 & ~n42501;
  assign n42510 = ~n42227 & ~n42508;
  assign n42511 = ~n42509 & n42510;
  assign n42512 = ~n39811 & ~n42485;
  assign n42513 = n39788 & n39811;
  assign n42514 = n42460 & n42513;
  assign n42515 = ~n42512 & ~n42514;
  assign n42516 = n42123 & n42515;
  assign n42517 = P1_P2_REIP_REG_14_ & n42091;
  assign n42518 = P1_P2_PHYADDRPOINTER_REG_14_ & n42120;
  assign n42519 = ~n42517 & ~n42518;
  assign n42520 = ~n39811 & n42117;
  assign n42521 = n42519 & ~n42520;
  assign n42522 = ~n42502 & ~n42503;
  assign n42523 = n42511 & n42522;
  assign n42524 = ~n42516 & n42523;
  assign n7576 = ~n42521 | ~n42524;
  assign n42526 = P1_P2_REIP_REG_14_ & n42498;
  assign n42527 = ~P1_P2_REIP_REG_15_ & n42526;
  assign n42528 = P1_P2_REIP_REG_15_ & ~n42526;
  assign n42529 = ~n42527 & ~n42528;
  assign n42530 = n42114 & ~n42529;
  assign n42531 = P1_P2_EBX_REG_15_ & ~n42101;
  assign n42532 = ~P1_P2_EBX_REG_15_ & n42506;
  assign n42533 = P1_P2_EBX_REG_15_ & ~n42506;
  assign n42534 = ~n42532 & ~n42533;
  assign n42535 = n42105 & n42534;
  assign n42536 = n42103 & ~n42529;
  assign n42537 = ~n42227 & ~n42535;
  assign n42538 = ~n42536 & n42537;
  assign n42539 = n39834 & n42514;
  assign n42540 = ~n39834 & ~n42514;
  assign n42541 = ~n42539 & ~n42540;
  assign n42542 = n42123 & n42541;
  assign n42543 = P1_P2_REIP_REG_15_ & n42091;
  assign n42544 = P1_P2_PHYADDRPOINTER_REG_15_ & n42120;
  assign n42545 = ~n42543 & ~n42544;
  assign n42546 = ~n39834 & n42117;
  assign n42547 = n42545 & ~n42546;
  assign n42548 = ~n42530 & ~n42531;
  assign n42549 = n42538 & n42548;
  assign n42550 = ~n42542 & n42549;
  assign n7581 = ~n42547 | ~n42550;
  assign n42552 = P1_P2_REIP_REG_15_ & n42526;
  assign n42553 = ~P1_P2_REIP_REG_16_ & n42552;
  assign n42554 = P1_P2_REIP_REG_16_ & ~n42552;
  assign n42555 = ~n42553 & ~n42554;
  assign n42556 = n42114 & ~n42555;
  assign n42557 = P1_P2_EBX_REG_16_ & ~n42101;
  assign n42558 = P1_P2_EBX_REG_16_ & ~n42532;
  assign n42559 = ~P1_P2_EBX_REG_15_ & ~P1_P2_EBX_REG_16_;
  assign n42560 = n42506 & n42559;
  assign n42561 = ~n42558 & ~n42560;
  assign n42562 = n42105 & n42561;
  assign n42563 = n42103 & ~n42555;
  assign n42564 = ~n42227 & ~n42562;
  assign n42565 = ~n42563 & n42564;
  assign n42566 = ~n39857 & ~n42539;
  assign n42567 = n39834 & n39857;
  assign n42568 = n42514 & n42567;
  assign n42569 = ~n42566 & ~n42568;
  assign n42570 = n42123 & n42569;
  assign n42571 = P1_P2_REIP_REG_16_ & n42091;
  assign n42572 = P1_P2_PHYADDRPOINTER_REG_16_ & n42120;
  assign n42573 = ~n42571 & ~n42572;
  assign n42574 = ~n39857 & n42117;
  assign n42575 = n42573 & ~n42574;
  assign n42576 = ~n42556 & ~n42557;
  assign n42577 = n42565 & n42576;
  assign n42578 = ~n42570 & n42577;
  assign n7586 = ~n42575 | ~n42578;
  assign n42580 = P1_P2_REIP_REG_16_ & n42552;
  assign n42581 = ~P1_P2_REIP_REG_17_ & n42580;
  assign n42582 = P1_P2_REIP_REG_17_ & ~n42580;
  assign n42583 = ~n42581 & ~n42582;
  assign n42584 = n42114 & ~n42583;
  assign n42585 = P1_P2_EBX_REG_17_ & ~n42101;
  assign n42586 = ~P1_P2_EBX_REG_17_ & n42560;
  assign n42587 = P1_P2_EBX_REG_17_ & ~n42560;
  assign n42588 = ~n42586 & ~n42587;
  assign n42589 = n42105 & n42588;
  assign n42590 = n42103 & ~n42583;
  assign n42591 = ~n42227 & ~n42589;
  assign n42592 = ~n42590 & n42591;
  assign n42593 = n39880 & n42568;
  assign n42594 = ~n39880 & ~n42568;
  assign n42595 = ~n42593 & ~n42594;
  assign n42596 = n42123 & n42595;
  assign n42597 = P1_P2_REIP_REG_17_ & n42091;
  assign n42598 = P1_P2_PHYADDRPOINTER_REG_17_ & n42120;
  assign n42599 = ~n42597 & ~n42598;
  assign n42600 = ~n39880 & n42117;
  assign n42601 = n42599 & ~n42600;
  assign n42602 = ~n42584 & ~n42585;
  assign n42603 = n42592 & n42602;
  assign n42604 = ~n42596 & n42603;
  assign n7591 = ~n42601 | ~n42604;
  assign n42606 = P1_P2_REIP_REG_17_ & n42580;
  assign n42607 = ~P1_P2_REIP_REG_18_ & n42606;
  assign n42608 = P1_P2_REIP_REG_18_ & ~n42606;
  assign n42609 = ~n42607 & ~n42608;
  assign n42610 = n42114 & ~n42609;
  assign n42611 = P1_P2_EBX_REG_18_ & ~n42101;
  assign n42612 = P1_P2_EBX_REG_18_ & ~n42586;
  assign n42613 = ~P1_P2_EBX_REG_17_ & ~P1_P2_EBX_REG_18_;
  assign n42614 = n42560 & n42613;
  assign n42615 = ~n42612 & ~n42614;
  assign n42616 = n42105 & n42615;
  assign n42617 = n42103 & ~n42609;
  assign n42618 = ~n42227 & ~n42616;
  assign n42619 = ~n42617 & n42618;
  assign n42620 = ~n39903 & ~n42593;
  assign n42621 = n39880 & n39903;
  assign n42622 = n42568 & n42621;
  assign n42623 = ~n42620 & ~n42622;
  assign n42624 = n42123 & n42623;
  assign n42625 = P1_P2_REIP_REG_18_ & n42091;
  assign n42626 = P1_P2_PHYADDRPOINTER_REG_18_ & n42120;
  assign n42627 = ~n42625 & ~n42626;
  assign n42628 = ~n39903 & n42117;
  assign n42629 = n42627 & ~n42628;
  assign n42630 = ~n42610 & ~n42611;
  assign n42631 = n42619 & n42630;
  assign n42632 = ~n42624 & n42631;
  assign n7596 = ~n42629 | ~n42632;
  assign n42634 = P1_P2_REIP_REG_18_ & n42606;
  assign n42635 = ~P1_P2_REIP_REG_19_ & n42634;
  assign n42636 = P1_P2_REIP_REG_19_ & ~n42634;
  assign n42637 = ~n42635 & ~n42636;
  assign n42638 = n42114 & ~n42637;
  assign n42639 = P1_P2_EBX_REG_19_ & ~n42101;
  assign n42640 = ~P1_P2_EBX_REG_19_ & n42614;
  assign n42641 = P1_P2_EBX_REG_19_ & ~n42614;
  assign n42642 = ~n42640 & ~n42641;
  assign n42643 = n42105 & n42642;
  assign n42644 = n42103 & ~n42637;
  assign n42645 = ~n42227 & ~n42643;
  assign n42646 = ~n42644 & n42645;
  assign n42647 = n39926 & n42622;
  assign n42648 = ~n39926 & ~n42622;
  assign n42649 = ~n42647 & ~n42648;
  assign n42650 = n42123 & n42649;
  assign n42651 = P1_P2_REIP_REG_19_ & n42091;
  assign n42652 = P1_P2_PHYADDRPOINTER_REG_19_ & n42120;
  assign n42653 = ~n42651 & ~n42652;
  assign n42654 = ~n39926 & n42117;
  assign n42655 = n42653 & ~n42654;
  assign n42656 = ~n42638 & ~n42639;
  assign n42657 = n42646 & n42656;
  assign n42658 = ~n42650 & n42657;
  assign n7601 = ~n42655 | ~n42658;
  assign n42660 = P1_P2_REIP_REG_19_ & n42634;
  assign n42661 = ~P1_P2_REIP_REG_20_ & n42660;
  assign n42662 = P1_P2_REIP_REG_20_ & ~n42660;
  assign n42663 = ~n42661 & ~n42662;
  assign n42664 = n42114 & ~n42663;
  assign n42665 = P1_P2_EBX_REG_20_ & ~n42101;
  assign n42666 = n42103 & ~n42663;
  assign n42667 = P1_P2_EBX_REG_20_ & ~n42640;
  assign n42668 = ~P1_P2_EBX_REG_19_ & ~P1_P2_EBX_REG_20_;
  assign n42669 = n42614 & n42668;
  assign n42670 = ~n42667 & ~n42669;
  assign n42671 = n42105 & n42670;
  assign n42672 = ~n42666 & ~n42671;
  assign n42673 = ~n39949 & ~n42647;
  assign n42674 = n39926 & n39949;
  assign n42675 = n42622 & n42674;
  assign n42676 = ~n42673 & ~n42675;
  assign n42677 = n42123 & n42676;
  assign n42678 = P1_P2_REIP_REG_20_ & n42091;
  assign n42679 = P1_P2_PHYADDRPOINTER_REG_20_ & n42120;
  assign n42680 = ~n42678 & ~n42679;
  assign n42681 = ~n39949 & n42117;
  assign n42682 = n42680 & ~n42681;
  assign n42683 = ~n42664 & ~n42665;
  assign n42684 = n42672 & n42683;
  assign n42685 = ~n42677 & n42684;
  assign n7606 = ~n42682 | ~n42685;
  assign n42687 = P1_P2_REIP_REG_20_ & n42660;
  assign n42688 = ~P1_P2_REIP_REG_21_ & n42687;
  assign n42689 = P1_P2_REIP_REG_21_ & ~n42687;
  assign n42690 = ~n42688 & ~n42689;
  assign n42691 = n42114 & ~n42690;
  assign n42692 = P1_P2_EBX_REG_21_ & ~n42101;
  assign n42693 = n42103 & ~n42690;
  assign n42694 = ~P1_P2_EBX_REG_21_ & n42669;
  assign n42695 = P1_P2_EBX_REG_21_ & ~n42669;
  assign n42696 = ~n42694 & ~n42695;
  assign n42697 = n42105 & n42696;
  assign n42698 = ~n42693 & ~n42697;
  assign n42699 = n39972 & n42675;
  assign n42700 = ~n39972 & ~n42675;
  assign n42701 = ~n42699 & ~n42700;
  assign n42702 = n42123 & n42701;
  assign n42703 = P1_P2_REIP_REG_21_ & n42091;
  assign n42704 = P1_P2_PHYADDRPOINTER_REG_21_ & n42120;
  assign n42705 = ~n42703 & ~n42704;
  assign n42706 = ~n39972 & n42117;
  assign n42707 = n42705 & ~n42706;
  assign n42708 = ~n42691 & ~n42692;
  assign n42709 = n42698 & n42708;
  assign n42710 = ~n42702 & n42709;
  assign n7611 = ~n42707 | ~n42710;
  assign n42712 = P1_P2_REIP_REG_21_ & n42687;
  assign n42713 = ~P1_P2_REIP_REG_22_ & n42712;
  assign n42714 = P1_P2_REIP_REG_22_ & ~n42712;
  assign n42715 = ~n42713 & ~n42714;
  assign n42716 = n42114 & ~n42715;
  assign n42717 = P1_P2_EBX_REG_22_ & ~n42101;
  assign n42718 = n42103 & ~n42715;
  assign n42719 = P1_P2_EBX_REG_22_ & ~n42694;
  assign n42720 = ~P1_P2_EBX_REG_21_ & ~P1_P2_EBX_REG_22_;
  assign n42721 = n42669 & n42720;
  assign n42722 = ~n42719 & ~n42721;
  assign n42723 = n42105 & n42722;
  assign n42724 = ~n42718 & ~n42723;
  assign n42725 = ~n39996 & ~n42699;
  assign n42726 = n39972 & n39996;
  assign n42727 = n42675 & n42726;
  assign n42728 = ~n42725 & ~n42727;
  assign n42729 = n42123 & n42728;
  assign n42730 = P1_P2_REIP_REG_22_ & n42091;
  assign n42731 = P1_P2_PHYADDRPOINTER_REG_22_ & n42120;
  assign n42732 = ~n42730 & ~n42731;
  assign n42733 = ~n39996 & n42117;
  assign n42734 = n42732 & ~n42733;
  assign n42735 = ~n42716 & ~n42717;
  assign n42736 = n42724 & n42735;
  assign n42737 = ~n42729 & n42736;
  assign n7616 = ~n42734 | ~n42737;
  assign n42739 = P1_P2_REIP_REG_22_ & n42712;
  assign n42740 = ~P1_P2_REIP_REG_23_ & n42739;
  assign n42741 = P1_P2_REIP_REG_23_ & ~n42739;
  assign n42742 = ~n42740 & ~n42741;
  assign n42743 = n42114 & ~n42742;
  assign n42744 = P1_P2_EBX_REG_23_ & ~n42101;
  assign n42745 = n42103 & ~n42742;
  assign n42746 = ~P1_P2_EBX_REG_23_ & n42721;
  assign n42747 = P1_P2_EBX_REG_23_ & ~n42721;
  assign n42748 = ~n42746 & ~n42747;
  assign n42749 = n42105 & n42748;
  assign n42750 = ~n42745 & ~n42749;
  assign n42751 = n40019 & n42727;
  assign n42752 = ~n40019 & ~n42727;
  assign n42753 = ~n42751 & ~n42752;
  assign n42754 = n42123 & n42753;
  assign n42755 = P1_P2_REIP_REG_23_ & n42091;
  assign n42756 = P1_P2_PHYADDRPOINTER_REG_23_ & n42120;
  assign n42757 = ~n42755 & ~n42756;
  assign n42758 = ~n40019 & n42117;
  assign n42759 = n42757 & ~n42758;
  assign n42760 = ~n42743 & ~n42744;
  assign n42761 = n42750 & n42760;
  assign n42762 = ~n42754 & n42761;
  assign n7621 = ~n42759 | ~n42762;
  assign n42764 = P1_P2_REIP_REG_23_ & n42739;
  assign n42765 = ~P1_P2_REIP_REG_24_ & n42764;
  assign n42766 = P1_P2_REIP_REG_24_ & ~n42764;
  assign n42767 = ~n42765 & ~n42766;
  assign n42768 = n42114 & ~n42767;
  assign n42769 = P1_P2_EBX_REG_24_ & ~n42101;
  assign n42770 = n42103 & ~n42767;
  assign n42771 = P1_P2_EBX_REG_24_ & ~n42746;
  assign n42772 = ~P1_P2_EBX_REG_23_ & ~P1_P2_EBX_REG_24_;
  assign n42773 = n42721 & n42772;
  assign n42774 = ~n42771 & ~n42773;
  assign n42775 = n42105 & n42774;
  assign n42776 = ~n42770 & ~n42775;
  assign n42777 = ~n40042 & ~n42751;
  assign n42778 = n40019 & n40042;
  assign n42779 = n42727 & n42778;
  assign n42780 = ~n42777 & ~n42779;
  assign n42781 = n42123 & n42780;
  assign n42782 = P1_P2_REIP_REG_24_ & n42091;
  assign n42783 = P1_P2_PHYADDRPOINTER_REG_24_ & n42120;
  assign n42784 = ~n42782 & ~n42783;
  assign n42785 = ~n40042 & n42117;
  assign n42786 = n42784 & ~n42785;
  assign n42787 = ~n42768 & ~n42769;
  assign n42788 = n42776 & n42787;
  assign n42789 = ~n42781 & n42788;
  assign n7626 = ~n42786 | ~n42789;
  assign n42791 = P1_P2_REIP_REG_24_ & n42764;
  assign n42792 = ~P1_P2_REIP_REG_25_ & n42791;
  assign n42793 = P1_P2_REIP_REG_25_ & ~n42791;
  assign n42794 = ~n42792 & ~n42793;
  assign n42795 = n42114 & ~n42794;
  assign n42796 = P1_P2_EBX_REG_25_ & ~n42101;
  assign n42797 = n42103 & ~n42794;
  assign n42798 = ~P1_P2_EBX_REG_25_ & n42773;
  assign n42799 = P1_P2_EBX_REG_25_ & ~n42773;
  assign n42800 = ~n42798 & ~n42799;
  assign n42801 = n42105 & n42800;
  assign n42802 = ~n42797 & ~n42801;
  assign n42803 = n40065 & n42779;
  assign n42804 = ~n40065 & ~n42779;
  assign n42805 = ~n42803 & ~n42804;
  assign n42806 = n42123 & n42805;
  assign n42807 = P1_P2_REIP_REG_25_ & n42091;
  assign n42808 = P1_P2_PHYADDRPOINTER_REG_25_ & n42120;
  assign n42809 = ~n42807 & ~n42808;
  assign n42810 = ~n40065 & n42117;
  assign n42811 = n42809 & ~n42810;
  assign n42812 = ~n42795 & ~n42796;
  assign n42813 = n42802 & n42812;
  assign n42814 = ~n42806 & n42813;
  assign n7631 = ~n42811 | ~n42814;
  assign n42816 = P1_P2_REIP_REG_25_ & n42791;
  assign n42817 = ~P1_P2_REIP_REG_26_ & n42816;
  assign n42818 = P1_P2_REIP_REG_26_ & ~n42816;
  assign n42819 = ~n42817 & ~n42818;
  assign n42820 = n42114 & ~n42819;
  assign n42821 = P1_P2_EBX_REG_26_ & ~n42101;
  assign n42822 = n42103 & ~n42819;
  assign n42823 = P1_P2_EBX_REG_26_ & ~n42798;
  assign n42824 = ~P1_P2_EBX_REG_25_ & ~P1_P2_EBX_REG_26_;
  assign n42825 = n42773 & n42824;
  assign n42826 = ~n42823 & ~n42825;
  assign n42827 = n42105 & n42826;
  assign n42828 = ~n42822 & ~n42827;
  assign n42829 = ~n40088 & ~n42803;
  assign n42830 = n40065 & n40088;
  assign n42831 = n42779 & n42830;
  assign n42832 = ~n42829 & ~n42831;
  assign n42833 = n42123 & n42832;
  assign n42834 = P1_P2_REIP_REG_26_ & n42091;
  assign n42835 = P1_P2_PHYADDRPOINTER_REG_26_ & n42120;
  assign n42836 = ~n42834 & ~n42835;
  assign n42837 = ~n40088 & n42117;
  assign n42838 = n42836 & ~n42837;
  assign n42839 = ~n42820 & ~n42821;
  assign n42840 = n42828 & n42839;
  assign n42841 = ~n42833 & n42840;
  assign n7636 = ~n42838 | ~n42841;
  assign n42843 = P1_P2_REIP_REG_26_ & n42816;
  assign n42844 = ~P1_P2_REIP_REG_27_ & n42843;
  assign n42845 = P1_P2_REIP_REG_27_ & ~n42843;
  assign n42846 = ~n42844 & ~n42845;
  assign n42847 = n42114 & ~n42846;
  assign n42848 = P1_P2_EBX_REG_27_ & ~n42101;
  assign n42849 = n42103 & ~n42846;
  assign n42850 = ~P1_P2_EBX_REG_27_ & n42825;
  assign n42851 = P1_P2_EBX_REG_27_ & ~n42825;
  assign n42852 = ~n42850 & ~n42851;
  assign n42853 = n42105 & n42852;
  assign n42854 = ~n42849 & ~n42853;
  assign n42855 = n40111 & n42831;
  assign n42856 = ~n40111 & ~n42831;
  assign n42857 = ~n42855 & ~n42856;
  assign n42858 = n42123 & n42857;
  assign n42859 = P1_P2_REIP_REG_27_ & n42091;
  assign n42860 = P1_P2_PHYADDRPOINTER_REG_27_ & n42120;
  assign n42861 = ~n42859 & ~n42860;
  assign n42862 = ~n40111 & n42117;
  assign n42863 = n42861 & ~n42862;
  assign n42864 = ~n42847 & ~n42848;
  assign n42865 = n42854 & n42864;
  assign n42866 = ~n42858 & n42865;
  assign n7641 = ~n42863 | ~n42866;
  assign n42868 = P1_P2_REIP_REG_27_ & n42843;
  assign n42869 = ~P1_P2_REIP_REG_28_ & n42868;
  assign n42870 = P1_P2_REIP_REG_28_ & ~n42868;
  assign n42871 = ~n42869 & ~n42870;
  assign n42872 = n42114 & ~n42871;
  assign n42873 = P1_P2_EBX_REG_28_ & ~n42101;
  assign n42874 = n42103 & ~n42871;
  assign n42875 = P1_P2_EBX_REG_28_ & ~n42850;
  assign n42876 = ~P1_P2_EBX_REG_27_ & ~P1_P2_EBX_REG_28_;
  assign n42877 = n42825 & n42876;
  assign n42878 = ~n42875 & ~n42877;
  assign n42879 = n42105 & n42878;
  assign n42880 = ~n42874 & ~n42879;
  assign n42881 = ~n40135 & ~n42855;
  assign n42882 = n40111 & n40135;
  assign n42883 = n42831 & n42882;
  assign n42884 = ~n42881 & ~n42883;
  assign n42885 = n42123 & n42884;
  assign n42886 = P1_P2_REIP_REG_28_ & n42091;
  assign n42887 = P1_P2_PHYADDRPOINTER_REG_28_ & n42120;
  assign n42888 = ~n42886 & ~n42887;
  assign n42889 = ~n40135 & n42117;
  assign n42890 = n42888 & ~n42889;
  assign n42891 = ~n42872 & ~n42873;
  assign n42892 = n42880 & n42891;
  assign n42893 = ~n42885 & n42892;
  assign n7646 = ~n42890 | ~n42893;
  assign n42895 = P1_P2_REIP_REG_28_ & n42868;
  assign n42896 = ~P1_P2_REIP_REG_29_ & n42895;
  assign n42897 = P1_P2_REIP_REG_29_ & ~n42895;
  assign n42898 = ~n42896 & ~n42897;
  assign n42899 = n42114 & ~n42898;
  assign n42900 = P1_P2_EBX_REG_29_ & ~n42101;
  assign n42901 = n42103 & ~n42898;
  assign n42902 = P1_P2_EBX_REG_29_ & ~n42877;
  assign n42903 = ~P1_P2_EBX_REG_29_ & n42877;
  assign n42904 = ~n42902 & ~n42903;
  assign n42905 = n42105 & n42904;
  assign n42906 = ~n42901 & ~n42905;
  assign n42907 = ~n40158 & ~n42883;
  assign n42908 = n40158 & n42883;
  assign n42909 = ~n42907 & ~n42908;
  assign n42910 = n42123 & n42909;
  assign n42911 = P1_P2_REIP_REG_29_ & n42091;
  assign n42912 = P1_P2_PHYADDRPOINTER_REG_29_ & n42120;
  assign n42913 = ~n42911 & ~n42912;
  assign n42914 = ~n40158 & n42117;
  assign n42915 = n42913 & ~n42914;
  assign n42916 = ~n42899 & ~n42900;
  assign n42917 = n42906 & n42916;
  assign n42918 = ~n42910 & n42917;
  assign n7651 = ~n42915 | ~n42918;
  assign n42920 = P1_P2_REIP_REG_29_ & n42895;
  assign n42921 = ~P1_P2_REIP_REG_30_ & n42920;
  assign n42922 = P1_P2_REIP_REG_30_ & ~n42920;
  assign n42923 = ~n42921 & ~n42922;
  assign n42924 = n42114 & ~n42923;
  assign n42925 = P1_P2_EBX_REG_30_ & ~n42101;
  assign n42926 = n42103 & ~n42923;
  assign n42927 = ~P1_P2_EBX_REG_30_ & n42903;
  assign n42928 = P1_P2_EBX_REG_30_ & ~n42903;
  assign n42929 = ~n42927 & ~n42928;
  assign n42930 = n42105 & n42929;
  assign n42931 = ~n42926 & ~n42930;
  assign n42932 = n40181 & n42908;
  assign n42933 = ~n40181 & ~n42908;
  assign n42934 = ~n42932 & ~n42933;
  assign n42935 = n42123 & n42934;
  assign n42936 = P1_P2_REIP_REG_30_ & n42091;
  assign n42937 = P1_P2_PHYADDRPOINTER_REG_30_ & n42120;
  assign n42938 = ~n42936 & ~n42937;
  assign n42939 = ~n40181 & n42117;
  assign n42940 = n42938 & ~n42939;
  assign n42941 = ~n42924 & ~n42925;
  assign n42942 = n42931 & n42941;
  assign n42943 = ~n42935 & n42942;
  assign n7656 = ~n42940 | ~n42943;
  assign n42945 = ~n40204 & n42932;
  assign n42946 = n40204 & ~n42932;
  assign n42947 = ~n42945 & ~n42946;
  assign n42948 = ~n40204 & n42117;
  assign n42949 = n42947 & ~n42948;
  assign n42950 = P1_P2_EBX_REG_31_ & ~n42101;
  assign n42951 = P1_P2_EBX_REG_31_ & n42927;
  assign n42952 = ~P1_P2_EBX_REG_31_ & ~n42927;
  assign n42953 = ~n42951 & ~n42952;
  assign n42954 = n42105 & ~n42953;
  assign n42955 = P1_P2_REIP_REG_30_ & n42920;
  assign n42956 = ~P1_P2_REIP_REG_31_ & n42955;
  assign n42957 = P1_P2_REIP_REG_31_ & ~n42955;
  assign n42958 = ~n42956 & ~n42957;
  assign n42959 = n42103 & ~n42958;
  assign n42960 = P1_P2_PHYADDRPOINTER_REG_31_ & n42120;
  assign n42961 = P1_P2_REIP_REG_31_ & n42091;
  assign n42962 = ~n42960 & ~n42961;
  assign n42963 = n42114 & ~n42958;
  assign n42964 = n42962 & ~n42963;
  assign n42965 = ~n42950 & ~n42954;
  assign n42966 = ~n42959 & n42965;
  assign n42967 = n42964 & n42966;
  assign n42968 = n42949 & n42967;
  assign n42969 = ~n42123 & ~n42948;
  assign n42970 = n42967 & n42969;
  assign n7661 = ~n42968 & ~n42970;
  assign n42972 = ~P1_P2_DATAWIDTH_REG_1_ & ~P1_P2_REIP_REG_1_;
  assign n42973 = ~P1_P2_DATAWIDTH_REG_30_ & ~P1_P2_DATAWIDTH_REG_31_;
  assign n42974 = P1_P2_DATAWIDTH_REG_0_ & P1_P2_DATAWIDTH_REG_1_;
  assign n42975 = ~P1_P2_DATAWIDTH_REG_28_ & ~P1_P2_DATAWIDTH_REG_29_;
  assign n42976 = ~P1_P2_DATAWIDTH_REG_26_ & ~P1_P2_DATAWIDTH_REG_27_;
  assign n42977 = n42973 & ~n42974;
  assign n42978 = n42975 & n42977;
  assign n42979 = n42976 & n42978;
  assign n42980 = ~P1_P2_DATAWIDTH_REG_22_ & ~P1_P2_DATAWIDTH_REG_23_;
  assign n42981 = ~P1_P2_DATAWIDTH_REG_24_ & n42980;
  assign n42982 = ~P1_P2_DATAWIDTH_REG_25_ & n42981;
  assign n42983 = ~P1_P2_DATAWIDTH_REG_18_ & ~P1_P2_DATAWIDTH_REG_19_;
  assign n42984 = ~P1_P2_DATAWIDTH_REG_20_ & n42983;
  assign n42985 = ~P1_P2_DATAWIDTH_REG_21_ & n42984;
  assign n42986 = n42982 & n42985;
  assign n42987 = ~P1_P2_DATAWIDTH_REG_14_ & ~P1_P2_DATAWIDTH_REG_15_;
  assign n42988 = ~P1_P2_DATAWIDTH_REG_16_ & n42987;
  assign n42989 = ~P1_P2_DATAWIDTH_REG_17_ & n42988;
  assign n42990 = ~P1_P2_DATAWIDTH_REG_10_ & ~P1_P2_DATAWIDTH_REG_11_;
  assign n42991 = ~P1_P2_DATAWIDTH_REG_12_ & n42990;
  assign n42992 = ~P1_P2_DATAWIDTH_REG_13_ & n42991;
  assign n42993 = n42989 & n42992;
  assign n42994 = ~P1_P2_DATAWIDTH_REG_6_ & ~P1_P2_DATAWIDTH_REG_7_;
  assign n42995 = ~P1_P2_DATAWIDTH_REG_8_ & n42994;
  assign n42996 = ~P1_P2_DATAWIDTH_REG_9_ & n42995;
  assign n42997 = ~P1_P2_DATAWIDTH_REG_2_ & ~P1_P2_DATAWIDTH_REG_3_;
  assign n42998 = ~P1_P2_DATAWIDTH_REG_4_ & n42997;
  assign n42999 = ~P1_P2_DATAWIDTH_REG_5_ & n42998;
  assign n43000 = n42996 & n42999;
  assign n43001 = n42979 & n42986;
  assign n43002 = n42993 & n43001;
  assign n43003 = n43000 & n43002;
  assign n43004 = n42972 & n43003;
  assign n43005 = P1_P2_BYTEENABLE_REG_3_ & ~n43003;
  assign n43006 = ~P1_P2_DATAWIDTH_REG_0_ & ~P1_P2_REIP_REG_0_;
  assign n43007 = ~P1_P2_DATAWIDTH_REG_1_ & n43006;
  assign n43008 = n43003 & n43007;
  assign n43009 = ~n43004 & ~n43005;
  assign n7666 = n43008 | ~n43009;
  assign n43011 = P1_P2_REIP_REG_0_ & P1_P2_REIP_REG_1_;
  assign n43012 = P1_P2_DATAWIDTH_REG_0_ & ~P1_P2_REIP_REG_0_;
  assign n43013 = ~P1_P2_DATAWIDTH_REG_0_ & ~P1_P2_DATAWIDTH_REG_1_;
  assign n43014 = ~n43012 & ~n43013;
  assign n43015 = ~P1_P2_REIP_REG_1_ & ~n43014;
  assign n43016 = ~n43011 & ~n43015;
  assign n43017 = n43003 & ~n43016;
  assign n43018 = P1_P2_BYTEENABLE_REG_2_ & ~n43003;
  assign n7671 = n43017 | n43018;
  assign n43020 = P1_P2_REIP_REG_1_ & n43003;
  assign n43021 = P1_P2_BYTEENABLE_REG_1_ & ~n43003;
  assign n43022 = ~n43020 & ~n43021;
  assign n7676 = n43008 | ~n43022;
  assign n43024 = ~P1_P2_REIP_REG_0_ & ~P1_P2_REIP_REG_1_;
  assign n43025 = n43003 & ~n43024;
  assign n43026 = P1_P2_BYTEENABLE_REG_0_ & ~n43003;
  assign n7681 = n43025 | n43026;
  assign n43028 = P1_P2_W_R_N_REG & ~n34039;
  assign n43029 = ~P1_P2_READREQUEST_REG & n34039;
  assign n7686 = n43028 | n43029;
  assign n43031 = n34703 & n34935;
  assign n43032 = ~n34651 & n34935;
  assign n43033 = P1_P2_FLUSH_REG & ~n43032;
  assign n7691 = n43031 | n43033;
  assign n43035 = P1_P2_MORE_REG & ~n43032;
  assign n43036 = ~n34697 & n43032;
  assign n7696 = n43035 | n43036;
  assign n43038 = BS & ~n34256;
  assign n43039 = P1_P2_STATEBS16_REG & n34256;
  assign n43040 = ~P1_P2_STATE_REG_0_ & n34211;
  assign n43041 = ~n43038 & ~n43039;
  assign n7701 = n43040 | ~n43041;
  assign n43043 = ~n34581 & ~n34654;
  assign n43044 = ~n34299 & ~n43043;
  assign n43045 = ~P1_P2_STATEBS16_REG & n34581;
  assign n43046 = ~n34208 & ~n43045;
  assign n43047 = P1_P2_STATE2_REG_2_ & ~n43044;
  assign n43048 = n43046 & n43047;
  assign n43049 = P1_P2_STATE2_REG_0_ & ~n43048;
  assign n43050 = ~n34951 & ~n43049;
  assign n43051 = ~n34208 & n34293;
  assign n43052 = ~n34941 & ~n43051;
  assign n43053 = ~P1_P2_STATE2_REG_0_ & ~n43052;
  assign n43054 = ~n35013 & ~n43053;
  assign n43055 = ~n42090 & n43054;
  assign n43056 = ~n43050 & ~n43055;
  assign n43057 = P1_P2_REQUESTPENDING_REG & n43055;
  assign n7706 = n43056 | n43057;
  assign n43059 = P1_P2_D_C_N_REG & ~n34039;
  assign n43060 = ~P1_P2_CODEFETCH_REG & n34039;
  assign n43061 = ~n43059 & ~n43060;
  assign n7711 = n43040 | ~n43061;
  assign n43063 = P1_P2_MEMORYFETCH_REG & n34039;
  assign n43064 = P1_P2_M_IO_N_REG & ~n34039;
  assign n7716 = n43063 | n43064;
  assign n43066 = P1_P2_STATE2_REG_0_ & n36620;
  assign n43067 = n34650 & n34935;
  assign n43068 = P1_P2_CODEFETCH_REG & ~n43067;
  assign n7721 = n43066 | n43068;
  assign n43070 = P1_P2_STATE_REG_0_ & P1_P2_ADS_N_REG;
  assign n7726 = ~n34256 | n43070;
  assign n43072 = P1_P2_STATE2_REG_2_ & ~n34663;
  assign n43073 = ~n34658 & n43072;
  assign n43074 = ~n36620 & ~n42090;
  assign n43075 = ~n43073 & ~n43074;
  assign n43076 = P1_P2_READREQUEST_REG & n43074;
  assign n7731 = n43075 | n43076;
  assign n43078 = P1_P2_STATE2_REG_2_ & n34580;
  assign n43079 = ~n43074 & ~n43078;
  assign n43080 = P1_P2_MEMORYFETCH_REG & n43074;
  assign n7736 = n43079 | n43080;
  assign n43082 = P1_P1_STATE_REG_1_ & ~P1_P1_STATE_REG_0_;
  assign n43083 = P1_P1_BYTEENABLE_REG_3_ & n43082;
  assign n43084 = P1_P1_BE_N_REG_3_ & ~n43082;
  assign n7741 = n43083 | n43084;
  assign n43086 = P1_P1_BYTEENABLE_REG_2_ & n43082;
  assign n43087 = P1_P1_BE_N_REG_2_ & ~n43082;
  assign n7746 = n43086 | n43087;
  assign n43089 = P1_P1_BYTEENABLE_REG_1_ & n43082;
  assign n43090 = P1_P1_BE_N_REG_1_ & ~n43082;
  assign n7751 = n43089 | n43090;
  assign n43092 = P1_P1_BYTEENABLE_REG_0_ & n43082;
  assign n43093 = P1_P1_BE_N_REG_0_ & ~n43082;
  assign n7756 = n43092 | n43093;
  assign n43095 = P1_P1_STATE_REG_2_ & n43082;
  assign n43096 = P1_P1_REIP_REG_30_ & n43095;
  assign n43097 = ~P1_P1_STATE_REG_2_ & n43082;
  assign n43098 = P1_P1_REIP_REG_31_ & n43097;
  assign n43099 = P1_P1_ADDRESS_REG_29_ & ~n43082;
  assign n43100 = ~n43096 & ~n43098;
  assign n7761 = n43099 | ~n43100;
  assign n43102 = P1_P1_REIP_REG_29_ & n43095;
  assign n43103 = P1_P1_REIP_REG_30_ & n43097;
  assign n43104 = P1_P1_ADDRESS_REG_28_ & ~n43082;
  assign n43105 = ~n43102 & ~n43103;
  assign n7766 = n43104 | ~n43105;
  assign n43107 = P1_P1_REIP_REG_28_ & n43095;
  assign n43108 = P1_P1_REIP_REG_29_ & n43097;
  assign n43109 = P1_P1_ADDRESS_REG_27_ & ~n43082;
  assign n43110 = ~n43107 & ~n43108;
  assign n7771 = n43109 | ~n43110;
  assign n43112 = P1_P1_REIP_REG_27_ & n43095;
  assign n43113 = P1_P1_REIP_REG_28_ & n43097;
  assign n43114 = P1_P1_ADDRESS_REG_26_ & ~n43082;
  assign n43115 = ~n43112 & ~n43113;
  assign n7776 = n43114 | ~n43115;
  assign n43117 = P1_P1_REIP_REG_26_ & n43095;
  assign n43118 = P1_P1_REIP_REG_27_ & n43097;
  assign n43119 = P1_P1_ADDRESS_REG_25_ & ~n43082;
  assign n43120 = ~n43117 & ~n43118;
  assign n7781 = n43119 | ~n43120;
  assign n43122 = P1_P1_REIP_REG_25_ & n43095;
  assign n43123 = P1_P1_REIP_REG_26_ & n43097;
  assign n43124 = P1_P1_ADDRESS_REG_24_ & ~n43082;
  assign n43125 = ~n43122 & ~n43123;
  assign n7786 = n43124 | ~n43125;
  assign n43127 = P1_P1_REIP_REG_24_ & n43095;
  assign n43128 = P1_P1_REIP_REG_25_ & n43097;
  assign n43129 = P1_P1_ADDRESS_REG_23_ & ~n43082;
  assign n43130 = ~n43127 & ~n43128;
  assign n7791 = n43129 | ~n43130;
  assign n43132 = P1_P1_REIP_REG_23_ & n43095;
  assign n43133 = P1_P1_REIP_REG_24_ & n43097;
  assign n43134 = P1_P1_ADDRESS_REG_22_ & ~n43082;
  assign n43135 = ~n43132 & ~n43133;
  assign n7796 = n43134 | ~n43135;
  assign n43137 = P1_P1_REIP_REG_22_ & n43095;
  assign n43138 = P1_P1_REIP_REG_23_ & n43097;
  assign n43139 = P1_P1_ADDRESS_REG_21_ & ~n43082;
  assign n43140 = ~n43137 & ~n43138;
  assign n7801 = n43139 | ~n43140;
  assign n43142 = P1_P1_REIP_REG_21_ & n43095;
  assign n43143 = P1_P1_REIP_REG_22_ & n43097;
  assign n43144 = P1_P1_ADDRESS_REG_20_ & ~n43082;
  assign n43145 = ~n43142 & ~n43143;
  assign n7806 = n43144 | ~n43145;
  assign n43147 = P1_P1_REIP_REG_20_ & n43095;
  assign n43148 = P1_P1_REIP_REG_21_ & n43097;
  assign n43149 = P1_P1_ADDRESS_REG_19_ & ~n43082;
  assign n43150 = ~n43147 & ~n43148;
  assign n7811 = n43149 | ~n43150;
  assign n43152 = P1_P1_REIP_REG_19_ & n43095;
  assign n43153 = P1_P1_REIP_REG_20_ & n43097;
  assign n43154 = P1_P1_ADDRESS_REG_18_ & ~n43082;
  assign n43155 = ~n43152 & ~n43153;
  assign n7816 = n43154 | ~n43155;
  assign n43157 = P1_P1_REIP_REG_18_ & n43095;
  assign n43158 = P1_P1_REIP_REG_19_ & n43097;
  assign n43159 = P1_P1_ADDRESS_REG_17_ & ~n43082;
  assign n43160 = ~n43157 & ~n43158;
  assign n7821 = n43159 | ~n43160;
  assign n43162 = P1_P1_REIP_REG_17_ & n43095;
  assign n43163 = P1_P1_REIP_REG_18_ & n43097;
  assign n43164 = P1_P1_ADDRESS_REG_16_ & ~n43082;
  assign n43165 = ~n43162 & ~n43163;
  assign n7826 = n43164 | ~n43165;
  assign n43167 = P1_P1_REIP_REG_16_ & n43095;
  assign n43168 = P1_P1_REIP_REG_17_ & n43097;
  assign n43169 = P1_P1_ADDRESS_REG_15_ & ~n43082;
  assign n43170 = ~n43167 & ~n43168;
  assign n7831 = n43169 | ~n43170;
  assign n43172 = P1_P1_REIP_REG_15_ & n43095;
  assign n43173 = P1_P1_REIP_REG_16_ & n43097;
  assign n43174 = P1_P1_ADDRESS_REG_14_ & ~n43082;
  assign n43175 = ~n43172 & ~n43173;
  assign n7836 = n43174 | ~n43175;
  assign n43177 = P1_P1_REIP_REG_14_ & n43095;
  assign n43178 = P1_P1_REIP_REG_15_ & n43097;
  assign n43179 = P1_P1_ADDRESS_REG_13_ & ~n43082;
  assign n43180 = ~n43177 & ~n43178;
  assign n7841 = n43179 | ~n43180;
  assign n43182 = P1_P1_REIP_REG_13_ & n43095;
  assign n43183 = P1_P1_REIP_REG_14_ & n43097;
  assign n43184 = P1_P1_ADDRESS_REG_12_ & ~n43082;
  assign n43185 = ~n43182 & ~n43183;
  assign n7846 = n43184 | ~n43185;
  assign n43187 = P1_P1_REIP_REG_12_ & n43095;
  assign n43188 = P1_P1_REIP_REG_13_ & n43097;
  assign n43189 = P1_P1_ADDRESS_REG_11_ & ~n43082;
  assign n43190 = ~n43187 & ~n43188;
  assign n7851 = n43189 | ~n43190;
  assign n43192 = P1_P1_REIP_REG_11_ & n43095;
  assign n43193 = P1_P1_REIP_REG_12_ & n43097;
  assign n43194 = P1_P1_ADDRESS_REG_10_ & ~n43082;
  assign n43195 = ~n43192 & ~n43193;
  assign n7856 = n43194 | ~n43195;
  assign n43197 = P1_P1_REIP_REG_10_ & n43095;
  assign n43198 = P1_P1_REIP_REG_11_ & n43097;
  assign n43199 = P1_P1_ADDRESS_REG_9_ & ~n43082;
  assign n43200 = ~n43197 & ~n43198;
  assign n7861 = n43199 | ~n43200;
  assign n43202 = P1_P1_REIP_REG_9_ & n43095;
  assign n43203 = P1_P1_REIP_REG_10_ & n43097;
  assign n43204 = P1_P1_ADDRESS_REG_8_ & ~n43082;
  assign n43205 = ~n43202 & ~n43203;
  assign n7866 = n43204 | ~n43205;
  assign n43207 = P1_P1_REIP_REG_8_ & n43095;
  assign n43208 = P1_P1_REIP_REG_9_ & n43097;
  assign n43209 = P1_P1_ADDRESS_REG_7_ & ~n43082;
  assign n43210 = ~n43207 & ~n43208;
  assign n7871 = n43209 | ~n43210;
  assign n43212 = P1_P1_REIP_REG_7_ & n43095;
  assign n43213 = P1_P1_REIP_REG_8_ & n43097;
  assign n43214 = P1_P1_ADDRESS_REG_6_ & ~n43082;
  assign n43215 = ~n43212 & ~n43213;
  assign n7876 = n43214 | ~n43215;
  assign n43217 = P1_P1_REIP_REG_6_ & n43095;
  assign n43218 = P1_P1_REIP_REG_7_ & n43097;
  assign n43219 = P1_P1_ADDRESS_REG_5_ & ~n43082;
  assign n43220 = ~n43217 & ~n43218;
  assign n7881 = n43219 | ~n43220;
  assign n43222 = P1_P1_REIP_REG_5_ & n43095;
  assign n43223 = P1_P1_REIP_REG_6_ & n43097;
  assign n43224 = P1_P1_ADDRESS_REG_4_ & ~n43082;
  assign n43225 = ~n43222 & ~n43223;
  assign n7886 = n43224 | ~n43225;
  assign n43227 = P1_P1_REIP_REG_4_ & n43095;
  assign n43228 = P1_P1_REIP_REG_5_ & n43097;
  assign n43229 = P1_P1_ADDRESS_REG_3_ & ~n43082;
  assign n43230 = ~n43227 & ~n43228;
  assign n7891 = n43229 | ~n43230;
  assign n43232 = P1_P1_REIP_REG_3_ & n43095;
  assign n43233 = P1_P1_REIP_REG_4_ & n43097;
  assign n43234 = P1_P1_ADDRESS_REG_2_ & ~n43082;
  assign n43235 = ~n43232 & ~n43233;
  assign n7896 = n43234 | ~n43235;
  assign n43237 = P1_P1_REIP_REG_2_ & n43095;
  assign n43238 = P1_P1_REIP_REG_3_ & n43097;
  assign n43239 = P1_P1_ADDRESS_REG_1_ & ~n43082;
  assign n43240 = ~n43237 & ~n43238;
  assign n7901 = n43239 | ~n43240;
  assign n43242 = P1_P1_REIP_REG_1_ & n43095;
  assign n43243 = P1_P1_REIP_REG_2_ & n43097;
  assign n43244 = P1_P1_ADDRESS_REG_0_ & ~n43082;
  assign n43245 = ~n43242 & ~n43243;
  assign n7906 = n43244 | ~n43245;
  assign n43247 = ~P1_P1_STATE_REG_2_ & P1_P1_STATE_REG_1_;
  assign n43248 = NA & n43247;
  assign n43249 = P1_P1_STATE_REG_0_ & ~n43248;
  assign n43250 = ~HOLD & ~P1_P1_REQUESTPENDING_REG;
  assign n43251 = P1_READY11_REG & P2_P1_ADS_N_REG;
  assign n43252 = ~n43250 & n43251;
  assign n43253 = n43247 & n43252;
  assign n43254 = ~P1_P1_STATE_REG_2_ & ~P1_P1_STATE_REG_1_;
  assign n43255 = HOLD & ~P1_P1_REQUESTPENDING_REG;
  assign n43256 = n43254 & n43255;
  assign n43257 = ~n43253 & ~n43256;
  assign n43258 = n43249 & ~n43257;
  assign n43259 = ~n43095 & ~n43258;
  assign n43260 = ~HOLD & P1_P1_REQUESTPENDING_REG;
  assign n43261 = P1_P1_STATE_REG_0_ & ~n43260;
  assign n43262 = ~n43250 & n43261;
  assign n43263 = ~NA & ~P1_P1_STATE_REG_0_;
  assign n43264 = n43250 & ~n43251;
  assign n43265 = ~n43251 & n43260;
  assign n43266 = P1_P1_STATE_REG_1_ & ~n43264;
  assign n43267 = ~n43265 & n43266;
  assign n43268 = ~n43262 & ~n43263;
  assign n43269 = ~n43267 & n43268;
  assign n43270 = P1_P1_STATE_REG_2_ & ~n43269;
  assign n7911 = ~n43259 | n43270;
  assign n43272 = P1_P1_STATE_REG_2_ & ~n43261;
  assign n43273 = P1_P1_STATE_REG_0_ & P1_P1_REQUESTPENDING_REG;
  assign n43274 = ~P1_P1_STATE_REG_2_ & n43273;
  assign n43275 = ~n43272 & ~n43274;
  assign n43276 = ~P1_P1_STATE_REG_1_ & ~n43275;
  assign n43277 = HOLD & ~n43251;
  assign n43278 = P1_P1_STATE_REG_0_ & ~n43277;
  assign n43279 = P1_P1_STATE_REG_2_ & ~n43278;
  assign n43280 = ~n43264 & ~n43279;
  assign n43281 = P1_P1_STATE_REG_1_ & n43280;
  assign n43282 = n43082 & n43251;
  assign n43283 = ~n43097 & ~n43282;
  assign n43284 = ~n43276 & ~n43281;
  assign n7916 = ~n43283 | ~n43284;
  assign n43286 = P1_P1_STATE_REG_1_ & ~n43265;
  assign n43287 = n43273 & ~n43286;
  assign n43288 = ~P1_P1_STATE_REG_2_ & ~n43287;
  assign n43289 = P1_P1_STATE_REG_2_ & n43261;
  assign n43290 = NA & ~P1_P1_STATE_REG_0_;
  assign n43291 = P1_P1_STATE_REG_2_ & ~n43260;
  assign n43292 = ~n43290 & ~n43291;
  assign n43293 = ~P1_P1_STATE_REG_1_ & ~n43292;
  assign n43294 = ~n43288 & ~n43289;
  assign n7921 = n43293 | ~n43294;
  assign n43296 = ~BS & ~n43254;
  assign n43297 = P1_P1_STATE_REG_0_ & n43247;
  assign n43298 = ~P1_P1_STATE_REG_1_ & ~P1_P1_STATE_REG_0_;
  assign n43299 = ~n43297 & ~n43298;
  assign n43300 = n43296 & ~n43299;
  assign n43301 = P1_P1_DATAWIDTH_REG_0_ & n43299;
  assign n7926 = n43300 | n43301;
  assign n43303 = P1_P1_DATAWIDTH_REG_1_ & n43299;
  assign n43304 = ~n43296 & ~n43299;
  assign n7931 = n43303 | n43304;
  assign n7936 = P1_P1_DATAWIDTH_REG_2_ & n43299;
  assign n7941 = P1_P1_DATAWIDTH_REG_3_ & n43299;
  assign n7946 = P1_P1_DATAWIDTH_REG_4_ & n43299;
  assign n7951 = P1_P1_DATAWIDTH_REG_5_ & n43299;
  assign n7956 = P1_P1_DATAWIDTH_REG_6_ & n43299;
  assign n7961 = P1_P1_DATAWIDTH_REG_7_ & n43299;
  assign n7966 = P1_P1_DATAWIDTH_REG_8_ & n43299;
  assign n7971 = P1_P1_DATAWIDTH_REG_9_ & n43299;
  assign n7976 = P1_P1_DATAWIDTH_REG_10_ & n43299;
  assign n7981 = P1_P1_DATAWIDTH_REG_11_ & n43299;
  assign n7986 = P1_P1_DATAWIDTH_REG_12_ & n43299;
  assign n7991 = P1_P1_DATAWIDTH_REG_13_ & n43299;
  assign n7996 = P1_P1_DATAWIDTH_REG_14_ & n43299;
  assign n8001 = P1_P1_DATAWIDTH_REG_15_ & n43299;
  assign n8006 = P1_P1_DATAWIDTH_REG_16_ & n43299;
  assign n8011 = P1_P1_DATAWIDTH_REG_17_ & n43299;
  assign n8016 = P1_P1_DATAWIDTH_REG_18_ & n43299;
  assign n8021 = P1_P1_DATAWIDTH_REG_19_ & n43299;
  assign n8026 = P1_P1_DATAWIDTH_REG_20_ & n43299;
  assign n8031 = P1_P1_DATAWIDTH_REG_21_ & n43299;
  assign n8036 = P1_P1_DATAWIDTH_REG_22_ & n43299;
  assign n8041 = P1_P1_DATAWIDTH_REG_23_ & n43299;
  assign n8046 = P1_P1_DATAWIDTH_REG_24_ & n43299;
  assign n8051 = P1_P1_DATAWIDTH_REG_25_ & n43299;
  assign n8056 = P1_P1_DATAWIDTH_REG_26_ & n43299;
  assign n8061 = P1_P1_DATAWIDTH_REG_27_ & n43299;
  assign n8066 = P1_P1_DATAWIDTH_REG_28_ & n43299;
  assign n8071 = P1_P1_DATAWIDTH_REG_29_ & n43299;
  assign n8076 = P1_P1_DATAWIDTH_REG_30_ & n43299;
  assign n8081 = P1_P1_DATAWIDTH_REG_31_ & n43299;
  assign n43336 = P1_P1_STATE2_REG_2_ & P1_P1_STATE2_REG_1_;
  assign n43337 = P1_P1_STATE2_REG_1_ & n43251;
  assign n43338 = ~P1_P1_STATE2_REG_0_ & ~n43337;
  assign n43339 = ~P1_P1_STATEBS16_REG & ~n43251;
  assign n43340 = P1_P1_STATE_REG_2_ & ~P1_P1_STATE_REG_1_;
  assign n43341 = ~n43247 & ~n43340;
  assign n43342 = ~P1_P1_STATE_REG_0_ & ~n43341;
  assign n43343 = n43339 & n43342;
  assign n43344 = P1_P1_INSTQUEUERD_ADDR_REG_1_ & P1_P1_INSTQUEUERD_ADDR_REG_0_;
  assign n43345 = ~P1_P1_INSTQUEUERD_ADDR_REG_2_ & n43344;
  assign n43346 = P1_P1_INSTQUEUERD_ADDR_REG_3_ & n43345;
  assign n43347 = P1_P1_INSTQUEUE_REG_11__5_ & n43346;
  assign n43348 = P1_P1_INSTQUEUERD_ADDR_REG_1_ & ~P1_P1_INSTQUEUERD_ADDR_REG_0_;
  assign n43349 = ~P1_P1_INSTQUEUERD_ADDR_REG_2_ & n43348;
  assign n43350 = P1_P1_INSTQUEUERD_ADDR_REG_3_ & n43349;
  assign n43351 = P1_P1_INSTQUEUE_REG_10__5_ & n43350;
  assign n43352 = ~n43347 & ~n43351;
  assign n43353 = ~P1_P1_INSTQUEUERD_ADDR_REG_1_ & P1_P1_INSTQUEUERD_ADDR_REG_0_;
  assign n43354 = ~P1_P1_INSTQUEUERD_ADDR_REG_2_ & n43353;
  assign n43355 = P1_P1_INSTQUEUERD_ADDR_REG_3_ & n43354;
  assign n43356 = P1_P1_INSTQUEUE_REG_9__5_ & n43355;
  assign n43357 = ~P1_P1_INSTQUEUERD_ADDR_REG_1_ & ~P1_P1_INSTQUEUERD_ADDR_REG_0_;
  assign n43358 = ~P1_P1_INSTQUEUERD_ADDR_REG_2_ & n43357;
  assign n43359 = P1_P1_INSTQUEUERD_ADDR_REG_3_ & n43358;
  assign n43360 = P1_P1_INSTQUEUE_REG_8__5_ & n43359;
  assign n43361 = ~n43356 & ~n43360;
  assign n43362 = P1_P1_INSTQUEUERD_ADDR_REG_3_ & P1_P1_INSTQUEUERD_ADDR_REG_2_;
  assign n43363 = n43344 & n43362;
  assign n43364 = P1_P1_INSTQUEUE_REG_15__5_ & n43363;
  assign n43365 = n43348 & n43362;
  assign n43366 = P1_P1_INSTQUEUE_REG_14__5_ & n43365;
  assign n43367 = n43353 & n43362;
  assign n43368 = P1_P1_INSTQUEUE_REG_13__5_ & n43367;
  assign n43369 = n43357 & n43362;
  assign n43370 = P1_P1_INSTQUEUE_REG_12__5_ & n43369;
  assign n43371 = ~n43364 & ~n43366;
  assign n43372 = ~n43368 & n43371;
  assign n43373 = ~n43370 & n43372;
  assign n43374 = ~P1_P1_INSTQUEUERD_ADDR_REG_3_ & P1_P1_INSTQUEUERD_ADDR_REG_2_;
  assign n43375 = n43344 & n43374;
  assign n43376 = P1_P1_INSTQUEUE_REG_7__5_ & n43375;
  assign n43377 = n43348 & n43374;
  assign n43378 = P1_P1_INSTQUEUE_REG_6__5_ & n43377;
  assign n43379 = n43353 & n43374;
  assign n43380 = P1_P1_INSTQUEUE_REG_5__5_ & n43379;
  assign n43381 = n43357 & n43374;
  assign n43382 = P1_P1_INSTQUEUE_REG_4__5_ & n43381;
  assign n43383 = ~n43376 & ~n43378;
  assign n43384 = ~n43380 & n43383;
  assign n43385 = ~n43382 & n43384;
  assign n43386 = ~P1_P1_INSTQUEUERD_ADDR_REG_3_ & n43345;
  assign n43387 = P1_P1_INSTQUEUE_REG_3__5_ & n43386;
  assign n43388 = ~P1_P1_INSTQUEUERD_ADDR_REG_3_ & ~P1_P1_INSTQUEUERD_ADDR_REG_2_;
  assign n43389 = n43348 & n43388;
  assign n43390 = P1_P1_INSTQUEUE_REG_2__5_ & n43389;
  assign n43391 = n43353 & n43388;
  assign n43392 = P1_P1_INSTQUEUE_REG_1__5_ & n43391;
  assign n43393 = ~P1_P1_INSTQUEUERD_ADDR_REG_3_ & n43358;
  assign n43394 = P1_P1_INSTQUEUE_REG_0__5_ & n43393;
  assign n43395 = ~n43387 & ~n43390;
  assign n43396 = ~n43392 & n43395;
  assign n43397 = ~n43394 & n43396;
  assign n43398 = n43352 & n43361;
  assign n43399 = n43373 & n43398;
  assign n43400 = n43385 & n43399;
  assign n43401 = n43397 & n43400;
  assign n43402 = P1_P1_INSTQUEUE_REG_11__6_ & n43346;
  assign n43403 = P1_P1_INSTQUEUE_REG_10__6_ & n43350;
  assign n43404 = ~n43402 & ~n43403;
  assign n43405 = P1_P1_INSTQUEUE_REG_9__6_ & n43355;
  assign n43406 = P1_P1_INSTQUEUE_REG_8__6_ & n43359;
  assign n43407 = ~n43405 & ~n43406;
  assign n43408 = P1_P1_INSTQUEUE_REG_15__6_ & n43363;
  assign n43409 = P1_P1_INSTQUEUE_REG_14__6_ & n43365;
  assign n43410 = P1_P1_INSTQUEUE_REG_13__6_ & n43367;
  assign n43411 = P1_P1_INSTQUEUE_REG_12__6_ & n43369;
  assign n43412 = ~n43408 & ~n43409;
  assign n43413 = ~n43410 & n43412;
  assign n43414 = ~n43411 & n43413;
  assign n43415 = P1_P1_INSTQUEUE_REG_7__6_ & n43375;
  assign n43416 = P1_P1_INSTQUEUE_REG_6__6_ & n43377;
  assign n43417 = P1_P1_INSTQUEUE_REG_5__6_ & n43379;
  assign n43418 = P1_P1_INSTQUEUE_REG_4__6_ & n43381;
  assign n43419 = ~n43415 & ~n43416;
  assign n43420 = ~n43417 & n43419;
  assign n43421 = ~n43418 & n43420;
  assign n43422 = P1_P1_INSTQUEUE_REG_3__6_ & n43386;
  assign n43423 = P1_P1_INSTQUEUE_REG_2__6_ & n43389;
  assign n43424 = P1_P1_INSTQUEUE_REG_1__6_ & n43391;
  assign n43425 = P1_P1_INSTQUEUE_REG_0__6_ & n43393;
  assign n43426 = ~n43422 & ~n43423;
  assign n43427 = ~n43424 & n43426;
  assign n43428 = ~n43425 & n43427;
  assign n43429 = n43404 & n43407;
  assign n43430 = n43414 & n43429;
  assign n43431 = n43421 & n43430;
  assign n43432 = n43428 & n43431;
  assign n43433 = n43401 & n43432;
  assign n43434 = P1_P1_INSTQUEUE_REG_11__4_ & n43346;
  assign n43435 = P1_P1_INSTQUEUE_REG_10__4_ & n43350;
  assign n43436 = ~n43434 & ~n43435;
  assign n43437 = P1_P1_INSTQUEUE_REG_9__4_ & n43355;
  assign n43438 = P1_P1_INSTQUEUE_REG_8__4_ & n43359;
  assign n43439 = ~n43437 & ~n43438;
  assign n43440 = P1_P1_INSTQUEUE_REG_15__4_ & n43363;
  assign n43441 = P1_P1_INSTQUEUE_REG_14__4_ & n43365;
  assign n43442 = P1_P1_INSTQUEUE_REG_13__4_ & n43367;
  assign n43443 = P1_P1_INSTQUEUE_REG_12__4_ & n43369;
  assign n43444 = ~n43440 & ~n43441;
  assign n43445 = ~n43442 & n43444;
  assign n43446 = ~n43443 & n43445;
  assign n43447 = P1_P1_INSTQUEUE_REG_7__4_ & n43375;
  assign n43448 = P1_P1_INSTQUEUE_REG_6__4_ & n43377;
  assign n43449 = P1_P1_INSTQUEUE_REG_5__4_ & n43379;
  assign n43450 = P1_P1_INSTQUEUE_REG_4__4_ & n43381;
  assign n43451 = ~n43447 & ~n43448;
  assign n43452 = ~n43449 & n43451;
  assign n43453 = ~n43450 & n43452;
  assign n43454 = P1_P1_INSTQUEUE_REG_3__4_ & n43386;
  assign n43455 = P1_P1_INSTQUEUE_REG_2__4_ & n43389;
  assign n43456 = P1_P1_INSTQUEUE_REG_1__4_ & n43391;
  assign n43457 = P1_P1_INSTQUEUE_REG_0__4_ & n43393;
  assign n43458 = ~n43454 & ~n43455;
  assign n43459 = ~n43456 & n43458;
  assign n43460 = ~n43457 & n43459;
  assign n43461 = n43436 & n43439;
  assign n43462 = n43446 & n43461;
  assign n43463 = n43453 & n43462;
  assign n43464 = n43460 & n43463;
  assign n43465 = P1_P1_INSTQUEUE_REG_11__7_ & n43346;
  assign n43466 = P1_P1_INSTQUEUE_REG_10__7_ & n43350;
  assign n43467 = ~n43465 & ~n43466;
  assign n43468 = P1_P1_INSTQUEUE_REG_9__7_ & n43355;
  assign n43469 = P1_P1_INSTQUEUE_REG_8__7_ & n43359;
  assign n43470 = ~n43468 & ~n43469;
  assign n43471 = P1_P1_INSTQUEUE_REG_15__7_ & n43363;
  assign n43472 = P1_P1_INSTQUEUE_REG_14__7_ & n43365;
  assign n43473 = P1_P1_INSTQUEUE_REG_13__7_ & n43367;
  assign n43474 = P1_P1_INSTQUEUE_REG_12__7_ & n43369;
  assign n43475 = ~n43471 & ~n43472;
  assign n43476 = ~n43473 & n43475;
  assign n43477 = ~n43474 & n43476;
  assign n43478 = P1_P1_INSTQUEUE_REG_7__7_ & n43375;
  assign n43479 = P1_P1_INSTQUEUE_REG_6__7_ & n43377;
  assign n43480 = P1_P1_INSTQUEUE_REG_5__7_ & n43379;
  assign n43481 = P1_P1_INSTQUEUE_REG_4__7_ & n43381;
  assign n43482 = ~n43478 & ~n43479;
  assign n43483 = ~n43480 & n43482;
  assign n43484 = ~n43481 & n43483;
  assign n43485 = P1_P1_INSTQUEUE_REG_3__7_ & n43386;
  assign n43486 = P1_P1_INSTQUEUE_REG_2__7_ & n43389;
  assign n43487 = P1_P1_INSTQUEUE_REG_1__7_ & n43391;
  assign n43488 = P1_P1_INSTQUEUE_REG_0__7_ & n43393;
  assign n43489 = ~n43485 & ~n43486;
  assign n43490 = ~n43487 & n43489;
  assign n43491 = ~n43488 & n43490;
  assign n43492 = n43467 & n43470;
  assign n43493 = n43477 & n43492;
  assign n43494 = n43484 & n43493;
  assign n43495 = n43491 & n43494;
  assign n43496 = P1_P1_INSTQUEUE_REG_11__3_ & n43346;
  assign n43497 = P1_P1_INSTQUEUE_REG_10__3_ & n43350;
  assign n43498 = ~n43496 & ~n43497;
  assign n43499 = P1_P1_INSTQUEUE_REG_9__3_ & n43355;
  assign n43500 = P1_P1_INSTQUEUE_REG_8__3_ & n43359;
  assign n43501 = ~n43499 & ~n43500;
  assign n43502 = P1_P1_INSTQUEUE_REG_15__3_ & n43363;
  assign n43503 = P1_P1_INSTQUEUE_REG_14__3_ & n43365;
  assign n43504 = P1_P1_INSTQUEUE_REG_13__3_ & n43367;
  assign n43505 = P1_P1_INSTQUEUE_REG_12__3_ & n43369;
  assign n43506 = ~n43502 & ~n43503;
  assign n43507 = ~n43504 & n43506;
  assign n43508 = ~n43505 & n43507;
  assign n43509 = P1_P1_INSTQUEUE_REG_7__3_ & n43375;
  assign n43510 = P1_P1_INSTQUEUE_REG_6__3_ & n43377;
  assign n43511 = P1_P1_INSTQUEUE_REG_5__3_ & n43379;
  assign n43512 = P1_P1_INSTQUEUE_REG_4__3_ & n43381;
  assign n43513 = ~n43509 & ~n43510;
  assign n43514 = ~n43511 & n43513;
  assign n43515 = ~n43512 & n43514;
  assign n43516 = P1_P1_INSTQUEUE_REG_3__3_ & n43386;
  assign n43517 = P1_P1_INSTQUEUE_REG_2__3_ & n43389;
  assign n43518 = P1_P1_INSTQUEUE_REG_1__3_ & n43391;
  assign n43519 = P1_P1_INSTQUEUE_REG_0__3_ & n43393;
  assign n43520 = ~n43516 & ~n43517;
  assign n43521 = ~n43518 & n43520;
  assign n43522 = ~n43519 & n43521;
  assign n43523 = n43498 & n43501;
  assign n43524 = n43508 & n43523;
  assign n43525 = n43515 & n43524;
  assign n43526 = n43522 & n43525;
  assign n43527 = P1_P1_INSTQUEUE_REG_11__2_ & n43346;
  assign n43528 = P1_P1_INSTQUEUE_REG_10__2_ & n43350;
  assign n43529 = ~n43527 & ~n43528;
  assign n43530 = P1_P1_INSTQUEUE_REG_9__2_ & n43355;
  assign n43531 = P1_P1_INSTQUEUE_REG_8__2_ & n43359;
  assign n43532 = ~n43530 & ~n43531;
  assign n43533 = P1_P1_INSTQUEUE_REG_15__2_ & n43363;
  assign n43534 = P1_P1_INSTQUEUE_REG_14__2_ & n43365;
  assign n43535 = P1_P1_INSTQUEUE_REG_13__2_ & n43367;
  assign n43536 = P1_P1_INSTQUEUE_REG_12__2_ & n43369;
  assign n43537 = ~n43533 & ~n43534;
  assign n43538 = ~n43535 & n43537;
  assign n43539 = ~n43536 & n43538;
  assign n43540 = P1_P1_INSTQUEUE_REG_7__2_ & n43375;
  assign n43541 = P1_P1_INSTQUEUE_REG_6__2_ & n43377;
  assign n43542 = P1_P1_INSTQUEUE_REG_5__2_ & n43379;
  assign n43543 = P1_P1_INSTQUEUE_REG_4__2_ & n43381;
  assign n43544 = ~n43540 & ~n43541;
  assign n43545 = ~n43542 & n43544;
  assign n43546 = ~n43543 & n43545;
  assign n43547 = P1_P1_INSTQUEUE_REG_3__2_ & n43386;
  assign n43548 = P1_P1_INSTQUEUE_REG_2__2_ & n43389;
  assign n43549 = P1_P1_INSTQUEUE_REG_1__2_ & n43391;
  assign n43550 = P1_P1_INSTQUEUE_REG_0__2_ & n43393;
  assign n43551 = ~n43547 & ~n43548;
  assign n43552 = ~n43549 & n43551;
  assign n43553 = ~n43550 & n43552;
  assign n43554 = n43529 & n43532;
  assign n43555 = n43539 & n43554;
  assign n43556 = n43546 & n43555;
  assign n43557 = n43553 & n43556;
  assign n43558 = ~n43495 & ~n43526;
  assign n43559 = n43557 & n43558;
  assign n43560 = n43433 & n43464;
  assign n43561 = n43559 & n43560;
  assign n43562 = P1_P1_INSTQUEUE_REG_11__1_ & n43346;
  assign n43563 = P1_P1_INSTQUEUE_REG_10__1_ & n43350;
  assign n43564 = ~n43562 & ~n43563;
  assign n43565 = P1_P1_INSTQUEUE_REG_9__1_ & n43355;
  assign n43566 = P1_P1_INSTQUEUE_REG_8__1_ & n43359;
  assign n43567 = ~n43565 & ~n43566;
  assign n43568 = P1_P1_INSTQUEUE_REG_15__1_ & n43363;
  assign n43569 = P1_P1_INSTQUEUE_REG_14__1_ & n43365;
  assign n43570 = P1_P1_INSTQUEUE_REG_13__1_ & n43367;
  assign n43571 = P1_P1_INSTQUEUE_REG_12__1_ & n43369;
  assign n43572 = ~n43568 & ~n43569;
  assign n43573 = ~n43570 & n43572;
  assign n43574 = ~n43571 & n43573;
  assign n43575 = P1_P1_INSTQUEUE_REG_7__1_ & n43375;
  assign n43576 = P1_P1_INSTQUEUE_REG_6__1_ & n43377;
  assign n43577 = P1_P1_INSTQUEUE_REG_5__1_ & n43379;
  assign n43578 = P1_P1_INSTQUEUE_REG_4__1_ & n43381;
  assign n43579 = ~n43575 & ~n43576;
  assign n43580 = ~n43577 & n43579;
  assign n43581 = ~n43578 & n43580;
  assign n43582 = P1_P1_INSTQUEUE_REG_3__1_ & n43386;
  assign n43583 = P1_P1_INSTQUEUE_REG_2__1_ & n43389;
  assign n43584 = P1_P1_INSTQUEUE_REG_1__1_ & n43391;
  assign n43585 = P1_P1_INSTQUEUE_REG_0__1_ & n43393;
  assign n43586 = ~n43582 & ~n43583;
  assign n43587 = ~n43584 & n43586;
  assign n43588 = ~n43585 & n43587;
  assign n43589 = n43564 & n43567;
  assign n43590 = n43574 & n43589;
  assign n43591 = n43581 & n43590;
  assign n43592 = n43588 & n43591;
  assign n43593 = P1_P1_INSTQUEUE_REG_11__0_ & n43346;
  assign n43594 = P1_P1_INSTQUEUE_REG_10__0_ & n43350;
  assign n43595 = ~n43593 & ~n43594;
  assign n43596 = P1_P1_INSTQUEUE_REG_9__0_ & n43355;
  assign n43597 = P1_P1_INSTQUEUE_REG_8__0_ & n43359;
  assign n43598 = ~n43596 & ~n43597;
  assign n43599 = P1_P1_INSTQUEUE_REG_15__0_ & n43363;
  assign n43600 = P1_P1_INSTQUEUE_REG_14__0_ & n43365;
  assign n43601 = P1_P1_INSTQUEUE_REG_13__0_ & n43367;
  assign n43602 = P1_P1_INSTQUEUE_REG_12__0_ & n43369;
  assign n43603 = ~n43599 & ~n43600;
  assign n43604 = ~n43601 & n43603;
  assign n43605 = ~n43602 & n43604;
  assign n43606 = P1_P1_INSTQUEUE_REG_7__0_ & n43375;
  assign n43607 = P1_P1_INSTQUEUE_REG_6__0_ & n43377;
  assign n43608 = P1_P1_INSTQUEUE_REG_5__0_ & n43379;
  assign n43609 = P1_P1_INSTQUEUE_REG_4__0_ & n43381;
  assign n43610 = ~n43606 & ~n43607;
  assign n43611 = ~n43608 & n43610;
  assign n43612 = ~n43609 & n43611;
  assign n43613 = P1_P1_INSTQUEUE_REG_3__0_ & n43386;
  assign n43614 = P1_P1_INSTQUEUE_REG_2__0_ & n43389;
  assign n43615 = P1_P1_INSTQUEUE_REG_1__0_ & n43391;
  assign n43616 = P1_P1_INSTQUEUE_REG_0__0_ & n43393;
  assign n43617 = ~n43613 & ~n43614;
  assign n43618 = ~n43615 & n43617;
  assign n43619 = ~n43616 & n43618;
  assign n43620 = n43595 & n43598;
  assign n43621 = n43605 & n43620;
  assign n43622 = n43612 & n43621;
  assign n43623 = n43619 & n43622;
  assign n43624 = n43592 & ~n43623;
  assign n43625 = n43561 & n43624;
  assign n43626 = n43343 & n43625;
  assign n43627 = ~P1_P1_STATE2_REG_1_ & ~n43626;
  assign n43628 = ~n43251 & n43342;
  assign n43629 = ~n43557 & ~n43592;
  assign n43630 = n43628 & n43629;
  assign n43631 = ~n43251 & ~n43557;
  assign n43632 = n43592 & n43631;
  assign n43633 = ~n43251 & n43557;
  assign n43634 = n43592 & ~n43628;
  assign n43635 = n43633 & ~n43634;
  assign n43636 = ~n43630 & ~n43632;
  assign n43637 = ~n43635 & n43636;
  assign n43638 = P1_P1_INSTQUEUERD_ADDR_REG_4_ & ~P1_P1_INSTQUEUEWR_ADDR_REG_4_;
  assign n43639 = ~P1_P1_INSTQUEUERD_ADDR_REG_3_ & P1_P1_INSTQUEUEWR_ADDR_REG_3_;
  assign n43640 = P1_P1_INSTQUEUERD_ADDR_REG_3_ & ~P1_P1_INSTQUEUEWR_ADDR_REG_3_;
  assign n43641 = ~P1_P1_INSTQUEUERD_ADDR_REG_2_ & P1_P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n43642 = P1_P1_INSTQUEUERD_ADDR_REG_2_ & ~P1_P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n43643 = P1_P1_INSTQUEUERD_ADDR_REG_0_ & ~P1_P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n43644 = P1_P1_INSTQUEUEWR_ADDR_REG_1_ & ~n43643;
  assign n43645 = ~P1_P1_INSTQUEUEWR_ADDR_REG_1_ & n43643;
  assign n43646 = ~P1_P1_INSTQUEUERD_ADDR_REG_1_ & ~n43645;
  assign n43647 = ~n43644 & ~n43646;
  assign n43648 = ~n43642 & ~n43647;
  assign n43649 = ~n43641 & ~n43648;
  assign n43650 = ~n43640 & ~n43649;
  assign n43651 = ~n43639 & ~n43650;
  assign n43652 = ~P1_P1_INSTQUEUERD_ADDR_REG_4_ & P1_P1_INSTQUEUEWR_ADDR_REG_4_;
  assign n43653 = n43651 & ~n43652;
  assign n43654 = ~n43638 & ~n43653;
  assign n43655 = ~n43638 & ~n43652;
  assign n43656 = ~n43651 & ~n43655;
  assign n43657 = n43651 & n43655;
  assign n43658 = ~n43656 & ~n43657;
  assign n43659 = ~n43639 & ~n43640;
  assign n43660 = ~n43649 & ~n43659;
  assign n43661 = n43649 & n43659;
  assign n43662 = ~n43660 & ~n43661;
  assign n43663 = ~P1_P1_INSTQUEUERD_ADDR_REG_1_ & P1_P1_INSTQUEUEWR_ADDR_REG_1_;
  assign n43664 = P1_P1_INSTQUEUERD_ADDR_REG_1_ & ~P1_P1_INSTQUEUEWR_ADDR_REG_1_;
  assign n43665 = ~n43663 & ~n43664;
  assign n43666 = ~n43643 & ~n43665;
  assign n43667 = n43643 & n43665;
  assign n43668 = ~n43666 & ~n43667;
  assign n43669 = ~n43641 & ~n43642;
  assign n43670 = ~n43647 & ~n43669;
  assign n43671 = n43647 & n43669;
  assign n43672 = ~n43670 & ~n43671;
  assign n43673 = n43658 & n43662;
  assign n43674 = n43668 & n43673;
  assign n43675 = n43672 & n43674;
  assign n43676 = n43654 & ~n43675;
  assign n43677 = ~n43592 & ~n43676;
  assign n43678 = n43592 & ~n43676;
  assign n43679 = ~n43677 & ~n43678;
  assign n43680 = ~n43495 & n43526;
  assign n43681 = ~n43401 & ~n43432;
  assign n43682 = n43464 & n43681;
  assign n43683 = n43680 & n43682;
  assign n43684 = n43623 & n43683;
  assign n43685 = n43679 & n43684;
  assign n43686 = ~n43557 & ~n43685;
  assign n43687 = ~n43526 & ~n43623;
  assign n43688 = ~n43495 & n43687;
  assign n43689 = n43560 & n43688;
  assign n43690 = ~n43677 & n43689;
  assign n43691 = ~n43678 & n43690;
  assign n43692 = n43557 & ~n43691;
  assign n43693 = ~n43686 & ~n43692;
  assign n43694 = n43637 & n43693;
  assign n43695 = ~P1_P1_FLUSH_REG & ~P1_P1_MORE_REG;
  assign n43696 = n43694 & ~n43695;
  assign n43697 = ~n43592 & n43623;
  assign n43698 = ~n43557 & n43697;
  assign n43699 = n43683 & n43698;
  assign n43700 = ~n43676 & n43699;
  assign n43701 = n43592 & n43623;
  assign n43702 = ~n43557 & n43701;
  assign n43703 = n43683 & n43702;
  assign n43704 = ~n43676 & n43703;
  assign n43705 = n43625 & ~n43676;
  assign n43706 = ~n43592 & ~n43623;
  assign n43707 = n43561 & n43706;
  assign n43708 = ~n43676 & n43707;
  assign n43709 = ~n43700 & ~n43704;
  assign n43710 = ~n43705 & n43709;
  assign n43711 = ~n43708 & n43710;
  assign n43712 = ~n43401 & n43432;
  assign n43713 = ~n43464 & n43712;
  assign n43714 = n43559 & n43713;
  assign n43715 = n43706 & n43714;
  assign n43716 = ~P1_P1_INSTQUEUERD_ADDR_REG_0_ & P1_P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n43717 = ~n43643 & ~n43716;
  assign n43718 = n43668 & n43717;
  assign n43719 = ~n43672 & ~n43718;
  assign n43720 = n43673 & ~n43719;
  assign n43721 = n43654 & ~n43720;
  assign n43722 = n43715 & ~n43721;
  assign n43723 = n43701 & n43714;
  assign n43724 = ~n43721 & n43723;
  assign n43725 = n43559 & n43682;
  assign n43726 = n43624 & n43725;
  assign n43727 = n43658 & ~n43719;
  assign n43728 = n43662 & n43727;
  assign n43729 = n43654 & ~n43728;
  assign n43730 = n43726 & ~n43729;
  assign n43731 = n43706 & n43725;
  assign n43732 = ~n43668 & ~n43717;
  assign n43733 = n43673 & ~n43732;
  assign n43734 = n43672 & n43733;
  assign n43735 = n43654 & ~n43734;
  assign n43736 = n43731 & ~n43735;
  assign n43737 = ~n43722 & ~n43724;
  assign n43738 = ~n43730 & n43737;
  assign n43739 = ~n43736 & n43738;
  assign n43740 = n43711 & n43739;
  assign n43741 = ~n43694 & ~n43740;
  assign n43742 = ~n43592 & ~n43735;
  assign n43743 = n43592 & ~n43729;
  assign n43744 = ~n43742 & ~n43743;
  assign n43745 = ~n43623 & n43725;
  assign n43746 = n43744 & n43745;
  assign n43747 = n43526 & n43557;
  assign n43748 = n43401 & ~n43432;
  assign n43749 = n43747 & n43748;
  assign n43750 = n43701 & n43749;
  assign n43751 = ~n43495 & n43750;
  assign n43752 = n43561 & ~n43623;
  assign n43753 = ~n43699 & ~n43751;
  assign n43754 = ~n43752 & n43753;
  assign n43755 = n43432 & n43526;
  assign n43756 = ~n43464 & n43557;
  assign n43757 = ~n43495 & n43701;
  assign n43758 = n43756 & n43757;
  assign n43759 = n43401 & ~n43557;
  assign n43760 = n43464 & n43495;
  assign n43761 = n43759 & n43760;
  assign n43762 = ~n43758 & ~n43761;
  assign n43763 = n43755 & ~n43762;
  assign n43764 = n43706 & n43760;
  assign n43765 = n43749 & n43764;
  assign n43766 = n43526 & ~n43557;
  assign n43767 = n43495 & n43697;
  assign n43768 = n43682 & n43766;
  assign n43769 = n43767 & n43768;
  assign n43770 = ~n43592 & n43725;
  assign n43771 = ~n43769 & ~n43770;
  assign n43772 = ~n43763 & ~n43765;
  assign n43773 = n43771 & n43772;
  assign n43774 = n43432 & ~n43495;
  assign n43775 = ~n43748 & ~n43774;
  assign n43776 = n43526 & n43775;
  assign n43777 = ~n43557 & ~n43776;
  assign n43778 = ~n43495 & ~n43748;
  assign n43779 = ~n43712 & n43778;
  assign n43780 = ~n43526 & n43779;
  assign n43781 = n43624 & ~n43780;
  assign n43782 = n43681 & n43701;
  assign n43783 = n43401 & n43495;
  assign n43784 = ~n43558 & ~n43783;
  assign n43785 = ~n43592 & n43784;
  assign n43786 = n43432 & n43464;
  assign n43787 = n43623 & n43786;
  assign n43788 = ~n43782 & ~n43785;
  assign n43789 = ~n43787 & n43788;
  assign n43790 = ~n43781 & n43789;
  assign n43791 = n43557 & ~n43790;
  assign n43792 = ~n43526 & ~n43786;
  assign n43793 = n43401 & n43792;
  assign n43794 = n43495 & n43592;
  assign n43795 = n43623 & ~n43794;
  assign n43796 = n43526 & ~n43795;
  assign n43797 = ~n43401 & n43796;
  assign n43798 = ~n43495 & ~n43681;
  assign n43799 = ~n43624 & n43798;
  assign n43800 = ~n43464 & ~n43799;
  assign n43801 = n43432 & ~n43592;
  assign n43802 = n43495 & n43801;
  assign n43803 = n43464 & ~n43592;
  assign n43804 = n43712 & n43803;
  assign n43805 = ~n43681 & n43697;
  assign n43806 = ~n43802 & ~n43804;
  assign n43807 = ~n43805 & n43806;
  assign n43808 = ~n43793 & ~n43797;
  assign n43809 = ~n43800 & n43808;
  assign n43810 = n43807 & n43809;
  assign n43811 = ~n43777 & ~n43791;
  assign n43812 = n43810 & n43811;
  assign n43813 = n43773 & n43812;
  assign n43814 = ~n43750 & n43813;
  assign n43815 = P1_P1_INSTQUEUERD_ADDR_REG_0_ & ~n43814;
  assign n43816 = n43754 & ~n43815;
  assign n43817 = ~P1_P1_INSTQUEUERD_ADDR_REG_2_ & ~n43816;
  assign n43818 = P1_P1_INSTQUEUERD_ADDR_REG_1_ & n43817;
  assign n43819 = P1_P1_INSTQUEUERD_ADDR_REG_2_ & ~n43754;
  assign n43820 = ~P1_P1_INSTQUEUERD_ADDR_REG_1_ & n43819;
  assign n43821 = ~P1_P1_INSTQUEUERD_ADDR_REG_2_ & P1_P1_INSTQUEUERD_ADDR_REG_1_;
  assign n43822 = P1_P1_INSTQUEUERD_ADDR_REG_2_ & ~P1_P1_INSTQUEUERD_ADDR_REG_1_;
  assign n43823 = ~n43821 & ~n43822;
  assign n43824 = n43703 & ~n43823;
  assign n43825 = P1_P1_INSTQUEUERD_ADDR_REG_2_ & ~n43344;
  assign n43826 = ~n43345 & ~n43825;
  assign n43827 = ~n43701 & ~n43706;
  assign n43828 = n43826 & ~n43827;
  assign n43829 = n43714 & n43828;
  assign n43830 = ~n43824 & ~n43829;
  assign n43831 = n43592 & n43755;
  assign n43832 = ~n43756 & ~n43761;
  assign n43833 = n43831 & ~n43832;
  assign n43834 = n43760 & ~n43827;
  assign n43835 = n43749 & n43834;
  assign n43836 = ~n43833 & ~n43835;
  assign n43837 = n43771 & n43836;
  assign n43838 = n43812 & n43837;
  assign n43839 = n43825 & ~n43838;
  assign n43840 = n43830 & ~n43839;
  assign n43841 = ~n43818 & ~n43820;
  assign n43842 = n43840 & n43841;
  assign n43843 = n43464 & n43623;
  assign n43844 = ~n43526 & ~n43697;
  assign n43845 = n43778 & ~n43843;
  assign n43846 = n43844 & n43845;
  assign n43847 = ~n43804 & n43846;
  assign n43848 = n43557 & ~n43847;
  assign n43849 = ~n43557 & ~n43684;
  assign n43850 = n43624 & ~n43779;
  assign n43851 = ~n43848 & ~n43849;
  assign n43852 = ~n43850 & n43851;
  assign n43853 = n43721 & n43723;
  assign n43854 = n43676 & n43703;
  assign n43855 = n43676 & n43707;
  assign n43856 = ~n43854 & ~n43855;
  assign n43857 = ~n43251 & ~n43856;
  assign n43858 = ~n43853 & ~n43857;
  assign n43859 = n43715 & n43721;
  assign n43860 = ~n43712 & n43756;
  assign n43861 = ~n43859 & ~n43860;
  assign n43862 = n43676 & n43699;
  assign n43863 = n43625 & n43676;
  assign n43864 = ~n43862 & ~n43863;
  assign n43865 = n43628 & ~n43864;
  assign n43866 = n43861 & ~n43865;
  assign n43867 = n43852 & n43858;
  assign n43868 = n43866 & n43867;
  assign n43869 = ~n43842 & ~n43868;
  assign n43870 = P1_P1_INSTQUEUERD_ADDR_REG_2_ & n43868;
  assign n43871 = ~n43869 & ~n43870;
  assign n43872 = P1_P1_INSTQUEUERD_ADDR_REG_1_ & n43374;
  assign n43873 = ~n43816 & n43872;
  assign n43874 = P1_P1_INSTQUEUERD_ADDR_REG_2_ & n43344;
  assign n43875 = P1_P1_INSTQUEUERD_ADDR_REG_3_ & ~n43874;
  assign n43876 = ~n43837 & n43875;
  assign n43877 = P1_P1_INSTQUEUERD_ADDR_REG_2_ & P1_P1_INSTQUEUERD_ADDR_REG_1_;
  assign n43878 = ~P1_P1_INSTQUEUERD_ADDR_REG_3_ & n43877;
  assign n43879 = P1_P1_INSTQUEUERD_ADDR_REG_3_ & ~n43877;
  assign n43880 = ~n43878 & ~n43879;
  assign n43881 = n43703 & ~n43880;
  assign n43882 = ~n43876 & ~n43881;
  assign n43883 = ~n43464 & n43751;
  assign n43884 = n43464 & n43751;
  assign n43885 = ~n43625 & ~n43707;
  assign n43886 = ~n43699 & n43885;
  assign n43887 = ~n43883 & ~n43884;
  assign n43888 = n43886 & n43887;
  assign n43889 = n43812 & n43888;
  assign n43890 = n43879 & ~n43889;
  assign n43891 = P1_P1_INSTQUEUERD_ADDR_REG_3_ & ~P1_P1_INSTQUEUERD_ADDR_REG_0_;
  assign n43892 = ~n43812 & n43891;
  assign n43893 = ~n43344 & n43388;
  assign n43894 = ~P1_P1_INSTQUEUERD_ADDR_REG_2_ & ~n43344;
  assign n43895 = P1_P1_INSTQUEUERD_ADDR_REG_3_ & ~n43894;
  assign n43896 = ~n43893 & ~n43895;
  assign n43897 = ~n43827 & n43896;
  assign n43898 = n43714 & n43897;
  assign n43899 = ~n43892 & ~n43898;
  assign n43900 = n43882 & ~n43890;
  assign n43901 = n43899 & n43900;
  assign n43902 = ~n43873 & n43901;
  assign n43903 = ~n43868 & ~n43902;
  assign n43904 = P1_P1_INSTQUEUERD_ADDR_REG_3_ & n43868;
  assign n43905 = ~n43903 & ~n43904;
  assign n43906 = ~n43871 & ~n43905;
  assign n43907 = P1_P1_INSTQUEUERD_ADDR_REG_4_ & n43868;
  assign n43908 = P1_P1_INSTQUEUERD_ADDR_REG_3_ & n43877;
  assign n43909 = ~P1_P1_INSTQUEUERD_ADDR_REG_4_ & n43908;
  assign n43910 = P1_P1_INSTQUEUERD_ADDR_REG_4_ & ~n43908;
  assign n43911 = ~n43909 & ~n43910;
  assign n43912 = n43703 & ~n43911;
  assign n43913 = ~n43868 & n43912;
  assign n43914 = ~n43907 & ~n43913;
  assign n43915 = ~n43906 & n43914;
  assign n43916 = ~P1_P1_INSTQUEUEWR_ADDR_REG_3_ & ~n43905;
  assign n43917 = ~P1_P1_INSTQUEUEWR_ADDR_REG_4_ & ~n43914;
  assign n43918 = ~n43916 & ~n43917;
  assign n43919 = P1_P1_INSTQUEUEWR_ADDR_REG_2_ & n43871;
  assign n43920 = P1_P1_INSTQUEUEWR_ADDR_REG_3_ & n43905;
  assign n43921 = ~n43919 & ~n43920;
  assign n43922 = ~P1_P1_INSTQUEUEWR_ADDR_REG_2_ & ~n43871;
  assign n43923 = n43712 & n43758;
  assign n43924 = ~n43715 & ~n43923;
  assign n43925 = n43750 & n43760;
  assign n43926 = n43813 & ~n43925;
  assign n43927 = n43924 & n43926;
  assign n43928 = ~P1_P1_INSTQUEUERD_ADDR_REG_0_ & ~n43927;
  assign n43929 = P1_P1_INSTQUEUERD_ADDR_REG_0_ & ~n43754;
  assign n43930 = P1_P1_INSTQUEUERD_ADDR_REG_0_ & n43703;
  assign n43931 = ~n43928 & ~n43929;
  assign n43932 = ~n43930 & n43931;
  assign n43933 = ~n43868 & ~n43932;
  assign n43934 = P1_P1_INSTQUEUERD_ADDR_REG_0_ & n43868;
  assign n43935 = ~n43933 & ~n43934;
  assign n43936 = P1_P1_INSTQUEUEWR_ADDR_REG_0_ & n43935;
  assign n43937 = ~P1_P1_INSTQUEUEWR_ADDR_REG_1_ & ~n43936;
  assign n43938 = ~P1_P1_INSTQUEUERD_ADDR_REG_1_ & ~n43816;
  assign n43939 = ~P1_P1_INSTQUEUERD_ADDR_REG_1_ & n43703;
  assign n43940 = ~n43344 & ~n43357;
  assign n43941 = ~n43924 & n43940;
  assign n43942 = ~n43939 & ~n43941;
  assign n43943 = n43348 & ~n43926;
  assign n43944 = n43942 & ~n43943;
  assign n43945 = ~n43938 & n43944;
  assign n43946 = ~n43868 & ~n43945;
  assign n43947 = P1_P1_INSTQUEUERD_ADDR_REG_1_ & n43868;
  assign n43948 = ~n43946 & ~n43947;
  assign n43949 = ~P1_P1_INSTQUEUEWR_ADDR_REG_1_ & ~n43948;
  assign n43950 = ~n43936 & ~n43948;
  assign n43951 = ~n43922 & ~n43937;
  assign n43952 = ~n43949 & n43951;
  assign n43953 = ~n43950 & n43952;
  assign n43954 = n43921 & ~n43953;
  assign n43955 = n43918 & ~n43954;
  assign n43956 = P1_P1_INSTQUEUEWR_ADDR_REG_4_ & n43914;
  assign n43957 = ~n43955 & ~n43956;
  assign n43958 = ~n43696 & ~n43741;
  assign n43959 = ~n43746 & n43958;
  assign n43960 = n43915 & n43959;
  assign n43961 = ~n43957 & n43960;
  assign n43962 = n43627 & n43961;
  assign n43963 = P1_P1_STATE2_REG_0_ & ~n43962;
  assign n43964 = ~n43338 & ~n43963;
  assign n43965 = P1_P1_STATE2_REG_2_ & n43964;
  assign n43966 = P1_P1_STATE2_REG_0_ & ~n43965;
  assign n43967 = n43336 & n43966;
  assign n43968 = P1_P1_STATE2_REG_3_ & ~n43966;
  assign n8086 = n43967 | n43968;
  assign n43970 = ~P1_P1_STATE2_REG_2_ & ~n43251;
  assign n43971 = P1_P1_STATE2_REG_0_ & ~n43970;
  assign n43972 = ~P1_P1_STATE2_REG_0_ & ~P1_P1_STATEBS16_REG;
  assign n43973 = ~n43971 & ~n43972;
  assign n43974 = P1_P1_STATE2_REG_1_ & n43973;
  assign n43975 = P1_P1_STATE2_REG_2_ & ~P1_P1_STATE2_REG_1_;
  assign n43976 = ~n43974 & ~n43975;
  assign n43977 = P1_P1_STATE2_REG_2_ & ~n43966;
  assign n8091 = ~n43976 | n43977;
  assign n43979 = P1_P1_STATE2_REG_0_ & n43975;
  assign n43980 = ~n43965 & n43979;
  assign n43981 = ~P1_P1_STATE2_REG_2_ & P1_P1_STATE2_REG_0_;
  assign n43982 = n43251 & n43981;
  assign n43983 = ~n43965 & ~n43982;
  assign n43984 = P1_P1_STATE2_REG_1_ & ~n43983;
  assign n43985 = ~P1_P1_STATE2_REG_3_ & ~P1_P1_STATE2_REG_1_;
  assign n43986 = ~n43251 & n43985;
  assign n43987 = n43966 & n43986;
  assign n43988 = P1_P1_STATE2_REG_1_ & ~P1_P1_STATE2_REG_0_;
  assign n43989 = ~P1_P1_STATE2_REG_2_ & n43988;
  assign n43990 = ~P1_P1_STATEBS16_REG & n43989;
  assign n43991 = ~n43980 & ~n43984;
  assign n43992 = ~n43987 & n43991;
  assign n8096 = n43990 | ~n43992;
  assign n43994 = P1_P1_STATE2_REG_3_ & ~P1_P1_INSTQUEUERD_ADDR_REG_4_;
  assign n43995 = ~P1_P1_STATE2_REG_2_ & ~P1_P1_STATE2_REG_1_;
  assign n43996 = n43994 & n43995;
  assign n43997 = ~n43965 & ~n43996;
  assign n43998 = ~P1_P1_STATE2_REG_0_ & n43997;
  assign n43999 = P1_P1_INSTADDRPOINTER_REG_0_ & P1_P1_INSTADDRPOINTER_REG_31_;
  assign n44000 = P1_P1_INSTADDRPOINTER_REG_0_ & ~P1_P1_INSTADDRPOINTER_REG_31_;
  assign n44001 = ~n43999 & ~n44000;
  assign n44002 = P1_P1_FLUSH_REG & n44001;
  assign n44003 = P1_P1_INSTQUEUERD_ADDR_REG_0_ & ~P1_P1_FLUSH_REG;
  assign n44004 = ~n44002 & ~n44003;
  assign n44005 = P1_P1_INSTADDRPOINTER_REG_0_ & ~P1_P1_INSTADDRPOINTER_REG_1_;
  assign n44006 = ~P1_P1_INSTADDRPOINTER_REG_0_ & P1_P1_INSTADDRPOINTER_REG_1_;
  assign n44007 = ~n44005 & ~n44006;
  assign n44008 = P1_P1_INSTADDRPOINTER_REG_31_ & ~n44007;
  assign n44009 = P1_P1_INSTADDRPOINTER_REG_1_ & ~P1_P1_INSTADDRPOINTER_REG_31_;
  assign n44010 = ~n44008 & ~n44009;
  assign n44011 = ~n44001 & n44010;
  assign n44012 = P1_P1_FLUSH_REG & n44011;
  assign n44013 = P1_P1_INSTQUEUERD_ADDR_REG_1_ & ~P1_P1_FLUSH_REG;
  assign n44014 = ~n44012 & ~n44013;
  assign n44015 = n44004 & n44014;
  assign n44016 = P1_P1_INSTQUEUERD_ADDR_REG_3_ & ~P1_P1_FLUSH_REG;
  assign n44017 = ~n44001 & ~n44010;
  assign n44018 = P1_P1_FLUSH_REG & n44017;
  assign n44019 = P1_P1_INSTQUEUERD_ADDR_REG_2_ & ~P1_P1_FLUSH_REG;
  assign n44020 = ~n44018 & ~n44019;
  assign n44021 = ~n44015 & n44016;
  assign n44022 = ~n44020 & n44021;
  assign n44023 = P1_P1_INSTQUEUERD_ADDR_REG_4_ & ~P1_P1_FLUSH_REG;
  assign n44024 = ~n44022 & ~n44023;
  assign n44025 = n43336 & n44024;
  assign n44026 = ~n43965 & ~n44025;
  assign n44027 = P1_P1_STATE2_REG_0_ & ~n44026;
  assign n44028 = P1_P1_STATE2_REG_3_ & P1_P1_STATE2_REG_0_;
  assign n44029 = n43995 & n44028;
  assign n44030 = ~n43982 & ~n44029;
  assign n44031 = ~n43961 & n43979;
  assign n44032 = n44030 & ~n44031;
  assign n44033 = ~n43998 & ~n44027;
  assign n8101 = ~n44032 | ~n44033;
  assign n44035 = P1_P1_INSTQUEUEWR_ADDR_REG_1_ & P1_P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n44036 = P1_P1_INSTQUEUEWR_ADDR_REG_2_ & n44035;
  assign n44037 = P1_P1_INSTQUEUEWR_ADDR_REG_3_ & n44036;
  assign n44038 = P1_P1_STATE2_REG_3_ & ~n44037;
  assign n44039 = ~P1_P1_STATE2_REG_2_ & P1_P1_STATE2_REG_1_;
  assign n44040 = ~n43975 & ~n44039;
  assign n44041 = ~n43994 & n44040;
  assign n44042 = ~P1_P1_STATE2_REG_0_ & ~n44041;
  assign n44043 = ~n44038 & n44042;
  assign n44044 = ~P1_P1_INSTQUEUEWR_ADDR_REG_2_ & n44035;
  assign n44045 = P1_P1_INSTQUEUEWR_ADDR_REG_2_ & ~n44035;
  assign n44046 = ~n44044 & ~n44045;
  assign n44047 = ~P1_P1_INSTQUEUEWR_ADDR_REG_3_ & n44036;
  assign n44048 = P1_P1_INSTQUEUEWR_ADDR_REG_3_ & ~n44036;
  assign n44049 = ~n44047 & ~n44048;
  assign n44050 = ~n44046 & ~n44049;
  assign n44051 = ~P1_P1_INSTQUEUEWR_ADDR_REG_1_ & P1_P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n44052 = P1_P1_INSTQUEUEWR_ADDR_REG_1_ & ~P1_P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n44053 = ~n44051 & ~n44052;
  assign n44054 = ~P1_P1_INSTQUEUEWR_ADDR_REG_0_ & ~n44053;
  assign n44055 = n44050 & n44054;
  assign n44056 = ~n44037 & ~n44055;
  assign n44057 = ~P1_P1_STATE2_REG_3_ & ~P1_P1_STATE2_REG_2_;
  assign n44058 = ~P1_P1_STATEBS16_REG & n44057;
  assign n44059 = ~P1_P1_STATE2_REG_2_ & ~n44058;
  assign n44060 = P1_P1_INSTQUEUEWR_ADDR_REG_0_ & ~n44053;
  assign n44061 = ~P1_P1_INSTQUEUEWR_ADDR_REG_0_ & n44053;
  assign n44062 = ~n44060 & ~n44061;
  assign n44063 = ~P1_P1_INSTQUEUEWR_ADDR_REG_0_ & ~n44062;
  assign n44064 = P1_P1_INSTQUEUEWR_ADDR_REG_0_ & n44062;
  assign n44065 = ~n44063 & ~n44064;
  assign n44066 = ~P1_P1_INSTQUEUEWR_ADDR_REG_0_ & ~n44065;
  assign n44067 = ~n44046 & ~n44054;
  assign n44068 = n44046 & n44054;
  assign n44069 = ~n44067 & ~n44068;
  assign n44070 = P1_P1_INSTQUEUEWR_ADDR_REG_0_ & ~n44062;
  assign n44071 = ~n44069 & ~n44070;
  assign n44072 = n44069 & n44070;
  assign n44073 = ~n44071 & ~n44072;
  assign n44074 = ~n44046 & n44049;
  assign n44075 = n44054 & n44074;
  assign n44076 = ~n44046 & n44054;
  assign n44077 = ~n44049 & ~n44076;
  assign n44078 = ~n44075 & ~n44077;
  assign n44079 = n44069 & ~n44078;
  assign n44080 = ~n44070 & ~n44078;
  assign n44081 = ~n44079 & ~n44080;
  assign n44082 = ~n44069 & n44078;
  assign n44083 = n44070 & n44082;
  assign n44084 = n44081 & ~n44083;
  assign n44085 = ~n44073 & ~n44084;
  assign n44086 = n44066 & n44085;
  assign n44087 = ~n44069 & ~n44078;
  assign n44088 = n44070 & n44087;
  assign n44089 = ~n44086 & ~n44088;
  assign n44090 = n44059 & ~n44089;
  assign n44091 = n44056 & ~n44090;
  assign n44092 = n44043 & ~n44091;
  assign n44093 = P1_P1_INSTQUEUE_REG_15__7_ & ~n44092;
  assign n44094 = P1_P1_STATE2_REG_3_ & n44042;
  assign n44095 = ~n43495 & n44094;
  assign n44096 = n44037 & n44095;
  assign n44097 = P1_P1_STATEBS16_REG & n44057;
  assign n44098 = n44089 & n44097;
  assign n44099 = n44059 & ~n44098;
  assign n44100 = ~n44056 & ~n44099;
  assign n44101 = P1_BUF1_REG_7_ & n12460;
  assign n44102 = SEL & DIN_6_;
  assign n44103 = P4_DATAO_REG_0_ & n44102;
  assign n44104 = SEL & DIN_5_;
  assign n44105 = P4_DATAO_REG_0_ & n44104;
  assign n44106 = SEL & DIN_3_;
  assign n44107 = P4_DATAO_REG_1_ & n44106;
  assign n44108 = SEL & DIN_2_;
  assign n44109 = P4_DATAO_REG_1_ & n44108;
  assign n44110 = SEL & DIN_1_;
  assign n44111 = P4_DATAO_REG_2_ & n44110;
  assign n44112 = SEL & DIN_0_;
  assign n44113 = P4_DATAO_REG_3_ & n44112;
  assign n44114 = n44111 & ~n44113;
  assign n44115 = ~n44111 & n44113;
  assign n44116 = ~n44114 & ~n44115;
  assign n44117 = n44109 & ~n44116;
  assign n44118 = P4_DATAO_REG_1_ & P4_DATAO_REG_2_;
  assign n44119 = n44110 & n44112;
  assign n44120 = n44118 & n44119;
  assign n44121 = ~n44109 & n44116;
  assign n44122 = n44120 & ~n44121;
  assign n44123 = ~n44117 & ~n44122;
  assign n44124 = n44107 & ~n44123;
  assign n44125 = P4_DATAO_REG_2_ & n44108;
  assign n44126 = P4_DATAO_REG_4_ & n44112;
  assign n44127 = P4_DATAO_REG_3_ & n44110;
  assign n44128 = n44126 & ~n44127;
  assign n44129 = ~n44126 & n44127;
  assign n44130 = ~n44128 & ~n44129;
  assign n44131 = n44125 & ~n44130;
  assign n44132 = ~n44125 & n44130;
  assign n44133 = P4_DATAO_REG_2_ & P4_DATAO_REG_3_;
  assign n44134 = n44119 & n44133;
  assign n44135 = ~n44131 & ~n44132;
  assign n44136 = ~n44134 & n44135;
  assign n44137 = n44134 & ~n44135;
  assign n44138 = ~n44136 & ~n44137;
  assign n44139 = n44107 & ~n44138;
  assign n44140 = ~n44123 & ~n44138;
  assign n44141 = ~n44124 & ~n44139;
  assign n44142 = ~n44140 & n44141;
  assign n44143 = SEL & DIN_4_;
  assign n44144 = P4_DATAO_REG_1_ & n44143;
  assign n44145 = ~n44132 & n44134;
  assign n44146 = ~n44131 & ~n44145;
  assign n44147 = P4_DATAO_REG_2_ & n44106;
  assign n44148 = P4_DATAO_REG_3_ & n44108;
  assign n44149 = P4_DATAO_REG_5_ & n44112;
  assign n44150 = P4_DATAO_REG_4_ & n44110;
  assign n44151 = n44149 & ~n44150;
  assign n44152 = ~n44149 & n44150;
  assign n44153 = ~n44151 & ~n44152;
  assign n44154 = n44148 & ~n44153;
  assign n44155 = ~n44148 & n44153;
  assign n44156 = P4_DATAO_REG_3_ & P4_DATAO_REG_4_;
  assign n44157 = n44119 & n44156;
  assign n44158 = ~n44154 & ~n44155;
  assign n44159 = ~n44157 & n44158;
  assign n44160 = n44155 & n44157;
  assign n44161 = n44148 & n44157;
  assign n44162 = ~n44153 & n44161;
  assign n44163 = ~n44159 & ~n44160;
  assign n44164 = ~n44162 & n44163;
  assign n44165 = n44147 & ~n44164;
  assign n44166 = ~n44147 & n44164;
  assign n44167 = ~n44165 & ~n44166;
  assign n44168 = n44146 & ~n44167;
  assign n44169 = ~n44147 & ~n44164;
  assign n44170 = ~n44146 & n44169;
  assign n44171 = ~n44146 & n44147;
  assign n44172 = n44164 & n44171;
  assign n44173 = ~n44168 & ~n44170;
  assign n44174 = ~n44172 & n44173;
  assign n44175 = n44144 & ~n44174;
  assign n44176 = ~n44144 & n44174;
  assign n44177 = ~n44175 & ~n44176;
  assign n44178 = n44142 & ~n44177;
  assign n44179 = n44144 & n44174;
  assign n44180 = ~n44144 & ~n44174;
  assign n44181 = ~n44179 & ~n44180;
  assign n44182 = ~n44142 & ~n44181;
  assign n44183 = ~n44178 & ~n44182;
  assign n44184 = n44105 & ~n44183;
  assign n44185 = ~n44105 & n44183;
  assign n44186 = P4_DATAO_REG_0_ & n44143;
  assign n44187 = P4_DATAO_REG_0_ & n44106;
  assign n44188 = ~n44117 & ~n44121;
  assign n44189 = ~n44120 & n44188;
  assign n44190 = n44120 & ~n44188;
  assign n44191 = ~n44189 & ~n44190;
  assign n44192 = n44187 & ~n44191;
  assign n44193 = ~n44187 & n44191;
  assign n44194 = P4_DATAO_REG_1_ & n44110;
  assign n44195 = P4_DATAO_REG_0_ & n44112;
  assign n44196 = n44194 & n44195;
  assign n44197 = P4_DATAO_REG_0_ & n44108;
  assign n44198 = n44196 & n44197;
  assign n44199 = ~n44196 & ~n44197;
  assign n44200 = P4_DATAO_REG_2_ & n44112;
  assign n44201 = n44194 & ~n44200;
  assign n44202 = ~n44194 & n44200;
  assign n44203 = ~n44201 & ~n44202;
  assign n44204 = ~n44199 & ~n44203;
  assign n44205 = ~n44198 & ~n44204;
  assign n44206 = ~n44193 & ~n44205;
  assign n44207 = ~n44192 & ~n44206;
  assign n44208 = n44186 & ~n44207;
  assign n44209 = ~n44107 & n44138;
  assign n44210 = ~n44139 & ~n44209;
  assign n44211 = n44123 & ~n44210;
  assign n44212 = ~n44107 & ~n44138;
  assign n44213 = ~n44123 & n44212;
  assign n44214 = n44124 & n44138;
  assign n44215 = ~n44211 & ~n44213;
  assign n44216 = ~n44214 & n44215;
  assign n44217 = ~n44186 & n44207;
  assign n44218 = n44216 & ~n44217;
  assign n44219 = ~n44208 & ~n44218;
  assign n44220 = ~n44185 & ~n44219;
  assign n44221 = ~n44184 & ~n44220;
  assign n44222 = n44103 & ~n44221;
  assign n44223 = ~n44142 & ~n44180;
  assign n44224 = ~n44179 & ~n44223;
  assign n44225 = P4_DATAO_REG_1_ & n44104;
  assign n44226 = P4_DATAO_REG_2_ & n44143;
  assign n44227 = ~n44148 & ~n44157;
  assign n44228 = ~n44153 & ~n44227;
  assign n44229 = ~n44161 & ~n44228;
  assign n44230 = P4_DATAO_REG_3_ & n44106;
  assign n44231 = P4_DATAO_REG_4_ & n44108;
  assign n44232 = P4_DATAO_REG_6_ & n44112;
  assign n44233 = P4_DATAO_REG_5_ & n44110;
  assign n44234 = n44232 & ~n44233;
  assign n44235 = ~n44232 & n44233;
  assign n44236 = ~n44234 & ~n44235;
  assign n44237 = n44231 & ~n44236;
  assign n44238 = ~n44231 & n44236;
  assign n44239 = P4_DATAO_REG_4_ & P4_DATAO_REG_5_;
  assign n44240 = n44119 & n44239;
  assign n44241 = ~n44237 & ~n44238;
  assign n44242 = ~n44240 & n44241;
  assign n44243 = n44238 & n44240;
  assign n44244 = n44231 & n44240;
  assign n44245 = ~n44236 & n44244;
  assign n44246 = ~n44242 & ~n44243;
  assign n44247 = ~n44245 & n44246;
  assign n44248 = n44230 & ~n44247;
  assign n44249 = ~n44230 & n44247;
  assign n44250 = ~n44248 & ~n44249;
  assign n44251 = n44229 & ~n44250;
  assign n44252 = ~n44230 & ~n44247;
  assign n44253 = ~n44229 & n44252;
  assign n44254 = ~n44229 & n44230;
  assign n44255 = n44247 & n44254;
  assign n44256 = ~n44251 & ~n44253;
  assign n44257 = ~n44255 & n44256;
  assign n44258 = n44226 & ~n44257;
  assign n44259 = ~n44226 & n44257;
  assign n44260 = ~n44258 & ~n44259;
  assign n44261 = ~n44146 & ~n44164;
  assign n44262 = ~n44165 & ~n44171;
  assign n44263 = ~n44261 & n44262;
  assign n44264 = ~n44260 & n44263;
  assign n44265 = ~n44226 & ~n44257;
  assign n44266 = ~n44263 & n44265;
  assign n44267 = n44226 & ~n44263;
  assign n44268 = n44257 & n44267;
  assign n44269 = ~n44264 & ~n44266;
  assign n44270 = ~n44268 & n44269;
  assign n44271 = n44225 & ~n44270;
  assign n44272 = ~n44225 & n44270;
  assign n44273 = ~n44271 & ~n44272;
  assign n44274 = n44224 & ~n44273;
  assign n44275 = ~n44225 & ~n44270;
  assign n44276 = ~n44224 & n44275;
  assign n44277 = ~n44224 & n44225;
  assign n44278 = n44270 & n44277;
  assign n44279 = ~n44274 & ~n44276;
  assign n44280 = ~n44278 & n44279;
  assign n44281 = ~n44103 & n44221;
  assign n44282 = n44280 & ~n44281;
  assign n44283 = ~n44222 & ~n44282;
  assign n44284 = ~n44224 & ~n44270;
  assign n44285 = ~n44271 & ~n44277;
  assign n44286 = ~n44284 & n44285;
  assign n44287 = P4_DATAO_REG_1_ & n44102;
  assign n44288 = ~n44226 & n44263;
  assign n44289 = n44257 & ~n44288;
  assign n44290 = ~n44267 & ~n44289;
  assign n44291 = P4_DATAO_REG_2_ & n44104;
  assign n44292 = P4_DATAO_REG_3_ & n44143;
  assign n44293 = ~n44231 & ~n44240;
  assign n44294 = ~n44236 & ~n44293;
  assign n44295 = ~n44244 & ~n44294;
  assign n44296 = P4_DATAO_REG_4_ & n44106;
  assign n44297 = P4_DATAO_REG_5_ & n44108;
  assign n44298 = P4_DATAO_REG_7_ & n44112;
  assign n44299 = P4_DATAO_REG_6_ & n44110;
  assign n44300 = n44298 & ~n44299;
  assign n44301 = ~n44298 & n44299;
  assign n44302 = ~n44300 & ~n44301;
  assign n44303 = n44297 & ~n44302;
  assign n44304 = ~n44297 & n44302;
  assign n44305 = P4_DATAO_REG_5_ & P4_DATAO_REG_6_;
  assign n44306 = n44119 & n44305;
  assign n44307 = ~n44303 & ~n44304;
  assign n44308 = ~n44306 & n44307;
  assign n44309 = n44304 & n44306;
  assign n44310 = n44297 & n44306;
  assign n44311 = ~n44302 & n44310;
  assign n44312 = ~n44308 & ~n44309;
  assign n44313 = ~n44311 & n44312;
  assign n44314 = n44296 & ~n44313;
  assign n44315 = ~n44296 & n44313;
  assign n44316 = ~n44314 & ~n44315;
  assign n44317 = n44295 & ~n44316;
  assign n44318 = ~n44296 & ~n44313;
  assign n44319 = ~n44295 & n44318;
  assign n44320 = ~n44295 & n44296;
  assign n44321 = n44313 & n44320;
  assign n44322 = ~n44317 & ~n44319;
  assign n44323 = ~n44321 & n44322;
  assign n44324 = n44292 & ~n44323;
  assign n44325 = ~n44292 & n44323;
  assign n44326 = ~n44324 & ~n44325;
  assign n44327 = ~n44229 & ~n44247;
  assign n44328 = ~n44248 & ~n44254;
  assign n44329 = ~n44327 & n44328;
  assign n44330 = ~n44326 & n44329;
  assign n44331 = ~n44292 & ~n44323;
  assign n44332 = ~n44329 & n44331;
  assign n44333 = n44292 & ~n44329;
  assign n44334 = n44323 & n44333;
  assign n44335 = ~n44330 & ~n44332;
  assign n44336 = ~n44334 & n44335;
  assign n44337 = n44291 & ~n44336;
  assign n44338 = ~n44291 & n44336;
  assign n44339 = ~n44337 & ~n44338;
  assign n44340 = n44290 & ~n44339;
  assign n44341 = ~n44291 & ~n44336;
  assign n44342 = ~n44290 & n44341;
  assign n44343 = ~n44290 & n44291;
  assign n44344 = n44336 & n44343;
  assign n44345 = ~n44340 & ~n44342;
  assign n44346 = ~n44344 & n44345;
  assign n44347 = n44287 & ~n44346;
  assign n44348 = ~n44287 & n44346;
  assign n44349 = ~n44347 & ~n44348;
  assign n44350 = n44286 & ~n44349;
  assign n44351 = n44287 & n44346;
  assign n44352 = ~n44287 & ~n44346;
  assign n44353 = ~n44351 & ~n44352;
  assign n44354 = ~n44286 & ~n44353;
  assign n44355 = ~n44350 & ~n44354;
  assign n44356 = SEL & DIN_7_;
  assign n44357 = P4_DATAO_REG_0_ & n44356;
  assign n44358 = ~n44355 & ~n44357;
  assign n44359 = n44355 & n44357;
  assign n44360 = ~n44358 & ~n44359;
  assign n44361 = n44283 & ~n44360;
  assign n44362 = n44355 & ~n44357;
  assign n44363 = ~n44355 & n44357;
  assign n44364 = ~n44362 & ~n44363;
  assign n44365 = ~n44283 & ~n44364;
  assign n44366 = ~n44361 & ~n44365;
  assign n44367 = ~n12460 & ~n44366;
  assign n44368 = ~n44101 & ~n44367;
  assign n44369 = n44042 & ~n44368;
  assign n44370 = n44100 & n44369;
  assign n44371 = P1_BUF1_REG_23_ & n12460;
  assign n44372 = SEL & DIN_23_;
  assign n44373 = P4_DATAO_REG_0_ & n44372;
  assign n44374 = SEL & DIN_21_;
  assign n44375 = P4_DATAO_REG_1_ & n44374;
  assign n44376 = SEL & DIN_20_;
  assign n44377 = P4_DATAO_REG_1_ & n44376;
  assign n44378 = SEL & DIN_19_;
  assign n44379 = P4_DATAO_REG_1_ & n44378;
  assign n44380 = SEL & DIN_18_;
  assign n44381 = P4_DATAO_REG_2_ & n44380;
  assign n44382 = SEL & DIN_17_;
  assign n44383 = P4_DATAO_REG_2_ & n44382;
  assign n44384 = SEL & DIN_15_;
  assign n44385 = P4_DATAO_REG_4_ & n44384;
  assign n44386 = SEL & DIN_14_;
  assign n44387 = P4_DATAO_REG_4_ & n44386;
  assign n44388 = SEL & DIN_13_;
  assign n44389 = P4_DATAO_REG_5_ & n44388;
  assign n44390 = SEL & DIN_12_;
  assign n44391 = P4_DATAO_REG_5_ & n44390;
  assign n44392 = SEL & DIN_11_;
  assign n44393 = P4_DATAO_REG_6_ & n44392;
  assign n44394 = SEL & DIN_10_;
  assign n44395 = P4_DATAO_REG_6_ & n44394;
  assign n44396 = P4_DATAO_REG_13_ & n44106;
  assign n44397 = P4_DATAO_REG_13_ & n44108;
  assign n44398 = P4_DATAO_REG_14_ & n44110;
  assign n44399 = P4_DATAO_REG_15_ & n44112;
  assign n44400 = n44398 & ~n44399;
  assign n44401 = ~n44398 & n44399;
  assign n44402 = ~n44400 & ~n44401;
  assign n44403 = n44397 & ~n44402;
  assign n44404 = P4_DATAO_REG_13_ & P4_DATAO_REG_14_;
  assign n44405 = n44119 & n44404;
  assign n44406 = ~n44397 & n44402;
  assign n44407 = n44405 & ~n44406;
  assign n44408 = ~n44403 & ~n44407;
  assign n44409 = n44396 & ~n44408;
  assign n44410 = ~n44396 & n44408;
  assign n44411 = ~n44409 & ~n44410;
  assign n44412 = P4_DATAO_REG_14_ & n44108;
  assign n44413 = P4_DATAO_REG_15_ & n44110;
  assign n44414 = P4_DATAO_REG_16_ & n44112;
  assign n44415 = n44413 & ~n44414;
  assign n44416 = ~n44413 & n44414;
  assign n44417 = ~n44415 & ~n44416;
  assign n44418 = n44412 & ~n44417;
  assign n44419 = ~n44412 & n44417;
  assign n44420 = P4_DATAO_REG_14_ & P4_DATAO_REG_15_;
  assign n44421 = n44119 & n44420;
  assign n44422 = ~n44418 & ~n44419;
  assign n44423 = ~n44421 & n44422;
  assign n44424 = n44421 & ~n44422;
  assign n44425 = ~n44423 & ~n44424;
  assign n44426 = ~n44411 & n44425;
  assign n44427 = n44411 & ~n44425;
  assign n44428 = ~n44426 & ~n44427;
  assign n44429 = P4_DATAO_REG_12_ & n44143;
  assign n44430 = ~n44428 & ~n44429;
  assign n44431 = n44428 & n44429;
  assign n44432 = P4_DATAO_REG_12_ & n44106;
  assign n44433 = P4_DATAO_REG_12_ & n44108;
  assign n44434 = P4_DATAO_REG_13_ & n44110;
  assign n44435 = P4_DATAO_REG_14_ & n44112;
  assign n44436 = n44434 & ~n44435;
  assign n44437 = ~n44434 & n44435;
  assign n44438 = ~n44436 & ~n44437;
  assign n44439 = n44433 & ~n44438;
  assign n44440 = P4_DATAO_REG_12_ & P4_DATAO_REG_13_;
  assign n44441 = n44119 & n44440;
  assign n44442 = ~n44433 & n44438;
  assign n44443 = n44441 & ~n44442;
  assign n44444 = ~n44439 & ~n44443;
  assign n44445 = n44432 & ~n44444;
  assign n44446 = ~n44403 & ~n44406;
  assign n44447 = ~n44405 & n44446;
  assign n44448 = n44405 & ~n44446;
  assign n44449 = ~n44447 & ~n44448;
  assign n44450 = n44432 & ~n44449;
  assign n44451 = ~n44444 & ~n44449;
  assign n44452 = ~n44445 & ~n44450;
  assign n44453 = ~n44451 & n44452;
  assign n44454 = ~n44430 & ~n44431;
  assign n44455 = n44453 & n44454;
  assign n44456 = ~n44453 & ~n44454;
  assign n44457 = ~n44455 & ~n44456;
  assign n44458 = P4_DATAO_REG_11_ & n44104;
  assign n44459 = n44457 & n44458;
  assign n44460 = ~n44457 & ~n44458;
  assign n44461 = ~n44459 & ~n44460;
  assign n44462 = P4_DATAO_REG_11_ & n44143;
  assign n44463 = ~n44432 & n44449;
  assign n44464 = ~n44450 & ~n44463;
  assign n44465 = n44444 & ~n44464;
  assign n44466 = ~n44432 & ~n44449;
  assign n44467 = ~n44444 & n44466;
  assign n44468 = n44445 & n44449;
  assign n44469 = ~n44465 & ~n44467;
  assign n44470 = ~n44468 & n44469;
  assign n44471 = n44462 & n44470;
  assign n44472 = ~n44462 & ~n44470;
  assign n44473 = P4_DATAO_REG_11_ & n44106;
  assign n44474 = P4_DATAO_REG_11_ & n44108;
  assign n44475 = P4_DATAO_REG_12_ & n44110;
  assign n44476 = P4_DATAO_REG_13_ & n44112;
  assign n44477 = n44475 & ~n44476;
  assign n44478 = ~n44475 & n44476;
  assign n44479 = ~n44477 & ~n44478;
  assign n44480 = n44474 & ~n44479;
  assign n44481 = P4_DATAO_REG_11_ & P4_DATAO_REG_12_;
  assign n44482 = n44119 & n44481;
  assign n44483 = ~n44474 & n44479;
  assign n44484 = n44482 & ~n44483;
  assign n44485 = ~n44480 & ~n44484;
  assign n44486 = n44473 & ~n44485;
  assign n44487 = ~n44439 & ~n44442;
  assign n44488 = ~n44441 & n44487;
  assign n44489 = n44441 & ~n44487;
  assign n44490 = ~n44488 & ~n44489;
  assign n44491 = n44473 & ~n44490;
  assign n44492 = ~n44485 & ~n44490;
  assign n44493 = ~n44486 & ~n44491;
  assign n44494 = ~n44492 & n44493;
  assign n44495 = ~n44472 & ~n44494;
  assign n44496 = ~n44471 & ~n44495;
  assign n44497 = ~n44461 & ~n44496;
  assign n44498 = n44461 & n44496;
  assign n44499 = ~n44497 & ~n44498;
  assign n44500 = P4_DATAO_REG_10_ & n44102;
  assign n44501 = ~n44499 & ~n44500;
  assign n44502 = n44499 & n44500;
  assign n44503 = P4_DATAO_REG_10_ & n44104;
  assign n44504 = P4_DATAO_REG_10_ & n44143;
  assign n44505 = ~n44473 & n44490;
  assign n44506 = ~n44491 & ~n44505;
  assign n44507 = n44485 & ~n44506;
  assign n44508 = ~n44473 & ~n44490;
  assign n44509 = ~n44485 & n44508;
  assign n44510 = n44486 & n44490;
  assign n44511 = ~n44507 & ~n44509;
  assign n44512 = ~n44510 & n44511;
  assign n44513 = n44504 & n44512;
  assign n44514 = ~n44504 & ~n44512;
  assign n44515 = P4_DATAO_REG_10_ & n44106;
  assign n44516 = P4_DATAO_REG_10_ & n44108;
  assign n44517 = P4_DATAO_REG_11_ & n44110;
  assign n44518 = P4_DATAO_REG_12_ & n44112;
  assign n44519 = n44517 & ~n44518;
  assign n44520 = ~n44517 & n44518;
  assign n44521 = ~n44519 & ~n44520;
  assign n44522 = n44516 & ~n44521;
  assign n44523 = P4_DATAO_REG_10_ & P4_DATAO_REG_11_;
  assign n44524 = n44119 & n44523;
  assign n44525 = ~n44516 & n44521;
  assign n44526 = n44524 & ~n44525;
  assign n44527 = ~n44522 & ~n44526;
  assign n44528 = n44515 & ~n44527;
  assign n44529 = ~n44480 & ~n44483;
  assign n44530 = ~n44482 & n44529;
  assign n44531 = n44482 & ~n44529;
  assign n44532 = ~n44530 & ~n44531;
  assign n44533 = n44515 & ~n44532;
  assign n44534 = ~n44527 & ~n44532;
  assign n44535 = ~n44528 & ~n44533;
  assign n44536 = ~n44534 & n44535;
  assign n44537 = ~n44514 & ~n44536;
  assign n44538 = ~n44513 & ~n44537;
  assign n44539 = n44503 & ~n44538;
  assign n44540 = n44462 & ~n44470;
  assign n44541 = ~n44462 & n44470;
  assign n44542 = ~n44540 & ~n44541;
  assign n44543 = n44494 & ~n44542;
  assign n44544 = ~n44471 & ~n44472;
  assign n44545 = ~n44494 & ~n44544;
  assign n44546 = ~n44543 & ~n44545;
  assign n44547 = n44503 & ~n44546;
  assign n44548 = ~n44538 & ~n44546;
  assign n44549 = ~n44539 & ~n44547;
  assign n44550 = ~n44548 & n44549;
  assign n44551 = ~n44501 & ~n44502;
  assign n44552 = n44550 & n44551;
  assign n44553 = ~n44550 & ~n44551;
  assign n44554 = ~n44552 & ~n44553;
  assign n44555 = P4_DATAO_REG_9_ & n44356;
  assign n44556 = n44554 & n44555;
  assign n44557 = ~n44554 & ~n44555;
  assign n44558 = ~n44556 & ~n44557;
  assign n44559 = ~n44503 & n44546;
  assign n44560 = ~n44547 & ~n44559;
  assign n44561 = n44538 & ~n44560;
  assign n44562 = ~n44503 & ~n44546;
  assign n44563 = ~n44538 & n44562;
  assign n44564 = n44539 & n44546;
  assign n44565 = ~n44561 & ~n44563;
  assign n44566 = ~n44564 & n44565;
  assign n44567 = P4_DATAO_REG_9_ & n44102;
  assign n44568 = n44566 & n44567;
  assign n44569 = ~n44566 & ~n44567;
  assign n44570 = P4_DATAO_REG_9_ & n44104;
  assign n44571 = ~n44515 & n44532;
  assign n44572 = ~n44533 & ~n44571;
  assign n44573 = n44527 & ~n44572;
  assign n44574 = ~n44515 & ~n44532;
  assign n44575 = ~n44527 & n44574;
  assign n44576 = n44528 & n44532;
  assign n44577 = ~n44573 & ~n44575;
  assign n44578 = ~n44576 & n44577;
  assign n44579 = P4_DATAO_REG_9_ & n44143;
  assign n44580 = n44578 & n44579;
  assign n44581 = ~n44578 & ~n44579;
  assign n44582 = P4_DATAO_REG_9_ & n44106;
  assign n44583 = P4_DATAO_REG_9_ & n44108;
  assign n44584 = P4_DATAO_REG_10_ & n44110;
  assign n44585 = P4_DATAO_REG_11_ & n44112;
  assign n44586 = n44584 & ~n44585;
  assign n44587 = ~n44584 & n44585;
  assign n44588 = ~n44586 & ~n44587;
  assign n44589 = n44583 & ~n44588;
  assign n44590 = P4_DATAO_REG_9_ & P4_DATAO_REG_10_;
  assign n44591 = n44119 & n44590;
  assign n44592 = ~n44583 & n44588;
  assign n44593 = n44591 & ~n44592;
  assign n44594 = ~n44589 & ~n44593;
  assign n44595 = n44582 & ~n44594;
  assign n44596 = ~n44522 & ~n44525;
  assign n44597 = ~n44524 & n44596;
  assign n44598 = n44524 & ~n44596;
  assign n44599 = ~n44597 & ~n44598;
  assign n44600 = n44582 & ~n44599;
  assign n44601 = ~n44594 & ~n44599;
  assign n44602 = ~n44595 & ~n44600;
  assign n44603 = ~n44601 & n44602;
  assign n44604 = ~n44581 & ~n44603;
  assign n44605 = ~n44580 & ~n44604;
  assign n44606 = n44570 & ~n44605;
  assign n44607 = n44504 & ~n44512;
  assign n44608 = ~n44504 & n44512;
  assign n44609 = ~n44607 & ~n44608;
  assign n44610 = n44536 & ~n44609;
  assign n44611 = ~n44513 & ~n44514;
  assign n44612 = ~n44536 & ~n44611;
  assign n44613 = ~n44610 & ~n44612;
  assign n44614 = n44570 & ~n44613;
  assign n44615 = ~n44605 & ~n44613;
  assign n44616 = ~n44606 & ~n44614;
  assign n44617 = ~n44615 & n44616;
  assign n44618 = ~n44569 & ~n44617;
  assign n44619 = ~n44568 & ~n44618;
  assign n44620 = ~n44558 & ~n44619;
  assign n44621 = n44558 & n44619;
  assign n44622 = ~n44620 & ~n44621;
  assign n44623 = SEL & DIN_8_;
  assign n44624 = P4_DATAO_REG_8_ & n44623;
  assign n44625 = ~n44622 & ~n44624;
  assign n44626 = n44622 & n44624;
  assign n44627 = P4_DATAO_REG_8_ & n44356;
  assign n44628 = ~n44566 & n44567;
  assign n44629 = n44566 & ~n44567;
  assign n44630 = ~n44628 & ~n44629;
  assign n44631 = n44617 & ~n44630;
  assign n44632 = ~n44568 & ~n44569;
  assign n44633 = ~n44617 & ~n44632;
  assign n44634 = ~n44631 & ~n44633;
  assign n44635 = n44627 & ~n44634;
  assign n44636 = ~n44627 & n44634;
  assign n44637 = P4_DATAO_REG_8_ & n44102;
  assign n44638 = P4_DATAO_REG_8_ & n44104;
  assign n44639 = ~n44578 & n44579;
  assign n44640 = n44578 & ~n44579;
  assign n44641 = ~n44639 & ~n44640;
  assign n44642 = n44603 & ~n44641;
  assign n44643 = ~n44580 & ~n44581;
  assign n44644 = ~n44603 & ~n44643;
  assign n44645 = ~n44642 & ~n44644;
  assign n44646 = n44638 & ~n44645;
  assign n44647 = ~n44582 & n44599;
  assign n44648 = ~n44600 & ~n44647;
  assign n44649 = n44594 & ~n44648;
  assign n44650 = ~n44582 & ~n44599;
  assign n44651 = ~n44594 & n44650;
  assign n44652 = n44595 & n44599;
  assign n44653 = ~n44649 & ~n44651;
  assign n44654 = ~n44652 & n44653;
  assign n44655 = P4_DATAO_REG_8_ & n44143;
  assign n44656 = n44654 & n44655;
  assign n44657 = ~n44654 & ~n44655;
  assign n44658 = P4_DATAO_REG_8_ & n44106;
  assign n44659 = P4_DATAO_REG_8_ & n44108;
  assign n44660 = P4_DATAO_REG_9_ & n44110;
  assign n44661 = P4_DATAO_REG_10_ & n44112;
  assign n44662 = n44660 & ~n44661;
  assign n44663 = ~n44660 & n44661;
  assign n44664 = ~n44662 & ~n44663;
  assign n44665 = n44659 & ~n44664;
  assign n44666 = P4_DATAO_REG_8_ & P4_DATAO_REG_9_;
  assign n44667 = n44119 & n44666;
  assign n44668 = ~n44659 & n44664;
  assign n44669 = n44667 & ~n44668;
  assign n44670 = ~n44665 & ~n44669;
  assign n44671 = n44658 & ~n44670;
  assign n44672 = ~n44589 & ~n44592;
  assign n44673 = ~n44591 & n44672;
  assign n44674 = n44591 & ~n44672;
  assign n44675 = ~n44673 & ~n44674;
  assign n44676 = n44658 & ~n44675;
  assign n44677 = ~n44670 & ~n44675;
  assign n44678 = ~n44671 & ~n44676;
  assign n44679 = ~n44677 & n44678;
  assign n44680 = ~n44657 & ~n44679;
  assign n44681 = ~n44656 & ~n44680;
  assign n44682 = n44638 & ~n44681;
  assign n44683 = ~n44645 & ~n44681;
  assign n44684 = ~n44646 & ~n44682;
  assign n44685 = ~n44683 & n44684;
  assign n44686 = n44637 & ~n44685;
  assign n44687 = ~n44570 & n44613;
  assign n44688 = ~n44614 & ~n44687;
  assign n44689 = n44605 & ~n44688;
  assign n44690 = ~n44570 & ~n44613;
  assign n44691 = ~n44605 & n44690;
  assign n44692 = n44606 & n44613;
  assign n44693 = ~n44689 & ~n44691;
  assign n44694 = ~n44692 & n44693;
  assign n44695 = ~n44637 & n44685;
  assign n44696 = n44694 & ~n44695;
  assign n44697 = ~n44686 & ~n44696;
  assign n44698 = ~n44636 & ~n44697;
  assign n44699 = ~n44635 & ~n44698;
  assign n44700 = ~n44625 & ~n44626;
  assign n44701 = n44699 & n44700;
  assign n44702 = ~n44699 & ~n44700;
  assign n44703 = ~n44701 & ~n44702;
  assign n44704 = SEL & DIN_9_;
  assign n44705 = P4_DATAO_REG_7_ & n44704;
  assign n44706 = n44703 & n44705;
  assign n44707 = ~n44703 & ~n44705;
  assign n44708 = ~n44706 & ~n44707;
  assign n44709 = P4_DATAO_REG_7_ & n44623;
  assign n44710 = n44627 & ~n44697;
  assign n44711 = ~n44627 & n44697;
  assign n44712 = ~n44710 & ~n44711;
  assign n44713 = n44634 & ~n44712;
  assign n44714 = ~n44634 & n44712;
  assign n44715 = ~n44713 & ~n44714;
  assign n44716 = n44709 & n44715;
  assign n44717 = ~n44709 & ~n44715;
  assign n44718 = P4_DATAO_REG_7_ & n44356;
  assign n44719 = ~n44638 & n44681;
  assign n44720 = ~n44682 & ~n44719;
  assign n44721 = n44645 & ~n44720;
  assign n44722 = ~n44638 & ~n44681;
  assign n44723 = ~n44645 & n44722;
  assign n44724 = n44646 & n44681;
  assign n44725 = ~n44721 & ~n44723;
  assign n44726 = ~n44724 & n44725;
  assign n44727 = P4_DATAO_REG_7_ & n44102;
  assign n44728 = n44726 & n44727;
  assign n44729 = ~n44726 & ~n44727;
  assign n44730 = P4_DATAO_REG_7_ & n44104;
  assign n44731 = ~n44658 & n44675;
  assign n44732 = ~n44676 & ~n44731;
  assign n44733 = n44670 & ~n44732;
  assign n44734 = ~n44658 & ~n44675;
  assign n44735 = ~n44670 & n44734;
  assign n44736 = n44671 & n44675;
  assign n44737 = ~n44733 & ~n44735;
  assign n44738 = ~n44736 & n44737;
  assign n44739 = P4_DATAO_REG_7_ & n44143;
  assign n44740 = n44738 & n44739;
  assign n44741 = ~n44738 & ~n44739;
  assign n44742 = P4_DATAO_REG_7_ & n44106;
  assign n44743 = P4_DATAO_REG_7_ & P4_DATAO_REG_8_;
  assign n44744 = n44119 & n44743;
  assign n44745 = P4_DATAO_REG_7_ & n44108;
  assign n44746 = n44744 & n44745;
  assign n44747 = ~n44744 & ~n44745;
  assign n44748 = P4_DATAO_REG_9_ & n44112;
  assign n44749 = P4_DATAO_REG_8_ & n44110;
  assign n44750 = n44748 & ~n44749;
  assign n44751 = ~n44748 & n44749;
  assign n44752 = ~n44750 & ~n44751;
  assign n44753 = ~n44747 & ~n44752;
  assign n44754 = ~n44746 & ~n44753;
  assign n44755 = n44742 & ~n44754;
  assign n44756 = ~n44665 & ~n44668;
  assign n44757 = ~n44667 & n44756;
  assign n44758 = n44667 & ~n44756;
  assign n44759 = ~n44757 & ~n44758;
  assign n44760 = n44742 & ~n44759;
  assign n44761 = ~n44754 & ~n44759;
  assign n44762 = ~n44755 & ~n44760;
  assign n44763 = ~n44761 & n44762;
  assign n44764 = ~n44741 & ~n44763;
  assign n44765 = ~n44740 & ~n44764;
  assign n44766 = n44730 & ~n44765;
  assign n44767 = ~n44654 & n44655;
  assign n44768 = n44654 & ~n44655;
  assign n44769 = ~n44767 & ~n44768;
  assign n44770 = n44679 & ~n44769;
  assign n44771 = ~n44656 & ~n44657;
  assign n44772 = ~n44679 & ~n44771;
  assign n44773 = ~n44770 & ~n44772;
  assign n44774 = n44730 & ~n44773;
  assign n44775 = ~n44765 & ~n44773;
  assign n44776 = ~n44766 & ~n44774;
  assign n44777 = ~n44775 & n44776;
  assign n44778 = ~n44729 & ~n44777;
  assign n44779 = ~n44728 & ~n44778;
  assign n44780 = n44718 & ~n44779;
  assign n44781 = ~n44686 & ~n44695;
  assign n44782 = ~n44694 & n44781;
  assign n44783 = n44694 & ~n44781;
  assign n44784 = ~n44782 & ~n44783;
  assign n44785 = n44718 & ~n44784;
  assign n44786 = ~n44779 & ~n44784;
  assign n44787 = ~n44780 & ~n44785;
  assign n44788 = ~n44786 & n44787;
  assign n44789 = ~n44717 & ~n44788;
  assign n44790 = ~n44716 & ~n44789;
  assign n44791 = ~n44708 & ~n44790;
  assign n44792 = n44708 & n44790;
  assign n44793 = ~n44791 & ~n44792;
  assign n44794 = n44395 & n44793;
  assign n44795 = ~n44395 & ~n44793;
  assign n44796 = P4_DATAO_REG_6_ & n44704;
  assign n44797 = ~n44718 & n44784;
  assign n44798 = ~n44785 & ~n44797;
  assign n44799 = n44779 & ~n44798;
  assign n44800 = ~n44718 & ~n44784;
  assign n44801 = ~n44779 & n44800;
  assign n44802 = n44780 & n44784;
  assign n44803 = ~n44799 & ~n44801;
  assign n44804 = ~n44802 & n44803;
  assign n44805 = P4_DATAO_REG_6_ & n44623;
  assign n44806 = n44804 & n44805;
  assign n44807 = ~n44804 & ~n44805;
  assign n44808 = P4_DATAO_REG_6_ & n44356;
  assign n44809 = ~n44726 & n44727;
  assign n44810 = n44726 & ~n44727;
  assign n44811 = ~n44809 & ~n44810;
  assign n44812 = n44777 & ~n44811;
  assign n44813 = ~n44728 & ~n44729;
  assign n44814 = ~n44777 & ~n44813;
  assign n44815 = ~n44812 & ~n44814;
  assign n44816 = n44808 & ~n44815;
  assign n44817 = ~n44730 & n44773;
  assign n44818 = ~n44774 & ~n44817;
  assign n44819 = n44765 & ~n44818;
  assign n44820 = ~n44730 & ~n44773;
  assign n44821 = ~n44765 & n44820;
  assign n44822 = n44766 & n44773;
  assign n44823 = ~n44819 & ~n44821;
  assign n44824 = ~n44822 & n44823;
  assign n44825 = P4_DATAO_REG_6_ & n44102;
  assign n44826 = n44824 & n44825;
  assign n44827 = ~n44824 & ~n44825;
  assign n44828 = P4_DATAO_REG_6_ & n44104;
  assign n44829 = ~n44738 & n44739;
  assign n44830 = n44738 & ~n44739;
  assign n44831 = ~n44829 & ~n44830;
  assign n44832 = n44763 & ~n44831;
  assign n44833 = ~n44740 & ~n44741;
  assign n44834 = ~n44763 & ~n44833;
  assign n44835 = ~n44832 & ~n44834;
  assign n44836 = n44828 & ~n44835;
  assign n44837 = ~n44742 & n44759;
  assign n44838 = ~n44760 & ~n44837;
  assign n44839 = n44754 & ~n44838;
  assign n44840 = ~n44742 & ~n44759;
  assign n44841 = ~n44754 & n44840;
  assign n44842 = n44755 & n44759;
  assign n44843 = ~n44839 & ~n44841;
  assign n44844 = ~n44842 & n44843;
  assign n44845 = P4_DATAO_REG_6_ & n44143;
  assign n44846 = n44844 & n44845;
  assign n44847 = ~n44844 & ~n44845;
  assign n44848 = P4_DATAO_REG_6_ & n44106;
  assign n44849 = n44745 & ~n44752;
  assign n44850 = ~n44745 & n44752;
  assign n44851 = ~n44849 & ~n44850;
  assign n44852 = ~n44744 & n44851;
  assign n44853 = n44744 & n44850;
  assign n44854 = n44746 & ~n44752;
  assign n44855 = ~n44852 & ~n44853;
  assign n44856 = ~n44854 & n44855;
  assign n44857 = n44848 & ~n44856;
  assign n44858 = P4_DATAO_REG_6_ & P4_DATAO_REG_7_;
  assign n44859 = n44119 & n44858;
  assign n44860 = P4_DATAO_REG_6_ & n44108;
  assign n44861 = n44859 & n44860;
  assign n44862 = ~n44859 & ~n44860;
  assign n44863 = P4_DATAO_REG_8_ & n44112;
  assign n44864 = P4_DATAO_REG_7_ & n44110;
  assign n44865 = n44863 & ~n44864;
  assign n44866 = ~n44863 & n44864;
  assign n44867 = ~n44865 & ~n44866;
  assign n44868 = ~n44862 & ~n44867;
  assign n44869 = ~n44861 & ~n44868;
  assign n44870 = n44848 & ~n44869;
  assign n44871 = ~n44856 & ~n44869;
  assign n44872 = ~n44857 & ~n44870;
  assign n44873 = ~n44871 & n44872;
  assign n44874 = ~n44847 & ~n44873;
  assign n44875 = ~n44846 & ~n44874;
  assign n44876 = n44828 & ~n44875;
  assign n44877 = ~n44835 & ~n44875;
  assign n44878 = ~n44836 & ~n44876;
  assign n44879 = ~n44877 & n44878;
  assign n44880 = ~n44827 & ~n44879;
  assign n44881 = ~n44826 & ~n44880;
  assign n44882 = n44808 & ~n44881;
  assign n44883 = ~n44815 & ~n44881;
  assign n44884 = ~n44816 & ~n44882;
  assign n44885 = ~n44883 & n44884;
  assign n44886 = ~n44807 & ~n44885;
  assign n44887 = ~n44806 & ~n44886;
  assign n44888 = n44796 & ~n44887;
  assign n44889 = ~n44716 & ~n44717;
  assign n44890 = n44788 & n44889;
  assign n44891 = ~n44788 & ~n44889;
  assign n44892 = ~n44890 & ~n44891;
  assign n44893 = n44796 & ~n44892;
  assign n44894 = ~n44887 & ~n44892;
  assign n44895 = ~n44888 & ~n44893;
  assign n44896 = ~n44894 & n44895;
  assign n44897 = ~n44795 & ~n44896;
  assign n44898 = ~n44794 & ~n44897;
  assign n44899 = n44393 & ~n44898;
  assign n44900 = ~n44393 & n44898;
  assign n44901 = ~n44899 & ~n44900;
  assign n44902 = ~n44703 & n44705;
  assign n44903 = n44703 & ~n44705;
  assign n44904 = ~n44790 & ~n44903;
  assign n44905 = ~n44902 & ~n44904;
  assign n44906 = P4_DATAO_REG_7_ & n44394;
  assign n44907 = ~n44625 & ~n44699;
  assign n44908 = ~n44626 & ~n44907;
  assign n44909 = P4_DATAO_REG_8_ & n44704;
  assign n44910 = P4_DATAO_REG_9_ & n44623;
  assign n44911 = ~n44554 & n44555;
  assign n44912 = n44554 & ~n44555;
  assign n44913 = ~n44619 & ~n44912;
  assign n44914 = ~n44911 & ~n44913;
  assign n44915 = n44910 & ~n44914;
  assign n44916 = ~n44910 & n44914;
  assign n44917 = ~n44915 & ~n44916;
  assign n44918 = ~n44501 & ~n44550;
  assign n44919 = ~n44502 & ~n44918;
  assign n44920 = P4_DATAO_REG_10_ & n44356;
  assign n44921 = ~n44457 & n44458;
  assign n44922 = n44457 & ~n44458;
  assign n44923 = ~n44496 & ~n44922;
  assign n44924 = ~n44921 & ~n44923;
  assign n44925 = P4_DATAO_REG_11_ & n44102;
  assign n44926 = ~n44430 & ~n44453;
  assign n44927 = ~n44431 & ~n44926;
  assign n44928 = P4_DATAO_REG_12_ & n44104;
  assign n44929 = n44396 & ~n44425;
  assign n44930 = ~n44396 & n44425;
  assign n44931 = ~n44408 & ~n44930;
  assign n44932 = ~n44929 & ~n44931;
  assign n44933 = P4_DATAO_REG_13_ & n44143;
  assign n44934 = ~n44419 & n44421;
  assign n44935 = ~n44418 & ~n44934;
  assign n44936 = P4_DATAO_REG_14_ & n44106;
  assign n44937 = P4_DATAO_REG_16_ & n44110;
  assign n44938 = P4_DATAO_REG_17_ & n44112;
  assign n44939 = n44937 & ~n44938;
  assign n44940 = ~n44937 & n44938;
  assign n44941 = ~n44939 & ~n44940;
  assign n44942 = P4_DATAO_REG_15_ & n44108;
  assign n44943 = P4_DATAO_REG_15_ & P4_DATAO_REG_16_;
  assign n44944 = n44119 & n44943;
  assign n44945 = n44942 & ~n44944;
  assign n44946 = ~n44942 & n44944;
  assign n44947 = ~n44945 & ~n44946;
  assign n44948 = n44941 & ~n44947;
  assign n44949 = ~n44942 & ~n44944;
  assign n44950 = n44942 & n44944;
  assign n44951 = ~n44949 & ~n44950;
  assign n44952 = ~n44941 & ~n44951;
  assign n44953 = ~n44948 & ~n44952;
  assign n44954 = n44936 & ~n44953;
  assign n44955 = ~n44936 & n44953;
  assign n44956 = ~n44954 & ~n44955;
  assign n44957 = n44935 & ~n44956;
  assign n44958 = ~n44936 & ~n44953;
  assign n44959 = ~n44935 & n44958;
  assign n44960 = ~n44935 & n44936;
  assign n44961 = n44953 & n44960;
  assign n44962 = ~n44957 & ~n44959;
  assign n44963 = ~n44961 & n44962;
  assign n44964 = n44933 & ~n44963;
  assign n44965 = ~n44933 & n44963;
  assign n44966 = ~n44964 & ~n44965;
  assign n44967 = n44932 & ~n44966;
  assign n44968 = n44933 & n44963;
  assign n44969 = ~n44933 & ~n44963;
  assign n44970 = ~n44968 & ~n44969;
  assign n44971 = ~n44932 & ~n44970;
  assign n44972 = ~n44967 & ~n44971;
  assign n44973 = n44928 & ~n44972;
  assign n44974 = ~n44928 & n44972;
  assign n44975 = ~n44973 & ~n44974;
  assign n44976 = n44927 & ~n44975;
  assign n44977 = ~n44928 & ~n44972;
  assign n44978 = ~n44927 & n44977;
  assign n44979 = ~n44927 & n44928;
  assign n44980 = n44972 & n44979;
  assign n44981 = ~n44976 & ~n44978;
  assign n44982 = ~n44980 & n44981;
  assign n44983 = n44925 & ~n44982;
  assign n44984 = ~n44925 & n44982;
  assign n44985 = ~n44983 & ~n44984;
  assign n44986 = n44924 & ~n44985;
  assign n44987 = n44925 & n44982;
  assign n44988 = ~n44925 & ~n44982;
  assign n44989 = ~n44987 & ~n44988;
  assign n44990 = ~n44924 & ~n44989;
  assign n44991 = ~n44986 & ~n44990;
  assign n44992 = n44920 & ~n44991;
  assign n44993 = ~n44920 & n44991;
  assign n44994 = ~n44992 & ~n44993;
  assign n44995 = n44919 & ~n44994;
  assign n44996 = ~n44920 & ~n44991;
  assign n44997 = ~n44919 & n44996;
  assign n44998 = ~n44919 & n44920;
  assign n44999 = n44991 & n44998;
  assign n45000 = ~n44995 & ~n44997;
  assign n45001 = ~n44999 & n45000;
  assign n45002 = ~n44917 & ~n45001;
  assign n45003 = n44917 & n45001;
  assign n45004 = ~n45002 & ~n45003;
  assign n45005 = n44909 & n45004;
  assign n45006 = ~n44909 & ~n45004;
  assign n45007 = ~n45005 & ~n45006;
  assign n45008 = n44908 & ~n45007;
  assign n45009 = ~n44909 & n45004;
  assign n45010 = ~n44908 & n45009;
  assign n45011 = ~n44908 & n44909;
  assign n45012 = ~n45004 & n45011;
  assign n45013 = ~n45008 & ~n45010;
  assign n45014 = ~n45012 & n45013;
  assign n45015 = n44906 & ~n45014;
  assign n45016 = ~n44906 & n45014;
  assign n45017 = ~n45015 & ~n45016;
  assign n45018 = n44905 & ~n45017;
  assign n45019 = n44906 & n45014;
  assign n45020 = ~n44906 & ~n45014;
  assign n45021 = ~n45019 & ~n45020;
  assign n45022 = ~n44905 & ~n45021;
  assign n45023 = ~n45018 & ~n45022;
  assign n45024 = ~n44901 & n45023;
  assign n45025 = n44901 & ~n45023;
  assign n45026 = ~n45024 & ~n45025;
  assign n45027 = n44391 & n45026;
  assign n45028 = ~n44391 & ~n45026;
  assign n45029 = P4_DATAO_REG_5_ & n44392;
  assign n45030 = ~n44796 & n44892;
  assign n45031 = ~n44893 & ~n45030;
  assign n45032 = n44887 & ~n45031;
  assign n45033 = ~n44796 & ~n44892;
  assign n45034 = ~n44887 & n45033;
  assign n45035 = n44888 & n44892;
  assign n45036 = ~n45032 & ~n45034;
  assign n45037 = ~n45035 & n45036;
  assign n45038 = P4_DATAO_REG_5_ & n44394;
  assign n45039 = n45037 & n45038;
  assign n45040 = ~n45037 & ~n45038;
  assign n45041 = P4_DATAO_REG_5_ & n44704;
  assign n45042 = ~n44808 & n44881;
  assign n45043 = ~n44882 & ~n45042;
  assign n45044 = n44815 & ~n45043;
  assign n45045 = ~n44808 & ~n44881;
  assign n45046 = ~n44815 & n45045;
  assign n45047 = n44816 & n44881;
  assign n45048 = ~n45044 & ~n45046;
  assign n45049 = ~n45047 & n45048;
  assign n45050 = P4_DATAO_REG_5_ & n44623;
  assign n45051 = n45049 & n45050;
  assign n45052 = ~n45049 & ~n45050;
  assign n45053 = P4_DATAO_REG_5_ & n44356;
  assign n45054 = ~n44828 & n44875;
  assign n45055 = ~n44876 & ~n45054;
  assign n45056 = n44835 & ~n45055;
  assign n45057 = ~n44828 & ~n44875;
  assign n45058 = ~n44835 & n45057;
  assign n45059 = n44836 & n44875;
  assign n45060 = ~n45056 & ~n45058;
  assign n45061 = ~n45059 & n45060;
  assign n45062 = P4_DATAO_REG_5_ & n44102;
  assign n45063 = n45061 & n45062;
  assign n45064 = ~n45061 & ~n45062;
  assign n45065 = P4_DATAO_REG_5_ & n44104;
  assign n45066 = P4_DATAO_REG_5_ & n44143;
  assign n45067 = P4_DATAO_REG_5_ & n44106;
  assign n45068 = n44860 & ~n44867;
  assign n45069 = ~n44860 & n44867;
  assign n45070 = ~n45068 & ~n45069;
  assign n45071 = ~n44859 & n45070;
  assign n45072 = n44859 & n45069;
  assign n45073 = n44861 & ~n44867;
  assign n45074 = ~n45071 & ~n45072;
  assign n45075 = ~n45073 & n45074;
  assign n45076 = n45067 & ~n45075;
  assign n45077 = ~n44297 & ~n44306;
  assign n45078 = ~n44302 & ~n45077;
  assign n45079 = ~n44310 & ~n45078;
  assign n45080 = n45067 & ~n45079;
  assign n45081 = ~n45075 & ~n45079;
  assign n45082 = ~n45076 & ~n45080;
  assign n45083 = ~n45081 & n45082;
  assign n45084 = n45066 & ~n45083;
  assign n45085 = ~n44848 & n44856;
  assign n45086 = ~n44857 & ~n45085;
  assign n45087 = n44869 & ~n45086;
  assign n45088 = ~n44848 & ~n44856;
  assign n45089 = ~n44869 & n45088;
  assign n45090 = n44856 & n44870;
  assign n45091 = ~n45087 & ~n45089;
  assign n45092 = ~n45090 & n45091;
  assign n45093 = ~n45066 & n45083;
  assign n45094 = n45092 & ~n45093;
  assign n45095 = ~n45084 & ~n45094;
  assign n45096 = n45065 & ~n45095;
  assign n45097 = ~n44844 & n44845;
  assign n45098 = n44844 & ~n44845;
  assign n45099 = ~n45097 & ~n45098;
  assign n45100 = n44873 & ~n45099;
  assign n45101 = ~n44846 & ~n44847;
  assign n45102 = ~n44873 & ~n45101;
  assign n45103 = ~n45100 & ~n45102;
  assign n45104 = n45065 & ~n45103;
  assign n45105 = ~n45095 & ~n45103;
  assign n45106 = ~n45096 & ~n45104;
  assign n45107 = ~n45105 & n45106;
  assign n45108 = ~n45064 & ~n45107;
  assign n45109 = ~n45063 & ~n45108;
  assign n45110 = n45053 & ~n45109;
  assign n45111 = ~n44824 & n44825;
  assign n45112 = n44824 & ~n44825;
  assign n45113 = ~n45111 & ~n45112;
  assign n45114 = n44879 & ~n45113;
  assign n45115 = ~n44826 & ~n44827;
  assign n45116 = ~n44879 & ~n45115;
  assign n45117 = ~n45114 & ~n45116;
  assign n45118 = n45053 & ~n45117;
  assign n45119 = ~n45109 & ~n45117;
  assign n45120 = ~n45110 & ~n45118;
  assign n45121 = ~n45119 & n45120;
  assign n45122 = ~n45052 & ~n45121;
  assign n45123 = ~n45051 & ~n45122;
  assign n45124 = n45041 & ~n45123;
  assign n45125 = ~n44804 & n44805;
  assign n45126 = n44804 & ~n44805;
  assign n45127 = ~n45125 & ~n45126;
  assign n45128 = n44885 & ~n45127;
  assign n45129 = ~n44806 & ~n44807;
  assign n45130 = ~n44885 & ~n45129;
  assign n45131 = ~n45128 & ~n45130;
  assign n45132 = n45041 & ~n45131;
  assign n45133 = ~n45123 & ~n45131;
  assign n45134 = ~n45124 & ~n45132;
  assign n45135 = ~n45133 & n45134;
  assign n45136 = ~n45040 & ~n45135;
  assign n45137 = ~n45039 & ~n45136;
  assign n45138 = n45029 & ~n45137;
  assign n45139 = ~n44794 & ~n44795;
  assign n45140 = n44896 & n45139;
  assign n45141 = ~n44896 & ~n45139;
  assign n45142 = ~n45140 & ~n45141;
  assign n45143 = n45029 & ~n45142;
  assign n45144 = ~n45137 & ~n45142;
  assign n45145 = ~n45138 & ~n45143;
  assign n45146 = ~n45144 & n45145;
  assign n45147 = ~n45028 & ~n45146;
  assign n45148 = ~n45027 & ~n45147;
  assign n45149 = n44389 & ~n45148;
  assign n45150 = ~n44389 & n45148;
  assign n45151 = ~n45149 & ~n45150;
  assign n45152 = P4_DATAO_REG_6_ & n44390;
  assign n45153 = n44393 & ~n45023;
  assign n45154 = ~n44393 & n45023;
  assign n45155 = ~n44898 & ~n45154;
  assign n45156 = ~n45153 & ~n45155;
  assign n45157 = n45152 & ~n45156;
  assign n45158 = ~n45152 & n45156;
  assign n45159 = ~n44905 & n44906;
  assign n45160 = ~n44905 & n45014;
  assign n45161 = ~n45019 & ~n45159;
  assign n45162 = ~n45160 & n45161;
  assign n45163 = P4_DATAO_REG_7_ & n44392;
  assign n45164 = ~n44908 & n45004;
  assign n45165 = ~n45005 & ~n45011;
  assign n45166 = ~n45164 & n45165;
  assign n45167 = n44394 & ~n45166;
  assign n45168 = ~n44394 & n45166;
  assign n45169 = P4_DATAO_REG_8_ & ~n45167;
  assign n45170 = ~n45168 & n45169;
  assign n45171 = ~n44910 & ~n45001;
  assign n45172 = ~n44919 & ~n44991;
  assign n45173 = ~n44992 & ~n44998;
  assign n45174 = ~n45172 & n45173;
  assign n45175 = P4_DATAO_REG_10_ & n44623;
  assign n45176 = ~n44927 & ~n44972;
  assign n45177 = ~n44973 & ~n44979;
  assign n45178 = ~n45176 & n45177;
  assign n45179 = P4_DATAO_REG_12_ & n44102;
  assign n45180 = ~n44932 & ~n44969;
  assign n45181 = ~n44968 & ~n45180;
  assign n45182 = P4_DATAO_REG_13_ & n44104;
  assign n45183 = P4_DATAO_REG_15_ & n44106;
  assign n45184 = ~n44941 & ~n44949;
  assign n45185 = ~n44950 & ~n45184;
  assign n45186 = n45183 & ~n45185;
  assign n45187 = ~n45183 & n45185;
  assign n45188 = ~n45186 & ~n45187;
  assign n45189 = P4_DATAO_REG_16_ & n44108;
  assign n45190 = P4_DATAO_REG_17_ & n44110;
  assign n45191 = P4_DATAO_REG_18_ & n44112;
  assign n45192 = n45190 & ~n45191;
  assign n45193 = ~n45190 & n45191;
  assign n45194 = ~n45192 & ~n45193;
  assign n45195 = n45189 & ~n45194;
  assign n45196 = ~n45189 & n45194;
  assign n45197 = P4_DATAO_REG_16_ & P4_DATAO_REG_17_;
  assign n45198 = n44119 & n45197;
  assign n45199 = ~n45195 & ~n45196;
  assign n45200 = ~n45198 & n45199;
  assign n45201 = ~n45189 & ~n45192;
  assign n45202 = ~n45195 & ~n45201;
  assign n45203 = n45198 & ~n45202;
  assign n45204 = ~n45200 & ~n45203;
  assign n45205 = ~n45188 & n45204;
  assign n45206 = n45188 & ~n45204;
  assign n45207 = ~n45205 & ~n45206;
  assign n45208 = P4_DATAO_REG_14_ & n44143;
  assign n45209 = ~n45207 & ~n45208;
  assign n45210 = n45207 & n45208;
  assign n45211 = ~n44935 & ~n44953;
  assign n45212 = ~n44954 & ~n44960;
  assign n45213 = ~n45211 & n45212;
  assign n45214 = ~n45209 & ~n45210;
  assign n45215 = n45213 & n45214;
  assign n45216 = ~n45213 & ~n45214;
  assign n45217 = ~n45215 & ~n45216;
  assign n45218 = n45182 & ~n45217;
  assign n45219 = ~n45182 & n45217;
  assign n45220 = ~n45218 & ~n45219;
  assign n45221 = n45181 & ~n45220;
  assign n45222 = ~n45182 & ~n45217;
  assign n45223 = ~n45181 & n45222;
  assign n45224 = ~n45181 & n45182;
  assign n45225 = n45217 & n45224;
  assign n45226 = ~n45221 & ~n45223;
  assign n45227 = ~n45225 & n45226;
  assign n45228 = n45179 & ~n45227;
  assign n45229 = ~n45179 & n45227;
  assign n45230 = ~n45228 & ~n45229;
  assign n45231 = n45178 & ~n45230;
  assign n45232 = n45179 & n45227;
  assign n45233 = ~n45179 & ~n45227;
  assign n45234 = ~n45232 & ~n45233;
  assign n45235 = ~n45178 & ~n45234;
  assign n45236 = ~n45231 & ~n45235;
  assign n45237 = P4_DATAO_REG_11_ & n44356;
  assign n45238 = ~n44924 & ~n44988;
  assign n45239 = ~n44987 & ~n45238;
  assign n45240 = ~n45236 & ~n45237;
  assign n45241 = ~n45239 & n45240;
  assign n45242 = ~n45236 & n45237;
  assign n45243 = n45236 & ~n45237;
  assign n45244 = ~n45242 & ~n45243;
  assign n45245 = n45239 & ~n45244;
  assign n45246 = ~n45241 & ~n45245;
  assign n45247 = n45237 & ~n45239;
  assign n45248 = n45236 & n45247;
  assign n45249 = n45246 & ~n45248;
  assign n45250 = n45175 & ~n45249;
  assign n45251 = ~n45175 & n45249;
  assign n45252 = ~n45250 & ~n45251;
  assign n45253 = n45174 & ~n45252;
  assign n45254 = n45175 & n45249;
  assign n45255 = ~n45175 & ~n45249;
  assign n45256 = ~n45254 & ~n45255;
  assign n45257 = ~n45174 & ~n45256;
  assign n45258 = ~n45253 & ~n45257;
  assign n45259 = P4_DATAO_REG_9_ & n44704;
  assign n45260 = n45258 & ~n45259;
  assign n45261 = n44914 & ~n45001;
  assign n45262 = ~n44916 & ~n45261;
  assign n45263 = ~n45171 & ~n45260;
  assign n45264 = n45262 & n45263;
  assign n45265 = ~n45258 & n45259;
  assign n45266 = n45264 & ~n45265;
  assign n45267 = ~n45258 & ~n45259;
  assign n45268 = n45258 & n45259;
  assign n45269 = n44910 & n45001;
  assign n45270 = ~n44914 & ~n45171;
  assign n45271 = ~n45269 & ~n45270;
  assign n45272 = ~n45267 & ~n45268;
  assign n45273 = n45271 & n45272;
  assign n45274 = ~n45266 & ~n45273;
  assign n45275 = n45170 & ~n45274;
  assign n45276 = ~n45170 & n45274;
  assign n45277 = ~n45275 & ~n45276;
  assign n45278 = n45163 & ~n45277;
  assign n45279 = ~n45163 & n45277;
  assign n45280 = ~n45278 & ~n45279;
  assign n45281 = n45162 & ~n45280;
  assign n45282 = ~n45163 & ~n45277;
  assign n45283 = ~n45162 & n45282;
  assign n45284 = ~n45162 & n45163;
  assign n45285 = n45277 & n45284;
  assign n45286 = ~n45281 & ~n45283;
  assign n45287 = ~n45285 & n45286;
  assign n45288 = ~n45157 & ~n45158;
  assign n45289 = ~n45287 & n45288;
  assign n45290 = n45287 & ~n45288;
  assign n45291 = ~n45289 & ~n45290;
  assign n45292 = ~n45151 & n45291;
  assign n45293 = n45151 & ~n45291;
  assign n45294 = ~n45292 & ~n45293;
  assign n45295 = n44387 & n45294;
  assign n45296 = ~n44387 & ~n45294;
  assign n45297 = P4_DATAO_REG_4_ & n44388;
  assign n45298 = P4_DATAO_REG_4_ & n44390;
  assign n45299 = P4_DATAO_REG_4_ & n44392;
  assign n45300 = ~n45037 & n45038;
  assign n45301 = n45037 & ~n45038;
  assign n45302 = ~n45300 & ~n45301;
  assign n45303 = n45135 & ~n45302;
  assign n45304 = ~n45039 & ~n45040;
  assign n45305 = ~n45135 & ~n45304;
  assign n45306 = ~n45303 & ~n45305;
  assign n45307 = n45299 & ~n45306;
  assign n45308 = ~n45041 & n45131;
  assign n45309 = ~n45132 & ~n45308;
  assign n45310 = n45123 & ~n45309;
  assign n45311 = ~n45041 & ~n45131;
  assign n45312 = ~n45123 & n45311;
  assign n45313 = n45124 & n45131;
  assign n45314 = ~n45310 & ~n45312;
  assign n45315 = ~n45313 & n45314;
  assign n45316 = P4_DATAO_REG_4_ & n44394;
  assign n45317 = n45315 & n45316;
  assign n45318 = ~n45315 & ~n45316;
  assign n45319 = P4_DATAO_REG_4_ & n44704;
  assign n45320 = ~n45053 & n45117;
  assign n45321 = ~n45118 & ~n45320;
  assign n45322 = n45109 & ~n45321;
  assign n45323 = ~n45053 & ~n45117;
  assign n45324 = ~n45109 & n45323;
  assign n45325 = n45110 & n45117;
  assign n45326 = ~n45322 & ~n45324;
  assign n45327 = ~n45325 & n45326;
  assign n45328 = P4_DATAO_REG_4_ & n44623;
  assign n45329 = n45327 & n45328;
  assign n45330 = ~n45327 & ~n45328;
  assign n45331 = P4_DATAO_REG_4_ & n44356;
  assign n45332 = ~n45065 & n45103;
  assign n45333 = ~n45104 & ~n45332;
  assign n45334 = n45095 & ~n45333;
  assign n45335 = ~n45065 & ~n45103;
  assign n45336 = ~n45095 & n45335;
  assign n45337 = n45096 & n45103;
  assign n45338 = ~n45334 & ~n45336;
  assign n45339 = ~n45337 & n45338;
  assign n45340 = P4_DATAO_REG_4_ & n44102;
  assign n45341 = n45339 & n45340;
  assign n45342 = ~n45339 & ~n45340;
  assign n45343 = P4_DATAO_REG_4_ & n44104;
  assign n45344 = n45066 & ~n45092;
  assign n45345 = ~n45066 & n45092;
  assign n45346 = ~n45344 & ~n45345;
  assign n45347 = n45083 & ~n45346;
  assign n45348 = ~n45066 & ~n45092;
  assign n45349 = ~n45083 & n45348;
  assign n45350 = n45084 & n45092;
  assign n45351 = ~n45347 & ~n45349;
  assign n45352 = ~n45350 & n45351;
  assign n45353 = n45343 & ~n45352;
  assign n45354 = P4_DATAO_REG_4_ & n44143;
  assign n45355 = ~n44295 & ~n44313;
  assign n45356 = ~n44314 & ~n44320;
  assign n45357 = ~n45355 & n45356;
  assign n45358 = n45354 & ~n45357;
  assign n45359 = ~n45067 & n45075;
  assign n45360 = ~n45076 & ~n45359;
  assign n45361 = n45079 & ~n45360;
  assign n45362 = ~n45067 & ~n45075;
  assign n45363 = ~n45079 & n45362;
  assign n45364 = n45075 & n45080;
  assign n45365 = ~n45361 & ~n45363;
  assign n45366 = ~n45364 & n45365;
  assign n45367 = ~n45354 & n45357;
  assign n45368 = n45366 & ~n45367;
  assign n45369 = ~n45358 & ~n45368;
  assign n45370 = n45343 & ~n45369;
  assign n45371 = ~n45352 & ~n45369;
  assign n45372 = ~n45353 & ~n45370;
  assign n45373 = ~n45371 & n45372;
  assign n45374 = ~n45342 & ~n45373;
  assign n45375 = ~n45341 & ~n45374;
  assign n45376 = n45331 & ~n45375;
  assign n45377 = ~n45061 & n45062;
  assign n45378 = n45061 & ~n45062;
  assign n45379 = ~n45377 & ~n45378;
  assign n45380 = n45107 & ~n45379;
  assign n45381 = ~n45063 & ~n45064;
  assign n45382 = ~n45107 & ~n45381;
  assign n45383 = ~n45380 & ~n45382;
  assign n45384 = n45331 & ~n45383;
  assign n45385 = ~n45375 & ~n45383;
  assign n45386 = ~n45376 & ~n45384;
  assign n45387 = ~n45385 & n45386;
  assign n45388 = ~n45330 & ~n45387;
  assign n45389 = ~n45329 & ~n45388;
  assign n45390 = n45319 & ~n45389;
  assign n45391 = ~n45049 & n45050;
  assign n45392 = n45049 & ~n45050;
  assign n45393 = ~n45391 & ~n45392;
  assign n45394 = n45121 & ~n45393;
  assign n45395 = ~n45051 & ~n45052;
  assign n45396 = ~n45121 & ~n45395;
  assign n45397 = ~n45394 & ~n45396;
  assign n45398 = n45319 & ~n45397;
  assign n45399 = ~n45389 & ~n45397;
  assign n45400 = ~n45390 & ~n45398;
  assign n45401 = ~n45399 & n45400;
  assign n45402 = ~n45318 & ~n45401;
  assign n45403 = ~n45317 & ~n45402;
  assign n45404 = n45299 & ~n45403;
  assign n45405 = ~n45306 & ~n45403;
  assign n45406 = ~n45307 & ~n45404;
  assign n45407 = ~n45405 & n45406;
  assign n45408 = n45298 & ~n45407;
  assign n45409 = ~n45029 & n45142;
  assign n45410 = ~n45143 & ~n45409;
  assign n45411 = n45137 & ~n45410;
  assign n45412 = ~n45029 & ~n45142;
  assign n45413 = ~n45137 & n45412;
  assign n45414 = n45138 & n45142;
  assign n45415 = ~n45411 & ~n45413;
  assign n45416 = ~n45414 & n45415;
  assign n45417 = ~n45298 & n45407;
  assign n45418 = n45416 & ~n45417;
  assign n45419 = ~n45408 & ~n45418;
  assign n45420 = n45297 & ~n45419;
  assign n45421 = ~n45027 & ~n45028;
  assign n45422 = n45146 & n45421;
  assign n45423 = ~n45146 & ~n45421;
  assign n45424 = ~n45422 & ~n45423;
  assign n45425 = n45297 & ~n45424;
  assign n45426 = ~n45419 & ~n45424;
  assign n45427 = ~n45420 & ~n45425;
  assign n45428 = ~n45426 & n45427;
  assign n45429 = ~n45296 & ~n45428;
  assign n45430 = ~n45295 & ~n45429;
  assign n45431 = n44385 & ~n45430;
  assign n45432 = ~n44385 & n45430;
  assign n45433 = ~n45431 & ~n45432;
  assign n45434 = n44389 & ~n45291;
  assign n45435 = ~n44389 & n45291;
  assign n45436 = ~n45148 & ~n45435;
  assign n45437 = ~n45434 & ~n45436;
  assign n45438 = P4_DATAO_REG_5_ & n44386;
  assign n45439 = ~n45158 & n45287;
  assign n45440 = ~n45157 & ~n45439;
  assign n45441 = P4_DATAO_REG_6_ & n44388;
  assign n45442 = ~n45162 & ~n45277;
  assign n45443 = ~n45278 & ~n45284;
  assign n45444 = ~n45442 & n45443;
  assign n45445 = P4_DATAO_REG_7_ & n44390;
  assign n45446 = P4_DATAO_REG_8_ & ~n45168;
  assign n45447 = n45274 & n45446;
  assign n45448 = ~n45167 & ~n45447;
  assign n45449 = P4_DATAO_REG_8_ & n44392;
  assign n45450 = P4_DATAO_REG_10_ & n44704;
  assign n45451 = ~n45174 & ~n45255;
  assign n45452 = ~n45254 & ~n45451;
  assign n45453 = n45450 & ~n45452;
  assign n45454 = ~n45450 & n45452;
  assign n45455 = ~n45453 & ~n45454;
  assign n45456 = P4_DATAO_REG_11_ & n44623;
  assign n45457 = ~n45236 & ~n45239;
  assign n45458 = ~n45242 & ~n45247;
  assign n45459 = ~n45457 & n45458;
  assign n45460 = n45456 & ~n45459;
  assign n45461 = ~n45456 & n45459;
  assign n45462 = ~n45460 & ~n45461;
  assign n45463 = ~n45178 & ~n45233;
  assign n45464 = ~n45232 & ~n45463;
  assign n45465 = P4_DATAO_REG_12_ & n44356;
  assign n45466 = ~n45181 & ~n45217;
  assign n45467 = ~n45218 & ~n45224;
  assign n45468 = ~n45466 & n45467;
  assign n45469 = P4_DATAO_REG_13_ & n44102;
  assign n45470 = n45183 & ~n45204;
  assign n45471 = ~n45183 & n45204;
  assign n45472 = ~n45185 & ~n45471;
  assign n45473 = ~n45470 & ~n45472;
  assign n45474 = P4_DATAO_REG_15_ & n44143;
  assign n45475 = P4_DATAO_REG_17_ & n44108;
  assign n45476 = P4_DATAO_REG_18_ & n44110;
  assign n45477 = P4_DATAO_REG_19_ & n44112;
  assign n45478 = n45476 & ~n45477;
  assign n45479 = ~n45476 & n45477;
  assign n45480 = ~n45478 & ~n45479;
  assign n45481 = n45475 & ~n45480;
  assign n45482 = ~n45475 & n45480;
  assign n45483 = P4_DATAO_REG_17_ & P4_DATAO_REG_18_;
  assign n45484 = n44119 & n45483;
  assign n45485 = ~n45481 & ~n45482;
  assign n45486 = ~n45484 & n45485;
  assign n45487 = n45475 & ~n45478;
  assign n45488 = ~n45475 & n45478;
  assign n45489 = ~n45487 & ~n45488;
  assign n45490 = n45484 & n45489;
  assign n45491 = ~n45486 & ~n45490;
  assign n45492 = P4_DATAO_REG_16_ & n44106;
  assign n45493 = ~n45196 & n45198;
  assign n45494 = ~n45195 & ~n45493;
  assign n45495 = ~n45491 & ~n45492;
  assign n45496 = ~n45494 & n45495;
  assign n45497 = n45491 & n45492;
  assign n45498 = ~n45495 & ~n45497;
  assign n45499 = n45494 & n45498;
  assign n45500 = ~n45496 & ~n45499;
  assign n45501 = n45492 & ~n45494;
  assign n45502 = n45491 & n45501;
  assign n45503 = n45500 & ~n45502;
  assign n45504 = n45474 & ~n45503;
  assign n45505 = ~n45474 & n45503;
  assign n45506 = ~n45504 & ~n45505;
  assign n45507 = n45473 & ~n45506;
  assign n45508 = n45474 & n45500;
  assign n45509 = ~n45502 & n45508;
  assign n45510 = ~n45474 & ~n45503;
  assign n45511 = ~n45509 & ~n45510;
  assign n45512 = ~n45473 & ~n45511;
  assign n45513 = ~n45507 & ~n45512;
  assign n45514 = P4_DATAO_REG_14_ & n44104;
  assign n45515 = ~n45209 & ~n45213;
  assign n45516 = ~n45210 & ~n45515;
  assign n45517 = ~n45513 & ~n45514;
  assign n45518 = ~n45516 & n45517;
  assign n45519 = ~n45513 & n45514;
  assign n45520 = n45513 & ~n45514;
  assign n45521 = ~n45519 & ~n45520;
  assign n45522 = n45516 & ~n45521;
  assign n45523 = ~n45518 & ~n45522;
  assign n45524 = n45514 & ~n45516;
  assign n45525 = n45513 & n45524;
  assign n45526 = n45523 & ~n45525;
  assign n45527 = n45469 & ~n45526;
  assign n45528 = ~n45469 & n45526;
  assign n45529 = ~n45527 & ~n45528;
  assign n45530 = n45468 & ~n45529;
  assign n45531 = n45469 & ~n45525;
  assign n45532 = n45523 & n45531;
  assign n45533 = ~n45469 & ~n45526;
  assign n45534 = ~n45532 & ~n45533;
  assign n45535 = ~n45468 & ~n45534;
  assign n45536 = ~n45530 & ~n45535;
  assign n45537 = n45465 & ~n45536;
  assign n45538 = ~n45465 & n45536;
  assign n45539 = ~n45537 & ~n45538;
  assign n45540 = n45464 & ~n45539;
  assign n45541 = ~n45465 & ~n45536;
  assign n45542 = ~n45464 & n45541;
  assign n45543 = ~n45464 & n45465;
  assign n45544 = n45536 & n45543;
  assign n45545 = ~n45540 & ~n45542;
  assign n45546 = ~n45544 & n45545;
  assign n45547 = n45462 & ~n45546;
  assign n45548 = ~n45462 & n45546;
  assign n45549 = ~n45547 & ~n45548;
  assign n45550 = ~n45455 & n45549;
  assign n45551 = n45455 & ~n45549;
  assign n45552 = ~n45550 & ~n45551;
  assign n45553 = P4_DATAO_REG_9_ & n44394;
  assign n45554 = n45552 & n45553;
  assign n45555 = ~n45552 & ~n45553;
  assign n45556 = ~n45554 & ~n45555;
  assign n45557 = ~n45264 & ~n45265;
  assign n45558 = ~n45556 & ~n45557;
  assign n45559 = n45556 & n45557;
  assign n45560 = ~n45558 & ~n45559;
  assign n45561 = n45449 & ~n45560;
  assign n45562 = ~n45449 & n45560;
  assign n45563 = ~n45561 & ~n45562;
  assign n45564 = n45448 & ~n45563;
  assign n45565 = ~n45449 & ~n45560;
  assign n45566 = ~n45448 & n45565;
  assign n45567 = ~n45448 & n45449;
  assign n45568 = n45560 & n45567;
  assign n45569 = ~n45564 & ~n45566;
  assign n45570 = ~n45568 & n45569;
  assign n45571 = n45445 & ~n45570;
  assign n45572 = ~n45445 & n45570;
  assign n45573 = ~n45571 & ~n45572;
  assign n45574 = n45444 & ~n45573;
  assign n45575 = n45445 & n45570;
  assign n45576 = ~n45445 & ~n45570;
  assign n45577 = ~n45575 & ~n45576;
  assign n45578 = ~n45444 & ~n45577;
  assign n45579 = ~n45574 & ~n45578;
  assign n45580 = n45441 & ~n45579;
  assign n45581 = ~n45441 & n45579;
  assign n45582 = ~n45580 & ~n45581;
  assign n45583 = n45440 & ~n45582;
  assign n45584 = ~n45441 & ~n45579;
  assign n45585 = ~n45440 & n45584;
  assign n45586 = ~n45440 & n45441;
  assign n45587 = n45579 & n45586;
  assign n45588 = ~n45583 & ~n45585;
  assign n45589 = ~n45587 & n45588;
  assign n45590 = n45438 & ~n45589;
  assign n45591 = ~n45438 & n45589;
  assign n45592 = ~n45590 & ~n45591;
  assign n45593 = n45437 & ~n45592;
  assign n45594 = n45438 & n45589;
  assign n45595 = ~n45438 & ~n45589;
  assign n45596 = ~n45594 & ~n45595;
  assign n45597 = ~n45437 & ~n45596;
  assign n45598 = ~n45593 & ~n45597;
  assign n45599 = ~n45433 & n45598;
  assign n45600 = n45433 & ~n45598;
  assign n45601 = ~n45599 & ~n45600;
  assign n45602 = SEL & DIN_16_;
  assign n45603 = P4_DATAO_REG_3_ & n45602;
  assign n45604 = ~n45601 & ~n45603;
  assign n45605 = n45601 & n45603;
  assign n45606 = P4_DATAO_REG_3_ & n44384;
  assign n45607 = ~n45295 & ~n45296;
  assign n45608 = ~n45428 & ~n45607;
  assign n45609 = n45428 & n45607;
  assign n45610 = ~n45608 & ~n45609;
  assign n45611 = n45606 & ~n45610;
  assign n45612 = ~n45606 & n45610;
  assign n45613 = ~n45297 & n45424;
  assign n45614 = ~n45425 & ~n45613;
  assign n45615 = n45419 & ~n45614;
  assign n45616 = ~n45297 & ~n45424;
  assign n45617 = ~n45419 & n45616;
  assign n45618 = n45420 & n45424;
  assign n45619 = ~n45615 & ~n45617;
  assign n45620 = ~n45618 & n45619;
  assign n45621 = P4_DATAO_REG_3_ & n44386;
  assign n45622 = n45620 & n45621;
  assign n45623 = ~n45620 & ~n45621;
  assign n45624 = P4_DATAO_REG_3_ & n44388;
  assign n45625 = ~n45299 & n45403;
  assign n45626 = ~n45404 & ~n45625;
  assign n45627 = n45306 & ~n45626;
  assign n45628 = ~n45299 & ~n45403;
  assign n45629 = ~n45306 & n45628;
  assign n45630 = n45307 & n45403;
  assign n45631 = ~n45627 & ~n45629;
  assign n45632 = ~n45630 & n45631;
  assign n45633 = P4_DATAO_REG_3_ & n44390;
  assign n45634 = n45632 & n45633;
  assign n45635 = ~n45632 & ~n45633;
  assign n45636 = P4_DATAO_REG_3_ & n44392;
  assign n45637 = ~n45319 & n45397;
  assign n45638 = ~n45398 & ~n45637;
  assign n45639 = n45389 & ~n45638;
  assign n45640 = ~n45319 & ~n45397;
  assign n45641 = ~n45389 & n45640;
  assign n45642 = n45390 & n45397;
  assign n45643 = ~n45639 & ~n45641;
  assign n45644 = ~n45642 & n45643;
  assign n45645 = P4_DATAO_REG_3_ & n44394;
  assign n45646 = n45644 & n45645;
  assign n45647 = ~n45644 & ~n45645;
  assign n45648 = P4_DATAO_REG_3_ & n44704;
  assign n45649 = ~n45331 & n45383;
  assign n45650 = ~n45384 & ~n45649;
  assign n45651 = n45375 & ~n45650;
  assign n45652 = ~n45331 & ~n45383;
  assign n45653 = ~n45375 & n45652;
  assign n45654 = n45376 & n45383;
  assign n45655 = ~n45651 & ~n45653;
  assign n45656 = ~n45654 & n45655;
  assign n45657 = P4_DATAO_REG_3_ & n44623;
  assign n45658 = n45656 & n45657;
  assign n45659 = ~n45656 & ~n45657;
  assign n45660 = P4_DATAO_REG_3_ & n44356;
  assign n45661 = P4_DATAO_REG_3_ & n44102;
  assign n45662 = P4_DATAO_REG_3_ & n44104;
  assign n45663 = n45354 & ~n45366;
  assign n45664 = ~n45354 & n45366;
  assign n45665 = ~n45663 & ~n45664;
  assign n45666 = n45357 & ~n45665;
  assign n45667 = ~n45354 & ~n45366;
  assign n45668 = ~n45357 & n45667;
  assign n45669 = n45358 & n45366;
  assign n45670 = ~n45666 & ~n45668;
  assign n45671 = ~n45669 & n45670;
  assign n45672 = n45662 & ~n45671;
  assign n45673 = ~n44292 & n44329;
  assign n45674 = n44323 & ~n45673;
  assign n45675 = ~n44333 & ~n45674;
  assign n45676 = n45662 & ~n45675;
  assign n45677 = ~n45671 & ~n45675;
  assign n45678 = ~n45672 & ~n45676;
  assign n45679 = ~n45677 & n45678;
  assign n45680 = n45661 & ~n45679;
  assign n45681 = ~n45343 & n45352;
  assign n45682 = ~n45353 & ~n45681;
  assign n45683 = n45369 & ~n45682;
  assign n45684 = ~n45343 & ~n45352;
  assign n45685 = ~n45369 & n45684;
  assign n45686 = n45352 & n45370;
  assign n45687 = ~n45683 & ~n45685;
  assign n45688 = ~n45686 & n45687;
  assign n45689 = ~n45661 & n45679;
  assign n45690 = n45688 & ~n45689;
  assign n45691 = ~n45680 & ~n45690;
  assign n45692 = n45660 & ~n45691;
  assign n45693 = ~n45339 & n45340;
  assign n45694 = n45339 & ~n45340;
  assign n45695 = ~n45693 & ~n45694;
  assign n45696 = n45373 & ~n45695;
  assign n45697 = ~n45341 & ~n45342;
  assign n45698 = ~n45373 & ~n45697;
  assign n45699 = ~n45696 & ~n45698;
  assign n45700 = n45660 & ~n45699;
  assign n45701 = ~n45691 & ~n45699;
  assign n45702 = ~n45692 & ~n45700;
  assign n45703 = ~n45701 & n45702;
  assign n45704 = ~n45659 & ~n45703;
  assign n45705 = ~n45658 & ~n45704;
  assign n45706 = n45648 & ~n45705;
  assign n45707 = ~n45327 & n45328;
  assign n45708 = n45327 & ~n45328;
  assign n45709 = ~n45707 & ~n45708;
  assign n45710 = n45387 & ~n45709;
  assign n45711 = ~n45329 & ~n45330;
  assign n45712 = ~n45387 & ~n45711;
  assign n45713 = ~n45710 & ~n45712;
  assign n45714 = n45648 & ~n45713;
  assign n45715 = ~n45705 & ~n45713;
  assign n45716 = ~n45706 & ~n45714;
  assign n45717 = ~n45715 & n45716;
  assign n45718 = ~n45647 & ~n45717;
  assign n45719 = ~n45646 & ~n45718;
  assign n45720 = n45636 & ~n45719;
  assign n45721 = ~n45315 & n45316;
  assign n45722 = n45315 & ~n45316;
  assign n45723 = ~n45721 & ~n45722;
  assign n45724 = n45401 & ~n45723;
  assign n45725 = ~n45317 & ~n45318;
  assign n45726 = ~n45401 & ~n45725;
  assign n45727 = ~n45724 & ~n45726;
  assign n45728 = n45636 & ~n45727;
  assign n45729 = ~n45719 & ~n45727;
  assign n45730 = ~n45720 & ~n45728;
  assign n45731 = ~n45729 & n45730;
  assign n45732 = ~n45635 & ~n45731;
  assign n45733 = ~n45634 & ~n45732;
  assign n45734 = n45624 & ~n45733;
  assign n45735 = ~n45408 & ~n45417;
  assign n45736 = ~n45416 & n45735;
  assign n45737 = n45416 & ~n45735;
  assign n45738 = ~n45736 & ~n45737;
  assign n45739 = n45624 & ~n45738;
  assign n45740 = ~n45733 & ~n45738;
  assign n45741 = ~n45734 & ~n45739;
  assign n45742 = ~n45740 & n45741;
  assign n45743 = ~n45623 & ~n45742;
  assign n45744 = ~n45622 & ~n45743;
  assign n45745 = ~n45612 & ~n45744;
  assign n45746 = ~n45611 & ~n45745;
  assign n45747 = ~n45604 & ~n45605;
  assign n45748 = n45746 & n45747;
  assign n45749 = ~n45746 & ~n45747;
  assign n45750 = ~n45748 & ~n45749;
  assign n45751 = n44383 & ~n45750;
  assign n45752 = ~n44383 & n45750;
  assign n45753 = P4_DATAO_REG_2_ & n45602;
  assign n45754 = n45606 & n45610;
  assign n45755 = ~n45606 & ~n45610;
  assign n45756 = ~n45754 & ~n45755;
  assign n45757 = ~n45744 & ~n45756;
  assign n45758 = n45744 & n45756;
  assign n45759 = ~n45757 & ~n45758;
  assign n45760 = n45753 & n45759;
  assign n45761 = ~n45753 & ~n45759;
  assign n45762 = P4_DATAO_REG_2_ & n44384;
  assign n45763 = ~n45620 & n45621;
  assign n45764 = n45620 & ~n45621;
  assign n45765 = ~n45763 & ~n45764;
  assign n45766 = n45742 & ~n45765;
  assign n45767 = ~n45622 & ~n45623;
  assign n45768 = ~n45742 & ~n45767;
  assign n45769 = ~n45766 & ~n45768;
  assign n45770 = n45762 & ~n45769;
  assign n45771 = ~n45624 & n45738;
  assign n45772 = ~n45739 & ~n45771;
  assign n45773 = n45733 & ~n45772;
  assign n45774 = ~n45624 & ~n45738;
  assign n45775 = ~n45733 & n45774;
  assign n45776 = n45734 & n45738;
  assign n45777 = ~n45773 & ~n45775;
  assign n45778 = ~n45776 & n45777;
  assign n45779 = P4_DATAO_REG_2_ & n44386;
  assign n45780 = n45778 & n45779;
  assign n45781 = ~n45778 & ~n45779;
  assign n45782 = P4_DATAO_REG_2_ & n44388;
  assign n45783 = ~n45636 & n45727;
  assign n45784 = ~n45728 & ~n45783;
  assign n45785 = n45719 & ~n45784;
  assign n45786 = ~n45636 & ~n45727;
  assign n45787 = ~n45719 & n45786;
  assign n45788 = n45720 & n45727;
  assign n45789 = ~n45785 & ~n45787;
  assign n45790 = ~n45788 & n45789;
  assign n45791 = P4_DATAO_REG_2_ & n44390;
  assign n45792 = n45790 & n45791;
  assign n45793 = ~n45790 & ~n45791;
  assign n45794 = P4_DATAO_REG_2_ & n44392;
  assign n45795 = ~n45648 & n45713;
  assign n45796 = ~n45714 & ~n45795;
  assign n45797 = n45705 & ~n45796;
  assign n45798 = ~n45648 & ~n45713;
  assign n45799 = ~n45705 & n45798;
  assign n45800 = n45706 & n45713;
  assign n45801 = ~n45797 & ~n45799;
  assign n45802 = ~n45800 & n45801;
  assign n45803 = P4_DATAO_REG_2_ & n44394;
  assign n45804 = n45802 & n45803;
  assign n45805 = ~n45802 & ~n45803;
  assign n45806 = P4_DATAO_REG_2_ & n44704;
  assign n45807 = ~n45660 & n45699;
  assign n45808 = ~n45700 & ~n45807;
  assign n45809 = n45691 & ~n45808;
  assign n45810 = ~n45660 & ~n45699;
  assign n45811 = ~n45691 & n45810;
  assign n45812 = n45692 & n45699;
  assign n45813 = ~n45809 & ~n45811;
  assign n45814 = ~n45812 & n45813;
  assign n45815 = P4_DATAO_REG_2_ & n44623;
  assign n45816 = n45814 & n45815;
  assign n45817 = ~n45814 & ~n45815;
  assign n45818 = P4_DATAO_REG_2_ & n44356;
  assign n45819 = ~n45662 & n45671;
  assign n45820 = ~n45672 & ~n45819;
  assign n45821 = n45675 & ~n45820;
  assign n45822 = ~n45662 & ~n45671;
  assign n45823 = ~n45675 & n45822;
  assign n45824 = n45671 & n45676;
  assign n45825 = ~n45821 & ~n45823;
  assign n45826 = ~n45824 & n45825;
  assign n45827 = P4_DATAO_REG_2_ & n44102;
  assign n45828 = n45826 & n45827;
  assign n45829 = ~n45826 & ~n45827;
  assign n45830 = ~n44290 & ~n44336;
  assign n45831 = ~n44337 & ~n44343;
  assign n45832 = ~n45830 & n45831;
  assign n45833 = ~n45829 & ~n45832;
  assign n45834 = ~n45828 & ~n45833;
  assign n45835 = n45818 & ~n45834;
  assign n45836 = n45661 & ~n45688;
  assign n45837 = ~n45661 & n45688;
  assign n45838 = ~n45836 & ~n45837;
  assign n45839 = n45679 & ~n45838;
  assign n45840 = ~n45661 & ~n45688;
  assign n45841 = ~n45679 & n45840;
  assign n45842 = n45680 & n45688;
  assign n45843 = ~n45839 & ~n45841;
  assign n45844 = ~n45842 & n45843;
  assign n45845 = n45818 & ~n45844;
  assign n45846 = ~n45834 & ~n45844;
  assign n45847 = ~n45835 & ~n45845;
  assign n45848 = ~n45846 & n45847;
  assign n45849 = ~n45817 & ~n45848;
  assign n45850 = ~n45816 & ~n45849;
  assign n45851 = n45806 & ~n45850;
  assign n45852 = ~n45656 & n45657;
  assign n45853 = n45656 & ~n45657;
  assign n45854 = ~n45852 & ~n45853;
  assign n45855 = n45703 & ~n45854;
  assign n45856 = ~n45658 & ~n45659;
  assign n45857 = ~n45703 & ~n45856;
  assign n45858 = ~n45855 & ~n45857;
  assign n45859 = n45806 & ~n45858;
  assign n45860 = ~n45850 & ~n45858;
  assign n45861 = ~n45851 & ~n45859;
  assign n45862 = ~n45860 & n45861;
  assign n45863 = ~n45805 & ~n45862;
  assign n45864 = ~n45804 & ~n45863;
  assign n45865 = n45794 & ~n45864;
  assign n45866 = ~n45644 & n45645;
  assign n45867 = n45644 & ~n45645;
  assign n45868 = ~n45866 & ~n45867;
  assign n45869 = n45717 & ~n45868;
  assign n45870 = ~n45646 & ~n45647;
  assign n45871 = ~n45717 & ~n45870;
  assign n45872 = ~n45869 & ~n45871;
  assign n45873 = n45794 & ~n45872;
  assign n45874 = ~n45864 & ~n45872;
  assign n45875 = ~n45865 & ~n45873;
  assign n45876 = ~n45874 & n45875;
  assign n45877 = ~n45793 & ~n45876;
  assign n45878 = ~n45792 & ~n45877;
  assign n45879 = n45782 & ~n45878;
  assign n45880 = ~n45632 & n45633;
  assign n45881 = n45632 & ~n45633;
  assign n45882 = ~n45880 & ~n45881;
  assign n45883 = n45731 & ~n45882;
  assign n45884 = ~n45634 & ~n45635;
  assign n45885 = ~n45731 & ~n45884;
  assign n45886 = ~n45883 & ~n45885;
  assign n45887 = n45782 & ~n45886;
  assign n45888 = ~n45878 & ~n45886;
  assign n45889 = ~n45879 & ~n45887;
  assign n45890 = ~n45888 & n45889;
  assign n45891 = ~n45781 & ~n45890;
  assign n45892 = ~n45780 & ~n45891;
  assign n45893 = n45762 & ~n45892;
  assign n45894 = ~n45769 & ~n45892;
  assign n45895 = ~n45770 & ~n45893;
  assign n45896 = ~n45894 & n45895;
  assign n45897 = ~n45761 & ~n45896;
  assign n45898 = ~n45760 & ~n45897;
  assign n45899 = ~n45752 & ~n45898;
  assign n45900 = ~n45751 & ~n45899;
  assign n45901 = n44381 & ~n45900;
  assign n45902 = ~n44381 & n45900;
  assign n45903 = ~n45901 & ~n45902;
  assign n45904 = ~n45604 & ~n45746;
  assign n45905 = ~n45605 & ~n45904;
  assign n45906 = P4_DATAO_REG_3_ & n44382;
  assign n45907 = n44385 & ~n45598;
  assign n45908 = ~n44385 & n45598;
  assign n45909 = ~n45430 & ~n45908;
  assign n45910 = ~n45907 & ~n45909;
  assign n45911 = P4_DATAO_REG_4_ & n45602;
  assign n45912 = ~n45437 & ~n45595;
  assign n45913 = ~n45594 & ~n45912;
  assign n45914 = P4_DATAO_REG_5_ & n44384;
  assign n45915 = ~n45440 & ~n45579;
  assign n45916 = ~n45580 & ~n45586;
  assign n45917 = ~n45915 & n45916;
  assign n45918 = P4_DATAO_REG_6_ & n44386;
  assign n45919 = n45553 & ~n45557;
  assign n45920 = ~n45553 & n45557;
  assign n45921 = n45552 & ~n45920;
  assign n45922 = ~n45919 & ~n45921;
  assign n45923 = P4_DATAO_REG_9_ & n44392;
  assign n45924 = n45450 & ~n45549;
  assign n45925 = ~n45450 & n45549;
  assign n45926 = ~n45452 & ~n45925;
  assign n45927 = ~n45924 & ~n45926;
  assign n45928 = P4_DATAO_REG_10_ & n44394;
  assign n45929 = ~n45464 & ~n45536;
  assign n45930 = ~n45537 & ~n45543;
  assign n45931 = ~n45929 & n45930;
  assign n45932 = P4_DATAO_REG_12_ & n44623;
  assign n45933 = P4_DATAO_REG_14_ & n44102;
  assign n45934 = ~n45513 & ~n45516;
  assign n45935 = ~n45519 & ~n45524;
  assign n45936 = ~n45934 & n45935;
  assign n45937 = n45933 & ~n45936;
  assign n45938 = ~n45933 & n45936;
  assign n45939 = ~n45937 & ~n45938;
  assign n45940 = ~n45473 & ~n45510;
  assign n45941 = ~n45509 & ~n45940;
  assign n45942 = P4_DATAO_REG_15_ & n44104;
  assign n45943 = ~n45491 & n45492;
  assign n45944 = ~n45491 & ~n45494;
  assign n45945 = ~n45501 & ~n45943;
  assign n45946 = ~n45944 & n45945;
  assign n45947 = P4_DATAO_REG_16_ & n44143;
  assign n45948 = P4_DATAO_REG_18_ & n44108;
  assign n45949 = P4_DATAO_REG_19_ & n44110;
  assign n45950 = P4_DATAO_REG_20_ & n44112;
  assign n45951 = n45949 & ~n45950;
  assign n45952 = ~n45949 & n45950;
  assign n45953 = ~n45951 & ~n45952;
  assign n45954 = n45948 & ~n45953;
  assign n45955 = ~n45948 & n45953;
  assign n45956 = P4_DATAO_REG_18_ & P4_DATAO_REG_19_;
  assign n45957 = n44119 & n45956;
  assign n45958 = ~n45954 & ~n45955;
  assign n45959 = ~n45957 & n45958;
  assign n45960 = ~n45948 & ~n45951;
  assign n45961 = ~n45954 & ~n45960;
  assign n45962 = n45957 & ~n45961;
  assign n45963 = ~n45959 & ~n45962;
  assign n45964 = P4_DATAO_REG_17_ & n44106;
  assign n45965 = ~n45482 & n45484;
  assign n45966 = ~n45481 & ~n45965;
  assign n45967 = ~n45963 & ~n45964;
  assign n45968 = ~n45966 & n45967;
  assign n45969 = ~n45963 & n45964;
  assign n45970 = n45963 & ~n45964;
  assign n45971 = ~n45969 & ~n45970;
  assign n45972 = n45966 & ~n45971;
  assign n45973 = ~n45968 & ~n45972;
  assign n45974 = n45964 & ~n45966;
  assign n45975 = n45963 & n45974;
  assign n45976 = n45973 & ~n45975;
  assign n45977 = n45947 & ~n45976;
  assign n45978 = ~n45947 & n45976;
  assign n45979 = ~n45977 & ~n45978;
  assign n45980 = n45946 & ~n45979;
  assign n45981 = n45947 & ~n45975;
  assign n45982 = n45973 & n45981;
  assign n45983 = ~n45947 & ~n45976;
  assign n45984 = ~n45982 & ~n45983;
  assign n45985 = ~n45946 & ~n45984;
  assign n45986 = ~n45980 & ~n45985;
  assign n45987 = n45942 & ~n45986;
  assign n45988 = ~n45942 & n45986;
  assign n45989 = ~n45987 & ~n45988;
  assign n45990 = n45941 & ~n45989;
  assign n45991 = ~n45942 & ~n45986;
  assign n45992 = ~n45941 & n45991;
  assign n45993 = ~n45941 & n45942;
  assign n45994 = n45986 & n45993;
  assign n45995 = ~n45990 & ~n45992;
  assign n45996 = ~n45994 & n45995;
  assign n45997 = n45939 & ~n45996;
  assign n45998 = ~n45939 & n45996;
  assign n45999 = ~n45997 & ~n45998;
  assign n46000 = P4_DATAO_REG_13_ & n44356;
  assign n46001 = ~n45468 & n45469;
  assign n46002 = ~n45532 & ~n46001;
  assign n46003 = ~n45468 & n45526;
  assign n46004 = n46002 & ~n46003;
  assign n46005 = ~n45999 & ~n46000;
  assign n46006 = ~n46004 & n46005;
  assign n46007 = n45999 & n46000;
  assign n46008 = ~n46005 & ~n46007;
  assign n46009 = n46004 & n46008;
  assign n46010 = ~n46006 & ~n46009;
  assign n46011 = n46000 & ~n46004;
  assign n46012 = n45999 & n46011;
  assign n46013 = n46010 & ~n46012;
  assign n46014 = n45932 & ~n46013;
  assign n46015 = ~n45932 & n46013;
  assign n46016 = ~n46014 & ~n46015;
  assign n46017 = n45931 & ~n46016;
  assign n46018 = n45932 & ~n46012;
  assign n46019 = n46010 & n46018;
  assign n46020 = ~n45932 & ~n46013;
  assign n46021 = ~n46019 & ~n46020;
  assign n46022 = ~n45931 & ~n46021;
  assign n46023 = ~n46017 & ~n46022;
  assign n46024 = P4_DATAO_REG_11_ & n44704;
  assign n46025 = ~n45461 & n45546;
  assign n46026 = ~n45460 & ~n46025;
  assign n46027 = ~n46023 & ~n46024;
  assign n46028 = ~n46026 & n46027;
  assign n46029 = ~n46023 & n46024;
  assign n46030 = n46023 & ~n46024;
  assign n46031 = ~n46029 & ~n46030;
  assign n46032 = n46026 & ~n46031;
  assign n46033 = ~n46028 & ~n46032;
  assign n46034 = n46024 & ~n46026;
  assign n46035 = n46023 & n46034;
  assign n46036 = n46033 & ~n46035;
  assign n46037 = n45928 & ~n46036;
  assign n46038 = ~n45928 & n46036;
  assign n46039 = ~n46037 & ~n46038;
  assign n46040 = n45927 & ~n46039;
  assign n46041 = n45928 & ~n46035;
  assign n46042 = n46033 & n46041;
  assign n46043 = ~n45928 & ~n46036;
  assign n46044 = ~n46042 & ~n46043;
  assign n46045 = ~n45927 & ~n46044;
  assign n46046 = ~n46040 & ~n46045;
  assign n46047 = n45923 & ~n46046;
  assign n46048 = ~n45923 & n46046;
  assign n46049 = ~n46047 & ~n46048;
  assign n46050 = n45922 & ~n46049;
  assign n46051 = ~n45922 & n46049;
  assign n46052 = ~n46050 & ~n46051;
  assign n46053 = P4_DATAO_REG_8_ & n44390;
  assign n46054 = ~n46052 & ~n46053;
  assign n46055 = n46052 & n46053;
  assign n46056 = ~n45448 & ~n45560;
  assign n46057 = ~n45561 & ~n45567;
  assign n46058 = ~n46056 & n46057;
  assign n46059 = ~n46054 & ~n46055;
  assign n46060 = n46058 & n46059;
  assign n46061 = ~n46058 & ~n46059;
  assign n46062 = ~n46060 & ~n46061;
  assign n46063 = ~n45444 & n45445;
  assign n46064 = ~n45444 & n45570;
  assign n46065 = ~n45575 & ~n46063;
  assign n46066 = ~n46064 & n46065;
  assign n46067 = P4_DATAO_REG_7_ & n44388;
  assign n46068 = ~n46062 & ~n46066;
  assign n46069 = ~n46067 & n46068;
  assign n46070 = ~n46062 & n46066;
  assign n46071 = n46067 & n46070;
  assign n46072 = ~n46066 & n46067;
  assign n46073 = n46066 & ~n46067;
  assign n46074 = ~n46072 & ~n46073;
  assign n46075 = n46062 & ~n46074;
  assign n46076 = ~n46069 & ~n46071;
  assign n46077 = ~n46075 & n46076;
  assign n46078 = n45918 & ~n46077;
  assign n46079 = ~n45918 & n46077;
  assign n46080 = ~n46078 & ~n46079;
  assign n46081 = n45917 & ~n46080;
  assign n46082 = n45918 & n46077;
  assign n46083 = ~n45918 & ~n46077;
  assign n46084 = ~n46082 & ~n46083;
  assign n46085 = ~n45917 & ~n46084;
  assign n46086 = ~n46081 & ~n46085;
  assign n46087 = n45914 & ~n46086;
  assign n46088 = ~n45914 & n46086;
  assign n46089 = ~n46087 & ~n46088;
  assign n46090 = n45913 & ~n46089;
  assign n46091 = ~n45914 & ~n46086;
  assign n46092 = ~n45913 & n46091;
  assign n46093 = ~n45913 & n45914;
  assign n46094 = n46086 & n46093;
  assign n46095 = ~n46090 & ~n46092;
  assign n46096 = ~n46094 & n46095;
  assign n46097 = n45911 & ~n46096;
  assign n46098 = ~n45911 & n46096;
  assign n46099 = ~n46097 & ~n46098;
  assign n46100 = n45910 & ~n46099;
  assign n46101 = n45911 & n46096;
  assign n46102 = ~n45911 & ~n46096;
  assign n46103 = ~n46101 & ~n46102;
  assign n46104 = ~n45910 & ~n46103;
  assign n46105 = ~n46100 & ~n46104;
  assign n46106 = n45906 & ~n46105;
  assign n46107 = ~n45906 & n46105;
  assign n46108 = ~n46106 & ~n46107;
  assign n46109 = n45905 & ~n46108;
  assign n46110 = ~n45906 & ~n46105;
  assign n46111 = ~n45905 & n46110;
  assign n46112 = ~n45905 & n45906;
  assign n46113 = n46105 & n46112;
  assign n46114 = ~n46109 & ~n46111;
  assign n46115 = ~n46113 & n46114;
  assign n46116 = n45903 & ~n46115;
  assign n46117 = ~n45903 & n46115;
  assign n46118 = ~n46116 & ~n46117;
  assign n46119 = n44379 & ~n46118;
  assign n46120 = ~n44379 & n46118;
  assign n46121 = P4_DATAO_REG_1_ & n44380;
  assign n46122 = n44383 & n45750;
  assign n46123 = ~n44383 & ~n45750;
  assign n46124 = ~n46122 & ~n46123;
  assign n46125 = ~n45898 & ~n46124;
  assign n46126 = n45898 & n46124;
  assign n46127 = ~n46125 & ~n46126;
  assign n46128 = n46121 & n46127;
  assign n46129 = ~n46121 & ~n46127;
  assign n46130 = P4_DATAO_REG_1_ & n44382;
  assign n46131 = ~n45762 & n45892;
  assign n46132 = ~n45893 & ~n46131;
  assign n46133 = n45769 & ~n46132;
  assign n46134 = ~n45762 & ~n45892;
  assign n46135 = ~n45769 & n46134;
  assign n46136 = n45770 & n45892;
  assign n46137 = ~n46133 & ~n46135;
  assign n46138 = ~n46136 & n46137;
  assign n46139 = P4_DATAO_REG_1_ & n45602;
  assign n46140 = n46138 & n46139;
  assign n46141 = ~n46138 & ~n46139;
  assign n46142 = P4_DATAO_REG_1_ & n44384;
  assign n46143 = P4_DATAO_REG_1_ & n44386;
  assign n46144 = P4_DATAO_REG_1_ & n44388;
  assign n46145 = ~n45790 & n45791;
  assign n46146 = n45790 & ~n45791;
  assign n46147 = ~n46145 & ~n46146;
  assign n46148 = n45876 & ~n46147;
  assign n46149 = ~n45792 & ~n45793;
  assign n46150 = ~n45876 & ~n46149;
  assign n46151 = ~n46148 & ~n46150;
  assign n46152 = n46144 & ~n46151;
  assign n46153 = ~n45794 & n45872;
  assign n46154 = ~n45873 & ~n46153;
  assign n46155 = n45864 & ~n46154;
  assign n46156 = ~n45794 & ~n45872;
  assign n46157 = ~n45864 & n46156;
  assign n46158 = n45865 & n45872;
  assign n46159 = ~n46155 & ~n46157;
  assign n46160 = ~n46158 & n46159;
  assign n46161 = P4_DATAO_REG_1_ & n44390;
  assign n46162 = n46160 & n46161;
  assign n46163 = ~n46160 & ~n46161;
  assign n46164 = P4_DATAO_REG_1_ & n44392;
  assign n46165 = ~n45802 & n45803;
  assign n46166 = n45802 & ~n45803;
  assign n46167 = ~n46165 & ~n46166;
  assign n46168 = n45862 & ~n46167;
  assign n46169 = ~n45804 & ~n45805;
  assign n46170 = ~n45862 & ~n46169;
  assign n46171 = ~n46168 & ~n46170;
  assign n46172 = n46164 & ~n46171;
  assign n46173 = ~n46164 & n46171;
  assign n46174 = P4_DATAO_REG_1_ & n44394;
  assign n46175 = P4_DATAO_REG_1_ & n44704;
  assign n46176 = ~n45818 & n45834;
  assign n46177 = ~n45835 & ~n46176;
  assign n46178 = n45844 & ~n46177;
  assign n46179 = ~n45818 & ~n45834;
  assign n46180 = ~n45844 & n46179;
  assign n46181 = n45834 & n45845;
  assign n46182 = ~n46178 & ~n46180;
  assign n46183 = ~n46181 & n46182;
  assign n46184 = P4_DATAO_REG_1_ & n44623;
  assign n46185 = n46183 & n46184;
  assign n46186 = ~n46183 & ~n46184;
  assign n46187 = P4_DATAO_REG_1_ & n44356;
  assign n46188 = n45827 & ~n45832;
  assign n46189 = ~n45827 & n45832;
  assign n46190 = ~n46188 & ~n46189;
  assign n46191 = ~n45826 & n46190;
  assign n46192 = n45826 & n46189;
  assign n46193 = ~n46191 & ~n46192;
  assign n46194 = n45828 & ~n45832;
  assign n46195 = n46193 & ~n46194;
  assign n46196 = n46187 & ~n46195;
  assign n46197 = ~n46187 & n46195;
  assign n46198 = ~n44286 & ~n44352;
  assign n46199 = ~n44351 & ~n46198;
  assign n46200 = ~n46197 & ~n46199;
  assign n46201 = ~n46196 & ~n46200;
  assign n46202 = ~n46186 & ~n46201;
  assign n46203 = ~n46185 & ~n46202;
  assign n46204 = n46175 & ~n46203;
  assign n46205 = ~n45814 & n45815;
  assign n46206 = n45814 & ~n45815;
  assign n46207 = ~n46205 & ~n46206;
  assign n46208 = n45848 & ~n46207;
  assign n46209 = ~n45816 & ~n45817;
  assign n46210 = ~n45848 & ~n46209;
  assign n46211 = ~n46208 & ~n46210;
  assign n46212 = n46175 & ~n46211;
  assign n46213 = ~n46203 & ~n46211;
  assign n46214 = ~n46204 & ~n46212;
  assign n46215 = ~n46213 & n46214;
  assign n46216 = n46174 & ~n46215;
  assign n46217 = ~n45806 & n45858;
  assign n46218 = ~n45859 & ~n46217;
  assign n46219 = n45850 & ~n46218;
  assign n46220 = ~n45806 & ~n45858;
  assign n46221 = ~n45850 & n46220;
  assign n46222 = n45851 & n45858;
  assign n46223 = ~n46219 & ~n46221;
  assign n46224 = ~n46222 & n46223;
  assign n46225 = ~n46174 & n46215;
  assign n46226 = n46224 & ~n46225;
  assign n46227 = ~n46216 & ~n46226;
  assign n46228 = ~n46173 & ~n46227;
  assign n46229 = ~n46172 & ~n46228;
  assign n46230 = ~n46163 & ~n46229;
  assign n46231 = ~n46162 & ~n46230;
  assign n46232 = n46144 & ~n46231;
  assign n46233 = ~n46151 & ~n46231;
  assign n46234 = ~n46152 & ~n46232;
  assign n46235 = ~n46233 & n46234;
  assign n46236 = n46143 & ~n46235;
  assign n46237 = ~n45782 & n45886;
  assign n46238 = ~n45887 & ~n46237;
  assign n46239 = n45878 & ~n46238;
  assign n46240 = ~n45782 & ~n45886;
  assign n46241 = ~n45878 & n46240;
  assign n46242 = n45879 & n45886;
  assign n46243 = ~n46239 & ~n46241;
  assign n46244 = ~n46242 & n46243;
  assign n46245 = ~n46143 & n46235;
  assign n46246 = n46244 & ~n46245;
  assign n46247 = ~n46236 & ~n46246;
  assign n46248 = n46142 & ~n46247;
  assign n46249 = ~n45778 & n45779;
  assign n46250 = n45778 & ~n45779;
  assign n46251 = ~n46249 & ~n46250;
  assign n46252 = n45890 & ~n46251;
  assign n46253 = ~n45780 & ~n45781;
  assign n46254 = ~n45890 & ~n46253;
  assign n46255 = ~n46252 & ~n46254;
  assign n46256 = n46142 & ~n46255;
  assign n46257 = ~n46247 & ~n46255;
  assign n46258 = ~n46248 & ~n46256;
  assign n46259 = ~n46257 & n46258;
  assign n46260 = ~n46141 & ~n46259;
  assign n46261 = ~n46140 & ~n46260;
  assign n46262 = n46130 & ~n46261;
  assign n46263 = ~n45760 & ~n45761;
  assign n46264 = n45896 & n46263;
  assign n46265 = ~n45896 & ~n46263;
  assign n46266 = ~n46264 & ~n46265;
  assign n46267 = n46130 & ~n46266;
  assign n46268 = ~n46261 & ~n46266;
  assign n46269 = ~n46262 & ~n46267;
  assign n46270 = ~n46268 & n46269;
  assign n46271 = ~n46129 & ~n46270;
  assign n46272 = ~n46128 & ~n46271;
  assign n46273 = ~n46120 & ~n46272;
  assign n46274 = ~n46119 & ~n46273;
  assign n46275 = n44377 & ~n46274;
  assign n46276 = P4_DATAO_REG_2_ & n44378;
  assign n46277 = ~n45902 & n46115;
  assign n46278 = ~n45901 & ~n46277;
  assign n46279 = n46276 & ~n46278;
  assign n46280 = ~n45905 & ~n46105;
  assign n46281 = ~n46106 & ~n46112;
  assign n46282 = ~n46280 & n46281;
  assign n46283 = P4_DATAO_REG_3_ & n44380;
  assign n46284 = ~n46062 & n46067;
  assign n46285 = ~n46072 & ~n46284;
  assign n46286 = ~n46068 & n46285;
  assign n46287 = P4_DATAO_REG_7_ & n44386;
  assign n46288 = P4_DATAO_REG_10_ & n44392;
  assign n46289 = ~n45927 & ~n46043;
  assign n46290 = ~n46042 & ~n46289;
  assign n46291 = n46288 & ~n46290;
  assign n46292 = ~n46288 & n46290;
  assign n46293 = ~n46291 & ~n46292;
  assign n46294 = ~n46023 & ~n46026;
  assign n46295 = ~n46029 & ~n46034;
  assign n46296 = ~n46294 & n46295;
  assign n46297 = P4_DATAO_REG_11_ & n44394;
  assign n46298 = P4_DATAO_REG_13_ & n44623;
  assign n46299 = ~n45999 & n46000;
  assign n46300 = ~n45999 & ~n46004;
  assign n46301 = ~n46011 & ~n46299;
  assign n46302 = ~n46300 & n46301;
  assign n46303 = n46298 & ~n46302;
  assign n46304 = ~n46298 & n46302;
  assign n46305 = ~n46303 & ~n46304;
  assign n46306 = ~n45941 & ~n45986;
  assign n46307 = ~n45987 & ~n45993;
  assign n46308 = ~n46306 & n46307;
  assign n46309 = P4_DATAO_REG_15_ & n44102;
  assign n46310 = ~n45963 & ~n45966;
  assign n46311 = ~n45969 & ~n45974;
  assign n46312 = ~n46310 & n46311;
  assign n46313 = P4_DATAO_REG_17_ & n44143;
  assign n46314 = P4_DATAO_REG_19_ & n44108;
  assign n46315 = P4_DATAO_REG_20_ & n44110;
  assign n46316 = P4_DATAO_REG_21_ & n44112;
  assign n46317 = n46315 & ~n46316;
  assign n46318 = ~n46315 & n46316;
  assign n46319 = ~n46317 & ~n46318;
  assign n46320 = n46314 & ~n46319;
  assign n46321 = ~n46314 & n46319;
  assign n46322 = P4_DATAO_REG_19_ & P4_DATAO_REG_20_;
  assign n46323 = n44119 & n46322;
  assign n46324 = ~n46320 & ~n46321;
  assign n46325 = ~n46323 & n46324;
  assign n46326 = n46314 & ~n46317;
  assign n46327 = ~n46314 & n46317;
  assign n46328 = ~n46326 & ~n46327;
  assign n46329 = n46323 & n46328;
  assign n46330 = ~n46325 & ~n46329;
  assign n46331 = P4_DATAO_REG_18_ & n44106;
  assign n46332 = ~n45955 & n45957;
  assign n46333 = ~n45954 & ~n46332;
  assign n46334 = ~n46330 & ~n46331;
  assign n46335 = ~n46333 & n46334;
  assign n46336 = n46330 & n46331;
  assign n46337 = ~n46334 & ~n46336;
  assign n46338 = n46333 & n46337;
  assign n46339 = ~n46335 & ~n46338;
  assign n46340 = n46331 & ~n46333;
  assign n46341 = n46330 & n46340;
  assign n46342 = n46339 & ~n46341;
  assign n46343 = n46313 & ~n46342;
  assign n46344 = ~n46313 & n46342;
  assign n46345 = ~n46343 & ~n46344;
  assign n46346 = n46312 & ~n46345;
  assign n46347 = ~n46313 & n46341;
  assign n46348 = ~n46313 & ~n46339;
  assign n46349 = n46313 & n46339;
  assign n46350 = ~n46341 & n46349;
  assign n46351 = ~n46347 & ~n46348;
  assign n46352 = ~n46350 & n46351;
  assign n46353 = ~n46312 & ~n46352;
  assign n46354 = ~n46346 & ~n46353;
  assign n46355 = P4_DATAO_REG_16_ & n44104;
  assign n46356 = ~n45946 & ~n45983;
  assign n46357 = ~n45982 & ~n46356;
  assign n46358 = ~n46354 & ~n46355;
  assign n46359 = ~n46357 & n46358;
  assign n46360 = n46354 & n46355;
  assign n46361 = ~n46358 & ~n46360;
  assign n46362 = n46357 & n46361;
  assign n46363 = ~n46359 & ~n46362;
  assign n46364 = n46355 & ~n46357;
  assign n46365 = n46354 & n46364;
  assign n46366 = n46363 & ~n46365;
  assign n46367 = n46309 & ~n46366;
  assign n46368 = ~n46309 & n46366;
  assign n46369 = ~n46367 & ~n46368;
  assign n46370 = n46308 & ~n46369;
  assign n46371 = ~n46309 & n46365;
  assign n46372 = ~n46309 & ~n46363;
  assign n46373 = n46309 & ~n46365;
  assign n46374 = n46363 & n46373;
  assign n46375 = ~n46371 & ~n46372;
  assign n46376 = ~n46374 & n46375;
  assign n46377 = ~n46308 & ~n46376;
  assign n46378 = ~n46370 & ~n46377;
  assign n46379 = P4_DATAO_REG_14_ & n44356;
  assign n46380 = ~n45938 & n45996;
  assign n46381 = ~n45937 & ~n46380;
  assign n46382 = ~n46378 & ~n46379;
  assign n46383 = ~n46381 & n46382;
  assign n46384 = ~n46378 & n46379;
  assign n46385 = n46378 & ~n46379;
  assign n46386 = ~n46384 & ~n46385;
  assign n46387 = n46381 & ~n46386;
  assign n46388 = ~n46383 & ~n46387;
  assign n46389 = n46379 & ~n46381;
  assign n46390 = n46378 & n46389;
  assign n46391 = n46388 & ~n46390;
  assign n46392 = n46305 & ~n46391;
  assign n46393 = ~n46298 & ~n46300;
  assign n46394 = ~n46011 & n46393;
  assign n46395 = ~n46299 & n46394;
  assign n46396 = ~n46303 & ~n46395;
  assign n46397 = n46391 & ~n46396;
  assign n46398 = ~n46392 & ~n46397;
  assign n46399 = P4_DATAO_REG_12_ & n44704;
  assign n46400 = ~n45931 & ~n46020;
  assign n46401 = ~n46019 & ~n46400;
  assign n46402 = ~n46398 & ~n46399;
  assign n46403 = ~n46401 & n46402;
  assign n46404 = ~n46398 & n46399;
  assign n46405 = n46398 & ~n46399;
  assign n46406 = ~n46404 & ~n46405;
  assign n46407 = n46401 & ~n46406;
  assign n46408 = ~n46403 & ~n46407;
  assign n46409 = n46399 & ~n46401;
  assign n46410 = n46398 & n46409;
  assign n46411 = n46408 & ~n46410;
  assign n46412 = n46297 & ~n46411;
  assign n46413 = ~n46297 & n46411;
  assign n46414 = ~n46412 & ~n46413;
  assign n46415 = n46296 & ~n46414;
  assign n46416 = n46297 & ~n46410;
  assign n46417 = n46408 & n46416;
  assign n46418 = ~n46297 & ~n46411;
  assign n46419 = ~n46417 & ~n46418;
  assign n46420 = ~n46296 & ~n46419;
  assign n46421 = ~n46415 & ~n46420;
  assign n46422 = ~n46293 & n46421;
  assign n46423 = n46293 & ~n46421;
  assign n46424 = ~n46422 & ~n46423;
  assign n46425 = P4_DATAO_REG_9_ & n44390;
  assign n46426 = ~n46424 & ~n46425;
  assign n46427 = n46424 & n46425;
  assign n46428 = ~n44392 & n46046;
  assign n46429 = ~n45922 & ~n46428;
  assign n46430 = ~n46047 & ~n46429;
  assign n46431 = ~n46426 & ~n46427;
  assign n46432 = n46430 & n46431;
  assign n46433 = ~n46430 & ~n46431;
  assign n46434 = ~n46432 & ~n46433;
  assign n46435 = P4_DATAO_REG_8_ & n44388;
  assign n46436 = n46053 & ~n46058;
  assign n46437 = n46052 & ~n46058;
  assign n46438 = ~n46055 & ~n46436;
  assign n46439 = ~n46437 & n46438;
  assign n46440 = ~n46434 & ~n46435;
  assign n46441 = ~n46439 & n46440;
  assign n46442 = ~n46434 & n46435;
  assign n46443 = n46434 & ~n46435;
  assign n46444 = ~n46442 & ~n46443;
  assign n46445 = n46439 & ~n46444;
  assign n46446 = ~n46441 & ~n46445;
  assign n46447 = n46435 & ~n46439;
  assign n46448 = n46434 & n46447;
  assign n46449 = n46446 & ~n46448;
  assign n46450 = n46287 & ~n46449;
  assign n46451 = ~n46287 & n46449;
  assign n46452 = ~n46450 & ~n46451;
  assign n46453 = n46286 & ~n46452;
  assign n46454 = n46287 & n46446;
  assign n46455 = ~n46448 & n46454;
  assign n46456 = ~n46287 & ~n46449;
  assign n46457 = ~n46455 & ~n46456;
  assign n46458 = ~n46286 & ~n46457;
  assign n46459 = ~n46453 & ~n46458;
  assign n46460 = P4_DATAO_REG_6_ & n44384;
  assign n46461 = ~n46459 & ~n46460;
  assign n46462 = n46459 & n46460;
  assign n46463 = ~n46461 & ~n46462;
  assign n46464 = ~n45917 & ~n46083;
  assign n46465 = ~n46082 & ~n46464;
  assign n46466 = ~n46463 & ~n46465;
  assign n46467 = ~n46459 & n46460;
  assign n46468 = n46459 & ~n46460;
  assign n46469 = ~n46467 & ~n46468;
  assign n46470 = n46465 & ~n46469;
  assign n46471 = ~n46466 & ~n46470;
  assign n46472 = P4_DATAO_REG_5_ & n45602;
  assign n46473 = ~n46471 & ~n46472;
  assign n46474 = n46471 & n46472;
  assign n46475 = ~n45913 & ~n46086;
  assign n46476 = ~n46087 & ~n46093;
  assign n46477 = ~n46475 & n46476;
  assign n46478 = ~n46473 & ~n46474;
  assign n46479 = n46477 & n46478;
  assign n46480 = ~n46477 & ~n46478;
  assign n46481 = ~n46479 & ~n46480;
  assign n46482 = P4_DATAO_REG_4_ & n44382;
  assign n46483 = ~n45910 & ~n46102;
  assign n46484 = ~n46101 & ~n46483;
  assign n46485 = ~n46481 & ~n46482;
  assign n46486 = ~n46484 & n46485;
  assign n46487 = ~n46481 & n46482;
  assign n46488 = n46481 & ~n46482;
  assign n46489 = ~n46487 & ~n46488;
  assign n46490 = n46484 & ~n46489;
  assign n46491 = ~n46486 & ~n46490;
  assign n46492 = n46482 & ~n46484;
  assign n46493 = n46481 & n46492;
  assign n46494 = n46491 & ~n46493;
  assign n46495 = n46283 & ~n46494;
  assign n46496 = ~n46283 & n46494;
  assign n46497 = ~n46495 & ~n46496;
  assign n46498 = n46282 & ~n46497;
  assign n46499 = n46283 & n46494;
  assign n46500 = ~n46283 & ~n46494;
  assign n46501 = ~n46499 & ~n46500;
  assign n46502 = ~n46282 & ~n46501;
  assign n46503 = ~n46498 & ~n46502;
  assign n46504 = n46279 & n46503;
  assign n46505 = ~n46276 & ~n46503;
  assign n46506 = ~n46278 & n46505;
  assign n46507 = n46276 & ~n46503;
  assign n46508 = ~n46276 & n46503;
  assign n46509 = ~n46507 & ~n46508;
  assign n46510 = n46278 & ~n46509;
  assign n46511 = ~n46506 & ~n46510;
  assign n46512 = ~n44377 & n46274;
  assign n46513 = ~n46504 & n46511;
  assign n46514 = ~n46512 & n46513;
  assign n46515 = ~n46275 & ~n46514;
  assign n46516 = n44375 & ~n46515;
  assign n46517 = ~n46278 & ~n46503;
  assign n46518 = ~n46279 & ~n46507;
  assign n46519 = ~n46517 & n46518;
  assign n46520 = P4_DATAO_REG_2_ & n44376;
  assign n46521 = ~n46282 & ~n46500;
  assign n46522 = ~n46499 & ~n46521;
  assign n46523 = P4_DATAO_REG_3_ & n44378;
  assign n46524 = P4_DATAO_REG_5_ & n44382;
  assign n46525 = ~n46473 & ~n46477;
  assign n46526 = ~n46474 & ~n46525;
  assign n46527 = n46524 & ~n46526;
  assign n46528 = ~n46524 & n46526;
  assign n46529 = ~n46527 & ~n46528;
  assign n46530 = ~n46465 & ~n46468;
  assign n46531 = ~n46467 & ~n46530;
  assign n46532 = P4_DATAO_REG_6_ & n45602;
  assign n46533 = ~n46286 & ~n46456;
  assign n46534 = ~n46455 & ~n46533;
  assign n46535 = P4_DATAO_REG_7_ & n44384;
  assign n46536 = P4_DATAO_REG_8_ & n44386;
  assign n46537 = ~n46434 & ~n46439;
  assign n46538 = ~n46442 & ~n46447;
  assign n46539 = ~n46537 & n46538;
  assign n46540 = n46536 & ~n46539;
  assign n46541 = ~n46536 & n46539;
  assign n46542 = n46288 & ~n46421;
  assign n46543 = ~n46288 & n46421;
  assign n46544 = ~n46290 & ~n46543;
  assign n46545 = ~n46542 & ~n46544;
  assign n46546 = P4_DATAO_REG_10_ & n44390;
  assign n46547 = P4_DATAO_REG_12_ & n44394;
  assign n46548 = ~n46398 & ~n46401;
  assign n46549 = ~n46404 & ~n46409;
  assign n46550 = ~n46548 & n46549;
  assign n46551 = n46547 & ~n46550;
  assign n46552 = ~n46547 & n46550;
  assign n46553 = ~n46551 & ~n46552;
  assign n46554 = P4_DATAO_REG_13_ & n44704;
  assign n46555 = ~n46304 & n46391;
  assign n46556 = ~n46303 & ~n46555;
  assign n46557 = ~n46554 & ~n46556;
  assign n46558 = ~n46378 & ~n46381;
  assign n46559 = ~n46384 & ~n46389;
  assign n46560 = ~n46558 & n46559;
  assign n46561 = P4_DATAO_REG_14_ & n44623;
  assign n46562 = ~n46309 & ~n46366;
  assign n46563 = ~n46308 & ~n46562;
  assign n46564 = ~n46374 & ~n46563;
  assign n46565 = ~n46354 & n46355;
  assign n46566 = ~n46354 & ~n46357;
  assign n46567 = ~n46364 & ~n46565;
  assign n46568 = ~n46566 & n46567;
  assign n46569 = P4_DATAO_REG_16_ & n44102;
  assign n46570 = ~n46330 & n46331;
  assign n46571 = ~n46330 & ~n46333;
  assign n46572 = ~n46340 & ~n46570;
  assign n46573 = ~n46571 & n46572;
  assign n46574 = P4_DATAO_REG_18_ & n44143;
  assign n46575 = P4_DATAO_REG_20_ & n44108;
  assign n46576 = P4_DATAO_REG_21_ & n44110;
  assign n46577 = P4_DATAO_REG_22_ & n44112;
  assign n46578 = n46576 & ~n46577;
  assign n46579 = ~n46576 & n46577;
  assign n46580 = ~n46578 & ~n46579;
  assign n46581 = n46575 & ~n46580;
  assign n46582 = ~n46575 & n46580;
  assign n46583 = P4_DATAO_REG_20_ & P4_DATAO_REG_21_;
  assign n46584 = n44119 & n46583;
  assign n46585 = ~n46581 & ~n46582;
  assign n46586 = ~n46584 & n46585;
  assign n46587 = ~n46575 & ~n46578;
  assign n46588 = n46575 & ~n46577;
  assign n46589 = ~n46587 & ~n46588;
  assign n46590 = n46584 & ~n46589;
  assign n46591 = ~n46586 & ~n46590;
  assign n46592 = P4_DATAO_REG_19_ & n44106;
  assign n46593 = ~n46321 & n46323;
  assign n46594 = ~n46320 & ~n46593;
  assign n46595 = ~n46591 & ~n46592;
  assign n46596 = ~n46594 & n46595;
  assign n46597 = n46591 & n46592;
  assign n46598 = ~n46595 & ~n46597;
  assign n46599 = n46594 & n46598;
  assign n46600 = ~n46596 & ~n46599;
  assign n46601 = n46592 & ~n46594;
  assign n46602 = n46591 & n46601;
  assign n46603 = n46600 & ~n46602;
  assign n46604 = n46574 & ~n46603;
  assign n46605 = ~n46574 & n46603;
  assign n46606 = ~n46604 & ~n46605;
  assign n46607 = n46573 & ~n46606;
  assign n46608 = ~n46574 & n46602;
  assign n46609 = ~n46574 & ~n46600;
  assign n46610 = n46574 & n46600;
  assign n46611 = ~n46602 & n46610;
  assign n46612 = ~n46608 & ~n46609;
  assign n46613 = ~n46611 & n46612;
  assign n46614 = ~n46573 & ~n46613;
  assign n46615 = ~n46607 & ~n46614;
  assign n46616 = P4_DATAO_REG_17_ & n44104;
  assign n46617 = ~n46313 & ~n46342;
  assign n46618 = ~n46312 & ~n46617;
  assign n46619 = ~n46350 & ~n46618;
  assign n46620 = ~n46615 & ~n46616;
  assign n46621 = ~n46619 & n46620;
  assign n46622 = n46615 & n46616;
  assign n46623 = ~n46620 & ~n46622;
  assign n46624 = n46619 & n46623;
  assign n46625 = ~n46621 & ~n46624;
  assign n46626 = n46616 & ~n46619;
  assign n46627 = n46615 & n46626;
  assign n46628 = n46625 & ~n46627;
  assign n46629 = n46569 & ~n46628;
  assign n46630 = ~n46569 & n46628;
  assign n46631 = ~n46629 & ~n46630;
  assign n46632 = n46568 & ~n46631;
  assign n46633 = n46569 & ~n46627;
  assign n46634 = n46625 & n46633;
  assign n46635 = ~n46569 & ~n46628;
  assign n46636 = ~n46634 & ~n46635;
  assign n46637 = ~n46568 & ~n46636;
  assign n46638 = ~n46632 & ~n46637;
  assign n46639 = P4_DATAO_REG_15_ & n44356;
  assign n46640 = n46564 & ~n46638;
  assign n46641 = n46639 & n46640;
  assign n46642 = n46564 & n46638;
  assign n46643 = ~n46639 & n46642;
  assign n46644 = ~n46641 & ~n46643;
  assign n46645 = ~n46564 & ~n46639;
  assign n46646 = ~n46638 & n46645;
  assign n46647 = ~n46564 & n46639;
  assign n46648 = n46638 & n46647;
  assign n46649 = ~n46646 & ~n46648;
  assign n46650 = n46644 & n46649;
  assign n46651 = n46561 & ~n46650;
  assign n46652 = ~n46561 & n46650;
  assign n46653 = ~n46651 & ~n46652;
  assign n46654 = n46560 & ~n46653;
  assign n46655 = n46561 & n46649;
  assign n46656 = n46644 & n46655;
  assign n46657 = ~n46561 & ~n46650;
  assign n46658 = ~n46656 & ~n46657;
  assign n46659 = ~n46560 & ~n46658;
  assign n46660 = ~n46654 & ~n46659;
  assign n46661 = n46557 & ~n46660;
  assign n46662 = n46554 & ~n46556;
  assign n46663 = ~n46303 & ~n46554;
  assign n46664 = ~n46555 & n46663;
  assign n46665 = ~n46662 & ~n46664;
  assign n46666 = n46660 & ~n46665;
  assign n46667 = ~n46661 & ~n46666;
  assign n46668 = n46554 & ~n46660;
  assign n46669 = n46556 & n46668;
  assign n46670 = n46667 & ~n46669;
  assign n46671 = n46553 & ~n46670;
  assign n46672 = ~n46547 & ~n46548;
  assign n46673 = ~n46409 & n46672;
  assign n46674 = ~n46404 & n46673;
  assign n46675 = ~n46551 & ~n46674;
  assign n46676 = n46670 & ~n46675;
  assign n46677 = ~n46671 & ~n46676;
  assign n46678 = P4_DATAO_REG_11_ & n44392;
  assign n46679 = ~n46677 & ~n46678;
  assign n46680 = ~n46296 & ~n46418;
  assign n46681 = ~n46417 & ~n46680;
  assign n46682 = n46679 & ~n46681;
  assign n46683 = ~n46677 & n46678;
  assign n46684 = n46677 & ~n46678;
  assign n46685 = ~n46683 & ~n46684;
  assign n46686 = n46681 & ~n46685;
  assign n46687 = ~n46682 & ~n46686;
  assign n46688 = n46678 & ~n46681;
  assign n46689 = n46677 & n46688;
  assign n46690 = n46687 & ~n46689;
  assign n46691 = n46546 & ~n46690;
  assign n46692 = ~n46546 & n46690;
  assign n46693 = ~n46691 & ~n46692;
  assign n46694 = n46545 & ~n46693;
  assign n46695 = n46546 & ~n46689;
  assign n46696 = n46687 & n46695;
  assign n46697 = ~n46546 & ~n46690;
  assign n46698 = ~n46696 & ~n46697;
  assign n46699 = ~n46545 & ~n46698;
  assign n46700 = ~n46694 & ~n46699;
  assign n46701 = P4_DATAO_REG_9_ & n44388;
  assign n46702 = ~n46426 & ~n46430;
  assign n46703 = ~n46427 & ~n46702;
  assign n46704 = ~n46700 & ~n46701;
  assign n46705 = ~n46703 & n46704;
  assign n46706 = ~n46700 & n46701;
  assign n46707 = n46700 & ~n46701;
  assign n46708 = ~n46706 & ~n46707;
  assign n46709 = n46703 & ~n46708;
  assign n46710 = ~n46705 & ~n46709;
  assign n46711 = n46701 & ~n46703;
  assign n46712 = n46700 & n46711;
  assign n46713 = n46710 & ~n46712;
  assign n46714 = ~n46540 & ~n46541;
  assign n46715 = ~n46713 & n46714;
  assign n46716 = ~n46536 & ~n46537;
  assign n46717 = ~n46447 & n46716;
  assign n46718 = ~n46442 & n46717;
  assign n46719 = ~n46540 & ~n46718;
  assign n46720 = n46713 & ~n46719;
  assign n46721 = ~n46715 & ~n46720;
  assign n46722 = n46535 & ~n46721;
  assign n46723 = ~n46535 & n46721;
  assign n46724 = ~n46722 & ~n46723;
  assign n46725 = n46534 & ~n46724;
  assign n46726 = ~n46535 & ~n46721;
  assign n46727 = ~n46534 & n46726;
  assign n46728 = ~n46534 & n46535;
  assign n46729 = n46721 & n46728;
  assign n46730 = ~n46725 & ~n46727;
  assign n46731 = ~n46729 & n46730;
  assign n46732 = n46532 & ~n46731;
  assign n46733 = ~n46532 & n46731;
  assign n46734 = ~n46732 & ~n46733;
  assign n46735 = n46531 & ~n46734;
  assign n46736 = n46532 & n46731;
  assign n46737 = ~n46532 & ~n46731;
  assign n46738 = ~n46736 & ~n46737;
  assign n46739 = ~n46531 & ~n46738;
  assign n46740 = ~n46735 & ~n46739;
  assign n46741 = ~n46529 & n46740;
  assign n46742 = n46529 & ~n46740;
  assign n46743 = ~n46741 & ~n46742;
  assign n46744 = P4_DATAO_REG_4_ & n44380;
  assign n46745 = ~n46743 & ~n46744;
  assign n46746 = n46743 & n46744;
  assign n46747 = ~n46481 & ~n46484;
  assign n46748 = ~n46487 & ~n46492;
  assign n46749 = ~n46747 & n46748;
  assign n46750 = ~n46745 & ~n46746;
  assign n46751 = n46749 & n46750;
  assign n46752 = ~n46749 & ~n46750;
  assign n46753 = ~n46751 & ~n46752;
  assign n46754 = n46523 & ~n46753;
  assign n46755 = ~n46523 & n46753;
  assign n46756 = ~n46754 & ~n46755;
  assign n46757 = n46522 & ~n46756;
  assign n46758 = ~n46523 & ~n46753;
  assign n46759 = ~n46522 & n46758;
  assign n46760 = n46523 & n46753;
  assign n46761 = ~n46522 & n46760;
  assign n46762 = ~n46757 & ~n46759;
  assign n46763 = ~n46761 & n46762;
  assign n46764 = n46520 & ~n46763;
  assign n46765 = ~n46520 & n46763;
  assign n46766 = ~n46764 & ~n46765;
  assign n46767 = n46519 & ~n46766;
  assign n46768 = n46520 & n46763;
  assign n46769 = ~n46520 & ~n46763;
  assign n46770 = ~n46768 & ~n46769;
  assign n46771 = ~n46519 & ~n46770;
  assign n46772 = ~n46767 & ~n46771;
  assign n46773 = n44375 & ~n46772;
  assign n46774 = ~n46515 & ~n46772;
  assign n46775 = ~n46516 & ~n46773;
  assign n46776 = ~n46774 & n46775;
  assign n46777 = SEL & DIN_22_;
  assign n46778 = P4_DATAO_REG_1_ & n46777;
  assign n46779 = n46776 & ~n46778;
  assign n46780 = ~n46776 & n46778;
  assign n46781 = P4_DATAO_REG_4_ & n44378;
  assign n46782 = ~n46745 & ~n46749;
  assign n46783 = ~n46746 & ~n46782;
  assign n46784 = n46781 & ~n46783;
  assign n46785 = ~n46781 & n46783;
  assign n46786 = ~n46784 & ~n46785;
  assign n46787 = n46524 & ~n46740;
  assign n46788 = ~n46524 & n46740;
  assign n46789 = ~n46526 & ~n46788;
  assign n46790 = ~n46787 & ~n46789;
  assign n46791 = P4_DATAO_REG_5_ & n44380;
  assign n46792 = P4_DATAO_REG_6_ & n44382;
  assign n46793 = ~n46531 & n46532;
  assign n46794 = ~n46531 & n46731;
  assign n46795 = ~n46736 & ~n46793;
  assign n46796 = ~n46794 & n46795;
  assign n46797 = ~n46792 & ~n46796;
  assign n46798 = ~n46534 & ~n46721;
  assign n46799 = ~n46722 & ~n46728;
  assign n46800 = ~n46798 & n46799;
  assign n46801 = P4_DATAO_REG_7_ & n45602;
  assign n46802 = ~n46700 & ~n46703;
  assign n46803 = ~n46706 & ~n46711;
  assign n46804 = ~n46802 & n46803;
  assign n46805 = P4_DATAO_REG_9_ & n44386;
  assign n46806 = ~n46677 & ~n46681;
  assign n46807 = ~n46683 & ~n46688;
  assign n46808 = ~n46806 & n46807;
  assign n46809 = P4_DATAO_REG_11_ & n44390;
  assign n46810 = ~n46556 & ~n46660;
  assign n46811 = ~n46662 & ~n46668;
  assign n46812 = ~n46810 & n46811;
  assign n46813 = P4_DATAO_REG_13_ & n44394;
  assign n46814 = ~n46560 & n46561;
  assign n46815 = ~n46560 & n46650;
  assign n46816 = ~n46656 & ~n46814;
  assign n46817 = ~n46815 & n46816;
  assign n46818 = P4_DATAO_REG_14_ & n44704;
  assign n46819 = n46817 & ~n46818;
  assign n46820 = ~n46638 & n46639;
  assign n46821 = ~n46564 & ~n46638;
  assign n46822 = ~n46647 & ~n46820;
  assign n46823 = ~n46821 & n46822;
  assign n46824 = P4_DATAO_REG_15_ & n44623;
  assign n46825 = P4_DATAO_REG_16_ & n44356;
  assign n46826 = ~n46615 & n46616;
  assign n46827 = ~n46615 & ~n46619;
  assign n46828 = ~n46626 & ~n46826;
  assign n46829 = ~n46827 & n46828;
  assign n46830 = P4_DATAO_REG_17_ & n44102;
  assign n46831 = ~n46591 & n46592;
  assign n46832 = ~n46591 & ~n46594;
  assign n46833 = ~n46601 & ~n46831;
  assign n46834 = ~n46832 & n46833;
  assign n46835 = P4_DATAO_REG_19_ & n44143;
  assign n46836 = P4_DATAO_REG_21_ & n44108;
  assign n46837 = P4_DATAO_REG_22_ & n44110;
  assign n46838 = P4_DATAO_REG_23_ & n44112;
  assign n46839 = n46837 & ~n46838;
  assign n46840 = ~n46837 & n46838;
  assign n46841 = ~n46839 & ~n46840;
  assign n46842 = n46836 & ~n46841;
  assign n46843 = ~n46836 & n46841;
  assign n46844 = P4_DATAO_REG_21_ & P4_DATAO_REG_22_;
  assign n46845 = n44119 & n46844;
  assign n46846 = ~n46842 & ~n46843;
  assign n46847 = ~n46845 & n46846;
  assign n46848 = ~n46836 & ~n46839;
  assign n46849 = n46836 & ~n46838;
  assign n46850 = ~n46848 & ~n46849;
  assign n46851 = n46845 & ~n46850;
  assign n46852 = ~n46847 & ~n46851;
  assign n46853 = P4_DATAO_REG_20_ & n44106;
  assign n46854 = ~n46582 & n46584;
  assign n46855 = ~n46581 & ~n46854;
  assign n46856 = ~n46852 & ~n46853;
  assign n46857 = ~n46855 & n46856;
  assign n46858 = n46852 & n46853;
  assign n46859 = ~n46856 & ~n46858;
  assign n46860 = n46855 & n46859;
  assign n46861 = ~n46857 & ~n46860;
  assign n46862 = n46853 & ~n46855;
  assign n46863 = n46852 & n46862;
  assign n46864 = n46861 & ~n46863;
  assign n46865 = n46835 & ~n46864;
  assign n46866 = ~n46835 & n46864;
  assign n46867 = ~n46865 & ~n46866;
  assign n46868 = n46834 & ~n46867;
  assign n46869 = ~n46835 & n46863;
  assign n46870 = ~n46835 & ~n46861;
  assign n46871 = n46835 & n46861;
  assign n46872 = ~n46863 & n46871;
  assign n46873 = ~n46869 & ~n46870;
  assign n46874 = ~n46872 & n46873;
  assign n46875 = ~n46834 & ~n46874;
  assign n46876 = ~n46868 & ~n46875;
  assign n46877 = P4_DATAO_REG_18_ & n44104;
  assign n46878 = ~n46574 & ~n46603;
  assign n46879 = ~n46573 & ~n46878;
  assign n46880 = ~n46611 & ~n46879;
  assign n46881 = ~n46876 & ~n46877;
  assign n46882 = ~n46880 & n46881;
  assign n46883 = n46876 & n46877;
  assign n46884 = ~n46881 & ~n46883;
  assign n46885 = n46880 & n46884;
  assign n46886 = ~n46882 & ~n46885;
  assign n46887 = n46877 & ~n46880;
  assign n46888 = n46876 & n46887;
  assign n46889 = n46886 & ~n46888;
  assign n46890 = n46830 & ~n46889;
  assign n46891 = ~n46830 & n46889;
  assign n46892 = ~n46890 & ~n46891;
  assign n46893 = n46829 & ~n46892;
  assign n46894 = ~n46830 & n46888;
  assign n46895 = n46830 & ~n46888;
  assign n46896 = n46886 & n46895;
  assign n46897 = ~n46830 & ~n46886;
  assign n46898 = ~n46894 & ~n46896;
  assign n46899 = ~n46897 & n46898;
  assign n46900 = ~n46829 & ~n46899;
  assign n46901 = ~n46893 & ~n46900;
  assign n46902 = n46825 & ~n46901;
  assign n46903 = ~n46569 & n46627;
  assign n46904 = ~n46568 & ~n46903;
  assign n46905 = ~n46569 & ~n46625;
  assign n46906 = n46904 & ~n46905;
  assign n46907 = ~n46634 & ~n46906;
  assign n46908 = n46902 & n46907;
  assign n46909 = ~n46825 & ~n46901;
  assign n46910 = ~n46907 & n46909;
  assign n46911 = ~n46908 & ~n46910;
  assign n46912 = n46825 & ~n46907;
  assign n46913 = ~n46634 & ~n46825;
  assign n46914 = ~n46906 & n46913;
  assign n46915 = ~n46912 & ~n46914;
  assign n46916 = n46901 & ~n46915;
  assign n46917 = n46911 & ~n46916;
  assign n46918 = n46824 & ~n46917;
  assign n46919 = ~n46824 & n46917;
  assign n46920 = ~n46918 & ~n46919;
  assign n46921 = n46823 & ~n46920;
  assign n46922 = ~n46824 & n46901;
  assign n46923 = ~n46915 & n46922;
  assign n46924 = ~n46824 & ~n46911;
  assign n46925 = n46824 & ~n46916;
  assign n46926 = n46911 & n46925;
  assign n46927 = ~n46923 & ~n46924;
  assign n46928 = ~n46926 & n46927;
  assign n46929 = ~n46823 & ~n46928;
  assign n46930 = ~n46921 & ~n46929;
  assign n46931 = n46819 & n46930;
  assign n46932 = ~n46817 & n46818;
  assign n46933 = n46930 & n46932;
  assign n46934 = ~n46931 & ~n46933;
  assign n46935 = n46818 & ~n46930;
  assign n46936 = n46817 & n46935;
  assign n46937 = ~n46818 & ~n46930;
  assign n46938 = ~n46817 & n46937;
  assign n46939 = ~n46936 & ~n46938;
  assign n46940 = n46934 & n46939;
  assign n46941 = n46813 & ~n46940;
  assign n46942 = ~n46813 & n46940;
  assign n46943 = ~n46941 & ~n46942;
  assign n46944 = n46812 & ~n46943;
  assign n46945 = ~n46813 & ~n46939;
  assign n46946 = ~n46813 & ~n46934;
  assign n46947 = n46813 & n46939;
  assign n46948 = n46934 & n46947;
  assign n46949 = ~n46945 & ~n46946;
  assign n46950 = ~n46948 & n46949;
  assign n46951 = ~n46812 & ~n46950;
  assign n46952 = ~n46944 & ~n46951;
  assign n46953 = P4_DATAO_REG_12_ & n44392;
  assign n46954 = ~n46669 & ~n46674;
  assign n46955 = n46667 & n46954;
  assign n46956 = ~n46551 & ~n46955;
  assign n46957 = ~n46952 & ~n46953;
  assign n46958 = ~n46956 & n46957;
  assign n46959 = n46952 & n46953;
  assign n46960 = ~n46957 & ~n46959;
  assign n46961 = n46956 & n46960;
  assign n46962 = ~n46958 & ~n46961;
  assign n46963 = n46953 & ~n46956;
  assign n46964 = n46952 & n46963;
  assign n46965 = n46962 & ~n46964;
  assign n46966 = n46809 & ~n46965;
  assign n46967 = ~n46809 & n46965;
  assign n46968 = ~n46966 & ~n46967;
  assign n46969 = n46808 & ~n46968;
  assign n46970 = ~n46809 & n46964;
  assign n46971 = n46809 & ~n46964;
  assign n46972 = n46962 & n46971;
  assign n46973 = ~n46809 & ~n46962;
  assign n46974 = ~n46970 & ~n46972;
  assign n46975 = ~n46973 & n46974;
  assign n46976 = ~n46808 & ~n46975;
  assign n46977 = ~n46969 & ~n46976;
  assign n46978 = P4_DATAO_REG_10_ & n44388;
  assign n46979 = ~n46545 & ~n46697;
  assign n46980 = ~n46696 & ~n46979;
  assign n46981 = ~n46977 & ~n46978;
  assign n46982 = ~n46980 & n46981;
  assign n46983 = n46977 & n46978;
  assign n46984 = ~n46981 & ~n46983;
  assign n46985 = n46980 & n46984;
  assign n46986 = ~n46982 & ~n46985;
  assign n46987 = n46978 & ~n46980;
  assign n46988 = n46977 & n46987;
  assign n46989 = n46986 & ~n46988;
  assign n46990 = n46805 & ~n46989;
  assign n46991 = ~n46805 & n46989;
  assign n46992 = ~n46990 & ~n46991;
  assign n46993 = n46804 & ~n46992;
  assign n46994 = ~n46805 & n46988;
  assign n46995 = n46805 & ~n46988;
  assign n46996 = n46986 & n46995;
  assign n46997 = ~n46805 & ~n46986;
  assign n46998 = ~n46994 & ~n46996;
  assign n46999 = ~n46997 & n46998;
  assign n47000 = ~n46804 & ~n46999;
  assign n47001 = ~n46993 & ~n47000;
  assign n47002 = P4_DATAO_REG_8_ & n44384;
  assign n47003 = ~n46541 & n46713;
  assign n47004 = ~n46540 & ~n47003;
  assign n47005 = ~n47001 & ~n47002;
  assign n47006 = ~n47004 & n47005;
  assign n47007 = ~n47001 & n47002;
  assign n47008 = n47001 & ~n47002;
  assign n47009 = ~n47007 & ~n47008;
  assign n47010 = n47004 & ~n47009;
  assign n47011 = ~n47006 & ~n47010;
  assign n47012 = n47002 & ~n47004;
  assign n47013 = n47001 & n47012;
  assign n47014 = n47011 & ~n47013;
  assign n47015 = n46801 & ~n47014;
  assign n47016 = ~n46801 & n47014;
  assign n47017 = ~n47015 & ~n47016;
  assign n47018 = n46800 & ~n47017;
  assign n47019 = n46801 & ~n47013;
  assign n47020 = n47011 & n47019;
  assign n47021 = ~n46801 & ~n47014;
  assign n47022 = ~n47020 & ~n47021;
  assign n47023 = ~n46800 & ~n47022;
  assign n47024 = ~n47018 & ~n47023;
  assign n47025 = n46797 & ~n47024;
  assign n47026 = n46792 & ~n46796;
  assign n47027 = ~n46792 & n46796;
  assign n47028 = ~n47026 & ~n47027;
  assign n47029 = n47024 & ~n47028;
  assign n47030 = ~n47025 & ~n47029;
  assign n47031 = n46792 & ~n47024;
  assign n47032 = n46796 & n47031;
  assign n47033 = n47030 & ~n47032;
  assign n47034 = n46791 & ~n47033;
  assign n47035 = ~n46791 & n47033;
  assign n47036 = ~n47034 & ~n47035;
  assign n47037 = n46790 & ~n47036;
  assign n47038 = n46791 & n47030;
  assign n47039 = ~n47032 & n47038;
  assign n47040 = ~n46791 & ~n47033;
  assign n47041 = ~n47039 & ~n47040;
  assign n47042 = ~n46790 & ~n47041;
  assign n47043 = ~n47037 & ~n47042;
  assign n47044 = ~n46786 & n47043;
  assign n47045 = n46786 & ~n47043;
  assign n47046 = ~n47044 & ~n47045;
  assign n47047 = P4_DATAO_REG_3_ & n44376;
  assign n47048 = ~n47046 & ~n47047;
  assign n47049 = n47046 & n47047;
  assign n47050 = ~n46522 & n46523;
  assign n47051 = ~n46522 & ~n46753;
  assign n47052 = ~n46754 & ~n47050;
  assign n47053 = ~n47051 & n47052;
  assign n47054 = ~n47048 & ~n47049;
  assign n47055 = n47053 & n47054;
  assign n47056 = ~n47053 & ~n47054;
  assign n47057 = ~n47055 & ~n47056;
  assign n47058 = P4_DATAO_REG_2_ & n44374;
  assign n47059 = ~n46519 & ~n46769;
  assign n47060 = ~n46768 & ~n47059;
  assign n47061 = ~n47057 & ~n47058;
  assign n47062 = ~n47060 & n47061;
  assign n47063 = ~n47057 & n47058;
  assign n47064 = n47057 & ~n47058;
  assign n47065 = ~n47063 & ~n47064;
  assign n47066 = n47060 & ~n47065;
  assign n47067 = ~n47062 & ~n47066;
  assign n47068 = n47058 & ~n47060;
  assign n47069 = n47057 & n47068;
  assign n47070 = n47067 & ~n47069;
  assign n47071 = ~n46779 & ~n46780;
  assign n47072 = ~n47070 & n47071;
  assign n47073 = n46779 & n47070;
  assign n47074 = n46778 & ~n47069;
  assign n47075 = n47067 & n47074;
  assign n47076 = ~n46776 & n47075;
  assign n47077 = ~n47072 & ~n47073;
  assign n47078 = ~n47076 & n47077;
  assign n47079 = n44373 & ~n47078;
  assign n47080 = ~n44373 & n47078;
  assign n47081 = P4_DATAO_REG_0_ & n46777;
  assign n47082 = P4_DATAO_REG_0_ & n44374;
  assign n47083 = ~n46275 & ~n46512;
  assign n47084 = ~n46513 & n47083;
  assign n47085 = n46513 & ~n47083;
  assign n47086 = ~n47084 & ~n47085;
  assign n47087 = n47082 & ~n47086;
  assign n47088 = ~n47082 & n47086;
  assign n47089 = P4_DATAO_REG_0_ & n44376;
  assign n47090 = P4_DATAO_REG_0_ & n44378;
  assign n47091 = ~n46128 & ~n46129;
  assign n47092 = n46270 & n47091;
  assign n47093 = ~n46270 & ~n47091;
  assign n47094 = ~n47092 & ~n47093;
  assign n47095 = n47090 & ~n47094;
  assign n47096 = ~n47090 & n47094;
  assign n47097 = P4_DATAO_REG_0_ & n44380;
  assign n47098 = P4_DATAO_REG_0_ & n44382;
  assign n47099 = ~n46142 & n46255;
  assign n47100 = ~n46256 & ~n47099;
  assign n47101 = n46247 & ~n47100;
  assign n47102 = ~n46142 & ~n46255;
  assign n47103 = ~n46247 & n47102;
  assign n47104 = n46248 & n46255;
  assign n47105 = ~n47101 & ~n47103;
  assign n47106 = ~n47104 & n47105;
  assign n47107 = P4_DATAO_REG_0_ & n45602;
  assign n47108 = n47106 & n47107;
  assign n47109 = ~n47106 & ~n47107;
  assign n47110 = P4_DATAO_REG_0_ & n44384;
  assign n47111 = ~n46236 & ~n46245;
  assign n47112 = ~n46244 & n47111;
  assign n47113 = n46244 & ~n47111;
  assign n47114 = ~n47112 & ~n47113;
  assign n47115 = n47110 & ~n47114;
  assign n47116 = ~n47110 & n47114;
  assign n47117 = ~n46144 & n46231;
  assign n47118 = ~n46232 & ~n47117;
  assign n47119 = n46151 & ~n47118;
  assign n47120 = ~n46144 & ~n46231;
  assign n47121 = ~n46151 & n47120;
  assign n47122 = n46152 & n46231;
  assign n47123 = ~n47119 & ~n47121;
  assign n47124 = ~n47122 & n47123;
  assign n47125 = P4_DATAO_REG_0_ & n44386;
  assign n47126 = n47124 & n47125;
  assign n47127 = ~n47124 & ~n47125;
  assign n47128 = P4_DATAO_REG_0_ & n44388;
  assign n47129 = ~n46160 & n46161;
  assign n47130 = n46160 & ~n46161;
  assign n47131 = ~n47129 & ~n47130;
  assign n47132 = n46229 & ~n47131;
  assign n47133 = ~n46162 & ~n46163;
  assign n47134 = ~n46229 & ~n47133;
  assign n47135 = ~n47132 & ~n47134;
  assign n47136 = n47128 & ~n47135;
  assign n47137 = ~n47128 & n47135;
  assign n47138 = P4_DATAO_REG_0_ & n44390;
  assign n47139 = n46164 & ~n46227;
  assign n47140 = ~n46164 & n46227;
  assign n47141 = ~n47139 & ~n47140;
  assign n47142 = n46171 & ~n47141;
  assign n47143 = ~n46171 & n47141;
  assign n47144 = ~n47142 & ~n47143;
  assign n47145 = n47138 & n47144;
  assign n47146 = ~n47138 & ~n47144;
  assign n47147 = P4_DATAO_REG_0_ & n44392;
  assign n47148 = ~n46216 & ~n46225;
  assign n47149 = ~n46224 & n47148;
  assign n47150 = n46224 & ~n47148;
  assign n47151 = ~n47149 & ~n47150;
  assign n47152 = n47147 & ~n47151;
  assign n47153 = ~n47147 & n47151;
  assign n47154 = ~n46175 & n46211;
  assign n47155 = ~n46212 & ~n47154;
  assign n47156 = n46203 & ~n47155;
  assign n47157 = ~n46175 & ~n46211;
  assign n47158 = ~n46203 & n47157;
  assign n47159 = n46204 & n46211;
  assign n47160 = ~n47156 & ~n47158;
  assign n47161 = ~n47159 & n47160;
  assign n47162 = P4_DATAO_REG_0_ & n44394;
  assign n47163 = n47161 & n47162;
  assign n47164 = ~n47161 & ~n47162;
  assign n47165 = P4_DATAO_REG_0_ & n44704;
  assign n47166 = n46184 & ~n46201;
  assign n47167 = ~n46184 & n46201;
  assign n47168 = ~n47166 & ~n47167;
  assign n47169 = ~n46183 & n47168;
  assign n47170 = n46183 & n47167;
  assign n47171 = n46185 & ~n46201;
  assign n47172 = ~n47169 & ~n47170;
  assign n47173 = ~n47171 & n47172;
  assign n47174 = n47165 & ~n47173;
  assign n47175 = ~n47165 & n47173;
  assign n47176 = P4_DATAO_REG_0_ & n44623;
  assign n47177 = ~n44283 & ~n44362;
  assign n47178 = ~n44363 & ~n47177;
  assign n47179 = n47176 & ~n47178;
  assign n47180 = n46187 & ~n46199;
  assign n47181 = ~n46187 & n46199;
  assign n47182 = ~n47180 & ~n47181;
  assign n47183 = ~n46195 & ~n47182;
  assign n47184 = n46195 & n47182;
  assign n47185 = ~n47183 & ~n47184;
  assign n47186 = ~n47176 & n47178;
  assign n47187 = ~n47185 & ~n47186;
  assign n47188 = ~n47179 & ~n47187;
  assign n47189 = ~n47175 & ~n47188;
  assign n47190 = ~n47174 & ~n47189;
  assign n47191 = ~n47164 & ~n47190;
  assign n47192 = ~n47163 & ~n47191;
  assign n47193 = ~n47153 & ~n47192;
  assign n47194 = ~n47152 & ~n47193;
  assign n47195 = ~n47146 & ~n47194;
  assign n47196 = ~n47145 & ~n47195;
  assign n47197 = ~n47137 & ~n47196;
  assign n47198 = ~n47136 & ~n47197;
  assign n47199 = ~n47127 & ~n47198;
  assign n47200 = ~n47126 & ~n47199;
  assign n47201 = ~n47116 & ~n47200;
  assign n47202 = ~n47115 & ~n47201;
  assign n47203 = ~n47109 & ~n47202;
  assign n47204 = ~n47108 & ~n47203;
  assign n47205 = n47098 & ~n47204;
  assign n47206 = ~n46138 & n46139;
  assign n47207 = n46138 & ~n46139;
  assign n47208 = ~n47206 & ~n47207;
  assign n47209 = n46259 & ~n47208;
  assign n47210 = ~n46140 & ~n46141;
  assign n47211 = ~n46259 & ~n47210;
  assign n47212 = ~n47209 & ~n47211;
  assign n47213 = ~n47098 & n47204;
  assign n47214 = ~n47212 & ~n47213;
  assign n47215 = ~n47205 & ~n47214;
  assign n47216 = n47097 & ~n47215;
  assign n47217 = ~n46130 & n46266;
  assign n47218 = ~n46267 & ~n47217;
  assign n47219 = n46261 & ~n47218;
  assign n47220 = ~n46130 & ~n46266;
  assign n47221 = ~n46261 & n47220;
  assign n47222 = n46262 & n46266;
  assign n47223 = ~n47219 & ~n47221;
  assign n47224 = ~n47222 & n47223;
  assign n47225 = ~n47097 & n47215;
  assign n47226 = n47224 & ~n47225;
  assign n47227 = ~n47216 & ~n47226;
  assign n47228 = ~n47096 & ~n47227;
  assign n47229 = ~n47095 & ~n47228;
  assign n47230 = n47089 & ~n47229;
  assign n47231 = n44379 & ~n46272;
  assign n47232 = ~n44379 & n46272;
  assign n47233 = ~n47231 & ~n47232;
  assign n47234 = n46118 & ~n47233;
  assign n47235 = ~n46118 & n47233;
  assign n47236 = ~n47234 & ~n47235;
  assign n47237 = ~n47089 & n47229;
  assign n47238 = n47236 & ~n47237;
  assign n47239 = ~n47230 & ~n47238;
  assign n47240 = ~n47088 & ~n47239;
  assign n47241 = ~n47087 & ~n47240;
  assign n47242 = n47081 & ~n47241;
  assign n47243 = ~n44375 & n46772;
  assign n47244 = ~n46773 & ~n47243;
  assign n47245 = n46515 & ~n47244;
  assign n47246 = ~n44375 & ~n46772;
  assign n47247 = ~n46515 & n47246;
  assign n47248 = n46516 & n46772;
  assign n47249 = ~n47245 & ~n47247;
  assign n47250 = ~n47248 & n47249;
  assign n47251 = ~n47081 & n47241;
  assign n47252 = n47250 & ~n47251;
  assign n47253 = ~n47242 & ~n47252;
  assign n47254 = ~n47079 & ~n47080;
  assign n47255 = n47253 & n47254;
  assign n47256 = ~n47253 & ~n47254;
  assign n47257 = ~n47255 & ~n47256;
  assign n47258 = ~n12460 & ~n47257;
  assign n47259 = ~n44371 & ~n47258;
  assign n47260 = n44042 & n44097;
  assign n47261 = ~n47259 & n47260;
  assign n47262 = n44088 & n47261;
  assign n47263 = ~n44093 & ~n44096;
  assign n47264 = ~n44370 & n47263;
  assign n47265 = ~n47262 & n47264;
  assign n47266 = P1_BUF1_REG_31_ & n12460;
  assign n47267 = SEL & DIN_29_;
  assign n47268 = P4_DATAO_REG_1_ & n47267;
  assign n47269 = SEL & DIN_28_;
  assign n47270 = P4_DATAO_REG_1_ & n47269;
  assign n47271 = SEL & DIN_27_;
  assign n47272 = P4_DATAO_REG_2_ & n47271;
  assign n47273 = SEL & DIN_26_;
  assign n47274 = P4_DATAO_REG_2_ & n47273;
  assign n47275 = SEL & DIN_25_;
  assign n47276 = P4_DATAO_REG_2_ & n47275;
  assign n47277 = SEL & DIN_24_;
  assign n47278 = P4_DATAO_REG_2_ & n47277;
  assign n47279 = P4_DATAO_REG_4_ & n44374;
  assign n47280 = P4_DATAO_REG_4_ & n44376;
  assign n47281 = P4_DATAO_REG_5_ & n44378;
  assign n47282 = ~n46790 & ~n47040;
  assign n47283 = ~n47039 & ~n47282;
  assign n47284 = n47281 & ~n47283;
  assign n47285 = ~n46796 & ~n47024;
  assign n47286 = ~n47026 & ~n47031;
  assign n47287 = ~n47285 & n47286;
  assign n47288 = P4_DATAO_REG_6_ & n44380;
  assign n47289 = ~n47001 & ~n47004;
  assign n47290 = ~n47007 & ~n47012;
  assign n47291 = ~n47289 & n47290;
  assign n47292 = P4_DATAO_REG_8_ & n45602;
  assign n47293 = P4_DATAO_REG_12_ & n44390;
  assign n47294 = ~n46952 & n46953;
  assign n47295 = ~n46952 & ~n46956;
  assign n47296 = ~n46963 & ~n47294;
  assign n47297 = ~n47295 & n47296;
  assign n47298 = n47293 & ~n47297;
  assign n47299 = ~n47293 & n47297;
  assign n47300 = P4_DATAO_REG_14_ & n44394;
  assign n47301 = ~n46817 & ~n46930;
  assign n47302 = ~n46932 & ~n46935;
  assign n47303 = ~n47301 & n47302;
  assign n47304 = n47300 & ~n47303;
  assign n47305 = ~n47300 & n47303;
  assign n47306 = ~n47304 & ~n47305;
  assign n47307 = ~n46901 & ~n46907;
  assign n47308 = ~n46902 & ~n46912;
  assign n47309 = ~n47307 & n47308;
  assign n47310 = P4_DATAO_REG_16_ & n44623;
  assign n47311 = ~n46876 & n46877;
  assign n47312 = ~n46876 & ~n46880;
  assign n47313 = ~n46887 & ~n47311;
  assign n47314 = ~n47312 & n47313;
  assign n47315 = P4_DATAO_REG_18_ & n44102;
  assign n47316 = ~n46852 & n46853;
  assign n47317 = ~n46852 & ~n46855;
  assign n47318 = ~n46862 & ~n47316;
  assign n47319 = ~n47317 & n47318;
  assign n47320 = P4_DATAO_REG_20_ & n44143;
  assign n47321 = P4_DATAO_REG_22_ & n44108;
  assign n47322 = P4_DATAO_REG_23_ & n44110;
  assign n47323 = P4_DATAO_REG_24_ & n44112;
  assign n47324 = n47322 & ~n47323;
  assign n47325 = ~n47322 & n47323;
  assign n47326 = ~n47324 & ~n47325;
  assign n47327 = n47321 & ~n47326;
  assign n47328 = ~n47321 & n47326;
  assign n47329 = P4_DATAO_REG_22_ & P4_DATAO_REG_23_;
  assign n47330 = n44119 & n47329;
  assign n47331 = ~n47327 & ~n47328;
  assign n47332 = ~n47330 & n47331;
  assign n47333 = n47321 & ~n47324;
  assign n47334 = ~n47321 & n47324;
  assign n47335 = ~n47333 & ~n47334;
  assign n47336 = n47330 & n47335;
  assign n47337 = ~n47332 & ~n47336;
  assign n47338 = P4_DATAO_REG_21_ & n44106;
  assign n47339 = ~n46843 & n46845;
  assign n47340 = ~n46842 & ~n47339;
  assign n47341 = ~n47337 & ~n47338;
  assign n47342 = ~n47340 & n47341;
  assign n47343 = n47337 & n47338;
  assign n47344 = ~n47341 & ~n47343;
  assign n47345 = n47340 & n47344;
  assign n47346 = ~n47342 & ~n47345;
  assign n47347 = n47338 & ~n47340;
  assign n47348 = n47337 & n47347;
  assign n47349 = n47346 & ~n47348;
  assign n47350 = n47320 & ~n47349;
  assign n47351 = ~n47320 & n47349;
  assign n47352 = ~n47350 & ~n47351;
  assign n47353 = n47319 & ~n47352;
  assign n47354 = ~n47320 & n47348;
  assign n47355 = ~n47320 & ~n47346;
  assign n47356 = n47320 & n47346;
  assign n47357 = ~n47348 & n47356;
  assign n47358 = ~n47354 & ~n47355;
  assign n47359 = ~n47357 & n47358;
  assign n47360 = ~n47319 & ~n47359;
  assign n47361 = ~n47353 & ~n47360;
  assign n47362 = P4_DATAO_REG_19_ & n44104;
  assign n47363 = ~n46835 & ~n46864;
  assign n47364 = ~n46834 & ~n47363;
  assign n47365 = ~n46872 & ~n47364;
  assign n47366 = ~n47361 & ~n47362;
  assign n47367 = ~n47365 & n47366;
  assign n47368 = n47361 & n47362;
  assign n47369 = ~n47366 & ~n47368;
  assign n47370 = n47365 & n47369;
  assign n47371 = ~n47367 & ~n47370;
  assign n47372 = n47362 & ~n47365;
  assign n47373 = n47361 & n47372;
  assign n47374 = n47371 & ~n47373;
  assign n47375 = n47315 & ~n47374;
  assign n47376 = ~n47315 & n47374;
  assign n47377 = ~n47375 & ~n47376;
  assign n47378 = n47314 & ~n47377;
  assign n47379 = ~n47315 & n47373;
  assign n47380 = n47315 & ~n47373;
  assign n47381 = n47371 & n47380;
  assign n47382 = ~n47315 & ~n47371;
  assign n47383 = ~n47379 & ~n47381;
  assign n47384 = ~n47382 & n47383;
  assign n47385 = ~n47314 & ~n47384;
  assign n47386 = ~n47378 & ~n47385;
  assign n47387 = P4_DATAO_REG_17_ & n44356;
  assign n47388 = ~n46830 & ~n46889;
  assign n47389 = ~n46829 & ~n47388;
  assign n47390 = ~n46896 & ~n47389;
  assign n47391 = ~n47386 & ~n47387;
  assign n47392 = ~n47390 & n47391;
  assign n47393 = n47386 & n47387;
  assign n47394 = ~n47391 & ~n47393;
  assign n47395 = n47390 & n47394;
  assign n47396 = ~n47392 & ~n47395;
  assign n47397 = n47387 & ~n47390;
  assign n47398 = n47386 & n47397;
  assign n47399 = n47396 & ~n47398;
  assign n47400 = n47310 & ~n47399;
  assign n47401 = ~n47310 & n47399;
  assign n47402 = ~n47400 & ~n47401;
  assign n47403 = n47309 & ~n47402;
  assign n47404 = ~n47310 & n47398;
  assign n47405 = n47310 & ~n47398;
  assign n47406 = n47396 & n47405;
  assign n47407 = ~n47310 & ~n47396;
  assign n47408 = ~n47404 & ~n47406;
  assign n47409 = ~n47407 & n47408;
  assign n47410 = ~n47309 & ~n47409;
  assign n47411 = ~n47403 & ~n47410;
  assign n47412 = P4_DATAO_REG_15_ & n44704;
  assign n47413 = ~n46824 & ~n46917;
  assign n47414 = ~n46823 & ~n47413;
  assign n47415 = ~n46926 & ~n47414;
  assign n47416 = ~n47411 & ~n47412;
  assign n47417 = ~n47415 & n47416;
  assign n47418 = ~n47411 & n47412;
  assign n47419 = n47411 & ~n47412;
  assign n47420 = ~n47418 & ~n47419;
  assign n47421 = n47415 & ~n47420;
  assign n47422 = ~n47417 & ~n47421;
  assign n47423 = n47412 & ~n47415;
  assign n47424 = n47411 & n47423;
  assign n47425 = n47422 & ~n47424;
  assign n47426 = n47306 & ~n47425;
  assign n47427 = ~n47300 & ~n47301;
  assign n47428 = ~n46932 & n47427;
  assign n47429 = ~n46935 & n47428;
  assign n47430 = ~n47304 & ~n47429;
  assign n47431 = n47425 & ~n47430;
  assign n47432 = ~n47426 & ~n47431;
  assign n47433 = P4_DATAO_REG_13_ & n44392;
  assign n47434 = ~n46812 & n46813;
  assign n47435 = ~n46812 & n46940;
  assign n47436 = ~n46948 & ~n47434;
  assign n47437 = ~n47435 & n47436;
  assign n47438 = ~n47432 & ~n47433;
  assign n47439 = ~n47437 & n47438;
  assign n47440 = n47432 & n47433;
  assign n47441 = ~n47438 & ~n47440;
  assign n47442 = n47437 & n47441;
  assign n47443 = ~n47439 & ~n47442;
  assign n47444 = n47433 & ~n47437;
  assign n47445 = n47432 & n47444;
  assign n47446 = n47443 & ~n47445;
  assign n47447 = ~n47298 & ~n47299;
  assign n47448 = ~n47446 & n47447;
  assign n47449 = ~n47293 & ~n47295;
  assign n47450 = ~n46963 & n47449;
  assign n47451 = ~n47294 & n47450;
  assign n47452 = ~n47298 & ~n47451;
  assign n47453 = n47446 & ~n47452;
  assign n47454 = ~n47448 & ~n47453;
  assign n47455 = P4_DATAO_REG_11_ & n44388;
  assign n47456 = ~n47454 & ~n47455;
  assign n47457 = ~n46809 & ~n46965;
  assign n47458 = ~n46808 & ~n47457;
  assign n47459 = ~n46972 & ~n47458;
  assign n47460 = n47456 & ~n47459;
  assign n47461 = ~n47454 & n47455;
  assign n47462 = n47454 & ~n47455;
  assign n47463 = ~n47461 & ~n47462;
  assign n47464 = n47459 & ~n47463;
  assign n47465 = ~n47460 & ~n47464;
  assign n47466 = n47455 & ~n47459;
  assign n47467 = n47454 & n47466;
  assign n47468 = n47465 & ~n47467;
  assign n47469 = ~n46977 & n46978;
  assign n47470 = ~n46977 & ~n46980;
  assign n47471 = P4_DATAO_REG_10_ & n44386;
  assign n47472 = ~n46987 & ~n47469;
  assign n47473 = ~n47470 & n47472;
  assign n47474 = ~n47471 & n47473;
  assign n47475 = n47471 & ~n47473;
  assign n47476 = ~n47474 & ~n47475;
  assign n47477 = n47468 & ~n47476;
  assign n47478 = ~n47468 & n47476;
  assign n47479 = ~n47477 & ~n47478;
  assign n47480 = P4_DATAO_REG_9_ & n44384;
  assign n47481 = ~n47479 & ~n47480;
  assign n47482 = ~n46805 & ~n46989;
  assign n47483 = ~n46804 & ~n47482;
  assign n47484 = ~n46996 & ~n47483;
  assign n47485 = n47481 & ~n47484;
  assign n47486 = n47479 & n47480;
  assign n47487 = ~n47481 & ~n47486;
  assign n47488 = n47484 & n47487;
  assign n47489 = ~n47485 & ~n47488;
  assign n47490 = n47480 & ~n47484;
  assign n47491 = n47479 & n47490;
  assign n47492 = n47489 & ~n47491;
  assign n47493 = n47292 & ~n47492;
  assign n47494 = ~n47292 & n47492;
  assign n47495 = ~n47493 & ~n47494;
  assign n47496 = n47291 & ~n47495;
  assign n47497 = ~n47292 & n47491;
  assign n47498 = ~n47292 & ~n47489;
  assign n47499 = n47292 & ~n47491;
  assign n47500 = n47489 & n47499;
  assign n47501 = ~n47497 & ~n47498;
  assign n47502 = ~n47500 & n47501;
  assign n47503 = ~n47291 & ~n47502;
  assign n47504 = ~n47496 & ~n47503;
  assign n47505 = P4_DATAO_REG_7_ & n44382;
  assign n47506 = ~n46800 & n46801;
  assign n47507 = ~n46800 & ~n47013;
  assign n47508 = n47011 & n47507;
  assign n47509 = ~n47020 & ~n47506;
  assign n47510 = ~n47508 & n47509;
  assign n47511 = ~n47504 & ~n47505;
  assign n47512 = ~n47510 & n47511;
  assign n47513 = n47504 & n47505;
  assign n47514 = ~n47511 & ~n47513;
  assign n47515 = n47510 & n47514;
  assign n47516 = ~n47512 & ~n47515;
  assign n47517 = ~n47510 & n47513;
  assign n47518 = n47516 & ~n47517;
  assign n47519 = n47288 & ~n47518;
  assign n47520 = ~n47288 & n47518;
  assign n47521 = ~n47519 & ~n47520;
  assign n47522 = n47287 & ~n47521;
  assign n47523 = n47288 & ~n47517;
  assign n47524 = n47516 & n47523;
  assign n47525 = ~n47288 & ~n47518;
  assign n47526 = ~n47524 & ~n47525;
  assign n47527 = ~n47287 & ~n47526;
  assign n47528 = ~n47522 & ~n47527;
  assign n47529 = n47284 & n47528;
  assign n47530 = n47280 & ~n47529;
  assign n47531 = ~n47281 & ~n47528;
  assign n47532 = ~n47283 & n47531;
  assign n47533 = n47281 & ~n47528;
  assign n47534 = ~n47281 & n47528;
  assign n47535 = ~n47533 & ~n47534;
  assign n47536 = n47283 & ~n47535;
  assign n47537 = ~n47532 & ~n47536;
  assign n47538 = n47530 & n47537;
  assign n47539 = ~n47529 & n47537;
  assign n47540 = ~n47280 & ~n47539;
  assign n47541 = n46781 & ~n47043;
  assign n47542 = ~n46781 & n47043;
  assign n47543 = ~n46783 & ~n47542;
  assign n47544 = ~n47541 & ~n47543;
  assign n47545 = ~n47540 & ~n47544;
  assign n47546 = ~n47538 & ~n47545;
  assign n47547 = n47279 & ~n47546;
  assign n47548 = P4_DATAO_REG_5_ & n44376;
  assign n47549 = n47505 & ~n47510;
  assign n47550 = ~n47504 & n47505;
  assign n47551 = ~n47504 & ~n47510;
  assign n47552 = ~n47549 & ~n47550;
  assign n47553 = ~n47551 & n47552;
  assign n47554 = P4_DATAO_REG_7_ & n44380;
  assign n47555 = P4_DATAO_REG_8_ & n44382;
  assign n47556 = ~n47291 & n47501;
  assign n47557 = ~n47500 & ~n47556;
  assign n47558 = ~n47555 & ~n47557;
  assign n47559 = ~n47479 & n47480;
  assign n47560 = ~n47479 & ~n47484;
  assign n47561 = ~n47490 & ~n47559;
  assign n47562 = ~n47560 & n47561;
  assign n47563 = P4_DATAO_REG_9_ & n45602;
  assign n47564 = ~n47454 & ~n47459;
  assign n47565 = ~n47461 & ~n47466;
  assign n47566 = ~n47564 & n47565;
  assign n47567 = P4_DATAO_REG_11_ & n44386;
  assign n47568 = P4_DATAO_REG_14_ & n44392;
  assign n47569 = ~n47305 & n47425;
  assign n47570 = ~n47304 & ~n47569;
  assign n47571 = ~n47411 & ~n47415;
  assign n47572 = ~n47418 & ~n47423;
  assign n47573 = ~n47571 & n47572;
  assign n47574 = P4_DATAO_REG_15_ & n44394;
  assign n47575 = P4_DATAO_REG_16_ & n44704;
  assign n47576 = ~n47310 & ~n47399;
  assign n47577 = ~n47309 & ~n47576;
  assign n47578 = ~n47406 & ~n47577;
  assign n47579 = ~n47386 & n47387;
  assign n47580 = ~n47386 & ~n47390;
  assign n47581 = ~n47397 & ~n47579;
  assign n47582 = ~n47580 & n47581;
  assign n47583 = P4_DATAO_REG_17_ & n44623;
  assign n47584 = P4_DATAO_REG_18_ & n44356;
  assign n47585 = ~n47314 & ~n47379;
  assign n47586 = ~n47382 & n47585;
  assign n47587 = ~n47381 & ~n47586;
  assign n47588 = ~n47584 & ~n47587;
  assign n47589 = ~n47361 & n47362;
  assign n47590 = ~n47361 & ~n47365;
  assign n47591 = ~n47372 & ~n47589;
  assign n47592 = ~n47590 & n47591;
  assign n47593 = P4_DATAO_REG_19_ & n44102;
  assign n47594 = P4_DATAO_REG_20_ & n44104;
  assign n47595 = ~n47337 & n47338;
  assign n47596 = ~n47337 & ~n47340;
  assign n47597 = ~n47347 & ~n47595;
  assign n47598 = ~n47596 & n47597;
  assign n47599 = P4_DATAO_REG_21_ & n44143;
  assign n47600 = P4_DATAO_REG_23_ & n44108;
  assign n47601 = P4_DATAO_REG_24_ & n44110;
  assign n47602 = P4_DATAO_REG_25_ & n44112;
  assign n47603 = n47601 & ~n47602;
  assign n47604 = ~n47601 & n47602;
  assign n47605 = ~n47603 & ~n47604;
  assign n47606 = n47600 & ~n47605;
  assign n47607 = ~n47600 & n47605;
  assign n47608 = P4_DATAO_REG_23_ & P4_DATAO_REG_24_;
  assign n47609 = n44119 & n47608;
  assign n47610 = ~n47606 & ~n47607;
  assign n47611 = ~n47609 & n47610;
  assign n47612 = n47600 & ~n47603;
  assign n47613 = ~n47600 & n47603;
  assign n47614 = ~n47612 & ~n47613;
  assign n47615 = n47609 & n47614;
  assign n47616 = ~n47611 & ~n47615;
  assign n47617 = P4_DATAO_REG_22_ & n44106;
  assign n47618 = ~n47328 & n47330;
  assign n47619 = ~n47327 & ~n47618;
  assign n47620 = ~n47616 & ~n47617;
  assign n47621 = ~n47619 & n47620;
  assign n47622 = n47616 & n47617;
  assign n47623 = ~n47620 & ~n47622;
  assign n47624 = n47619 & n47623;
  assign n47625 = ~n47621 & ~n47624;
  assign n47626 = n47617 & ~n47619;
  assign n47627 = n47616 & n47626;
  assign n47628 = n47625 & ~n47627;
  assign n47629 = n47599 & ~n47628;
  assign n47630 = ~n47599 & n47628;
  assign n47631 = ~n47629 & ~n47630;
  assign n47632 = n47598 & ~n47631;
  assign n47633 = ~n47599 & n47627;
  assign n47634 = ~n47599 & ~n47625;
  assign n47635 = n47599 & n47625;
  assign n47636 = ~n47627 & n47635;
  assign n47637 = ~n47633 & ~n47634;
  assign n47638 = ~n47636 & n47637;
  assign n47639 = ~n47598 & ~n47638;
  assign n47640 = ~n47632 & ~n47639;
  assign n47641 = n47594 & ~n47640;
  assign n47642 = ~n47320 & ~n47349;
  assign n47643 = ~n47319 & ~n47642;
  assign n47644 = ~n47357 & ~n47643;
  assign n47645 = n47641 & n47644;
  assign n47646 = ~n47594 & ~n47640;
  assign n47647 = ~n47644 & n47646;
  assign n47648 = ~n47645 & ~n47647;
  assign n47649 = n47594 & ~n47644;
  assign n47650 = ~n47594 & n47644;
  assign n47651 = ~n47649 & ~n47650;
  assign n47652 = n47640 & ~n47651;
  assign n47653 = n47648 & ~n47652;
  assign n47654 = n47593 & ~n47653;
  assign n47655 = ~n47593 & n47653;
  assign n47656 = ~n47654 & ~n47655;
  assign n47657 = n47592 & ~n47656;
  assign n47658 = n47593 & ~n47652;
  assign n47659 = n47648 & n47658;
  assign n47660 = ~n47593 & ~n47653;
  assign n47661 = ~n47659 & ~n47660;
  assign n47662 = ~n47592 & ~n47661;
  assign n47663 = ~n47657 & ~n47662;
  assign n47664 = n47588 & ~n47663;
  assign n47665 = ~n47584 & n47587;
  assign n47666 = n47584 & ~n47587;
  assign n47667 = ~n47665 & ~n47666;
  assign n47668 = n47663 & ~n47667;
  assign n47669 = ~n47664 & ~n47668;
  assign n47670 = n47584 & n47587;
  assign n47671 = ~n47663 & n47670;
  assign n47672 = n47669 & ~n47671;
  assign n47673 = n47583 & ~n47672;
  assign n47674 = ~n47583 & n47672;
  assign n47675 = ~n47673 & ~n47674;
  assign n47676 = n47582 & ~n47675;
  assign n47677 = n47583 & ~n47671;
  assign n47678 = n47669 & n47677;
  assign n47679 = ~n47583 & ~n47672;
  assign n47680 = ~n47678 & ~n47679;
  assign n47681 = ~n47582 & ~n47680;
  assign n47682 = ~n47676 & ~n47681;
  assign n47683 = ~n47575 & ~n47578;
  assign n47684 = ~n47682 & n47683;
  assign n47685 = n47575 & ~n47578;
  assign n47686 = n47682 & n47685;
  assign n47687 = ~n47684 & ~n47686;
  assign n47688 = ~n47575 & ~n47682;
  assign n47689 = n47575 & n47682;
  assign n47690 = ~n47688 & ~n47689;
  assign n47691 = n47578 & n47690;
  assign n47692 = n47687 & ~n47691;
  assign n47693 = n47574 & ~n47692;
  assign n47694 = ~n47574 & n47692;
  assign n47695 = ~n47693 & ~n47694;
  assign n47696 = n47573 & ~n47695;
  assign n47697 = n47574 & n47687;
  assign n47698 = ~n47691 & n47697;
  assign n47699 = ~n47574 & ~n47692;
  assign n47700 = ~n47698 & ~n47699;
  assign n47701 = ~n47573 & ~n47700;
  assign n47702 = ~n47696 & ~n47701;
  assign n47703 = ~n47568 & ~n47570;
  assign n47704 = ~n47702 & n47703;
  assign n47705 = n47568 & ~n47570;
  assign n47706 = ~n47304 & ~n47568;
  assign n47707 = ~n47569 & n47706;
  assign n47708 = ~n47705 & ~n47707;
  assign n47709 = n47702 & ~n47708;
  assign n47710 = ~n47704 & ~n47709;
  assign n47711 = n47568 & ~n47702;
  assign n47712 = n47570 & n47711;
  assign n47713 = n47710 & ~n47712;
  assign n47714 = ~n47432 & n47433;
  assign n47715 = ~n47432 & ~n47437;
  assign n47716 = P4_DATAO_REG_13_ & n44390;
  assign n47717 = ~n47444 & ~n47714;
  assign n47718 = ~n47715 & n47717;
  assign n47719 = ~n47716 & n47718;
  assign n47720 = n47716 & ~n47718;
  assign n47721 = ~n47719 & ~n47720;
  assign n47722 = n47713 & ~n47721;
  assign n47723 = ~n47713 & n47721;
  assign n47724 = ~n47722 & ~n47723;
  assign n47725 = P4_DATAO_REG_12_ & n44388;
  assign n47726 = n47293 & ~n47445;
  assign n47727 = n47443 & n47726;
  assign n47728 = ~n47297 & n47446;
  assign n47729 = ~n47298 & ~n47727;
  assign n47730 = ~n47728 & n47729;
  assign n47731 = ~n47724 & ~n47725;
  assign n47732 = ~n47730 & n47731;
  assign n47733 = n47724 & n47725;
  assign n47734 = ~n47731 & ~n47733;
  assign n47735 = n47730 & n47734;
  assign n47736 = ~n47732 & ~n47735;
  assign n47737 = n47725 & ~n47730;
  assign n47738 = n47724 & n47737;
  assign n47739 = n47736 & ~n47738;
  assign n47740 = n47567 & ~n47739;
  assign n47741 = ~n47567 & n47739;
  assign n47742 = ~n47740 & ~n47741;
  assign n47743 = n47566 & ~n47742;
  assign n47744 = ~n47567 & ~n47736;
  assign n47745 = n47567 & n47736;
  assign n47746 = ~n47738 & n47745;
  assign n47747 = ~n47567 & n47738;
  assign n47748 = ~n47744 & ~n47746;
  assign n47749 = ~n47747 & n47748;
  assign n47750 = ~n47566 & ~n47749;
  assign n47751 = ~n47743 & ~n47750;
  assign n47752 = P4_DATAO_REG_10_ & n44384;
  assign n47753 = ~n47470 & ~n47471;
  assign n47754 = ~n46987 & n47753;
  assign n47755 = ~n47469 & n47754;
  assign n47756 = ~n47467 & ~n47755;
  assign n47757 = n47465 & n47756;
  assign n47758 = ~n47475 & ~n47757;
  assign n47759 = ~n47751 & ~n47752;
  assign n47760 = ~n47758 & n47759;
  assign n47761 = n47751 & n47752;
  assign n47762 = ~n47759 & ~n47761;
  assign n47763 = n47758 & n47762;
  assign n47764 = ~n47760 & ~n47763;
  assign n47765 = n47752 & ~n47758;
  assign n47766 = n47751 & n47765;
  assign n47767 = n47764 & ~n47766;
  assign n47768 = n47563 & ~n47767;
  assign n47769 = ~n47563 & n47767;
  assign n47770 = ~n47768 & ~n47769;
  assign n47771 = n47562 & ~n47770;
  assign n47772 = ~n47563 & n47766;
  assign n47773 = ~n47563 & ~n47764;
  assign n47774 = n47563 & ~n47766;
  assign n47775 = n47764 & n47774;
  assign n47776 = ~n47772 & ~n47773;
  assign n47777 = ~n47775 & n47776;
  assign n47778 = ~n47562 & ~n47777;
  assign n47779 = ~n47771 & ~n47778;
  assign n47780 = n47558 & ~n47779;
  assign n47781 = n47500 & n47555;
  assign n47782 = ~n47555 & ~n47556;
  assign n47783 = ~n47500 & n47782;
  assign n47784 = n47555 & n47556;
  assign n47785 = ~n47781 & ~n47783;
  assign n47786 = ~n47784 & n47785;
  assign n47787 = n47779 & ~n47786;
  assign n47788 = ~n47780 & ~n47787;
  assign n47789 = n47555 & n47557;
  assign n47790 = ~n47779 & n47789;
  assign n47791 = n47788 & ~n47790;
  assign n47792 = n47554 & ~n47791;
  assign n47793 = ~n47554 & n47791;
  assign n47794 = ~n47792 & ~n47793;
  assign n47795 = n47553 & ~n47794;
  assign n47796 = ~n47554 & n47790;
  assign n47797 = n47554 & ~n47790;
  assign n47798 = n47788 & n47797;
  assign n47799 = ~n47554 & ~n47788;
  assign n47800 = ~n47796 & ~n47798;
  assign n47801 = ~n47799 & n47800;
  assign n47802 = ~n47553 & ~n47801;
  assign n47803 = ~n47795 & ~n47802;
  assign n47804 = P4_DATAO_REG_6_ & n44378;
  assign n47805 = ~n47287 & ~n47525;
  assign n47806 = ~n47524 & ~n47805;
  assign n47807 = ~n47803 & ~n47804;
  assign n47808 = ~n47806 & n47807;
  assign n47809 = n47803 & n47804;
  assign n47810 = ~n47807 & ~n47809;
  assign n47811 = n47806 & n47810;
  assign n47812 = ~n47808 & ~n47811;
  assign n47813 = n47804 & ~n47806;
  assign n47814 = n47803 & n47813;
  assign n47815 = n47812 & ~n47814;
  assign n47816 = n47548 & ~n47815;
  assign n47817 = ~n47548 & n47815;
  assign n47818 = ~n47816 & ~n47817;
  assign n47819 = ~n47283 & ~n47528;
  assign n47820 = ~n47284 & ~n47533;
  assign n47821 = ~n47819 & n47820;
  assign n47822 = ~n47818 & n47821;
  assign n47823 = ~n47548 & n47814;
  assign n47824 = n47548 & ~n47814;
  assign n47825 = n47812 & n47824;
  assign n47826 = ~n47548 & ~n47812;
  assign n47827 = ~n47823 & ~n47825;
  assign n47828 = ~n47826 & n47827;
  assign n47829 = ~n47821 & ~n47828;
  assign n47830 = ~n47822 & ~n47829;
  assign n47831 = n47279 & ~n47830;
  assign n47832 = ~n47546 & ~n47830;
  assign n47833 = ~n47547 & ~n47831;
  assign n47834 = ~n47832 & n47833;
  assign n47835 = P4_DATAO_REG_4_ & n46777;
  assign n47836 = P4_DATAO_REG_7_ & n44378;
  assign n47837 = ~n47553 & n47554;
  assign n47838 = ~n47553 & n47791;
  assign n47839 = ~n47798 & ~n47837;
  assign n47840 = ~n47838 & n47839;
  assign n47841 = n47836 & ~n47840;
  assign n47842 = ~n47836 & n47840;
  assign n47843 = ~n47841 & ~n47842;
  assign n47844 = n47555 & ~n47779;
  assign n47845 = n47555 & ~n47557;
  assign n47846 = ~n47557 & ~n47779;
  assign n47847 = ~n47844 & ~n47845;
  assign n47848 = ~n47846 & n47847;
  assign n47849 = P4_DATAO_REG_8_ & n44380;
  assign n47850 = ~n47751 & n47752;
  assign n47851 = ~n47751 & ~n47758;
  assign n47852 = ~n47765 & ~n47850;
  assign n47853 = ~n47851 & n47852;
  assign n47854 = P4_DATAO_REG_10_ & n45602;
  assign n47855 = P4_DATAO_REG_11_ & n44384;
  assign n47856 = ~n47566 & n47567;
  assign n47857 = ~n47566 & n47739;
  assign n47858 = ~n47746 & ~n47856;
  assign n47859 = ~n47857 & n47858;
  assign n47860 = P4_DATAO_REG_14_ & n44390;
  assign n47861 = ~n47570 & ~n47702;
  assign n47862 = ~n47705 & ~n47711;
  assign n47863 = ~n47861 & n47862;
  assign n47864 = n47860 & ~n47863;
  assign n47865 = ~n47860 & n47863;
  assign n47866 = ~n47864 & ~n47865;
  assign n47867 = ~n47573 & ~n47699;
  assign n47868 = ~n47698 & ~n47867;
  assign n47869 = n47575 & ~n47682;
  assign n47870 = ~n47578 & ~n47682;
  assign n47871 = ~n47685 & ~n47869;
  assign n47872 = ~n47870 & n47871;
  assign n47873 = P4_DATAO_REG_16_ & n44394;
  assign n47874 = n47584 & ~n47663;
  assign n47875 = ~n47587 & ~n47663;
  assign n47876 = ~n47666 & ~n47874;
  assign n47877 = ~n47875 & n47876;
  assign n47878 = P4_DATAO_REG_18_ & n44623;
  assign n47879 = ~n47640 & ~n47644;
  assign n47880 = ~n47641 & ~n47649;
  assign n47881 = ~n47879 & n47880;
  assign n47882 = P4_DATAO_REG_20_ & n44102;
  assign n47883 = ~n47616 & n47617;
  assign n47884 = ~n47616 & ~n47619;
  assign n47885 = ~n47626 & ~n47883;
  assign n47886 = ~n47884 & n47885;
  assign n47887 = P4_DATAO_REG_22_ & n44143;
  assign n47888 = P4_DATAO_REG_24_ & n44108;
  assign n47889 = P4_DATAO_REG_25_ & n44110;
  assign n47890 = P4_DATAO_REG_26_ & n44112;
  assign n47891 = n47889 & ~n47890;
  assign n47892 = ~n47889 & n47890;
  assign n47893 = ~n47891 & ~n47892;
  assign n47894 = n47888 & ~n47893;
  assign n47895 = ~n47888 & n47893;
  assign n47896 = P4_DATAO_REG_24_ & P4_DATAO_REG_25_;
  assign n47897 = n44119 & n47896;
  assign n47898 = ~n47894 & ~n47895;
  assign n47899 = ~n47897 & n47898;
  assign n47900 = ~n47888 & ~n47891;
  assign n47901 = n47888 & ~n47890;
  assign n47902 = ~n47900 & ~n47901;
  assign n47903 = n47897 & ~n47902;
  assign n47904 = ~n47899 & ~n47903;
  assign n47905 = P4_DATAO_REG_23_ & n44106;
  assign n47906 = ~n47607 & n47609;
  assign n47907 = ~n47606 & ~n47906;
  assign n47908 = ~n47904 & ~n47905;
  assign n47909 = ~n47907 & n47908;
  assign n47910 = n47904 & n47905;
  assign n47911 = ~n47908 & ~n47910;
  assign n47912 = n47907 & n47911;
  assign n47913 = ~n47909 & ~n47912;
  assign n47914 = n47905 & ~n47907;
  assign n47915 = n47904 & n47914;
  assign n47916 = n47913 & ~n47915;
  assign n47917 = n47887 & ~n47916;
  assign n47918 = ~n47887 & n47916;
  assign n47919 = ~n47917 & ~n47918;
  assign n47920 = n47886 & ~n47919;
  assign n47921 = ~n47887 & n47915;
  assign n47922 = ~n47887 & ~n47913;
  assign n47923 = n47887 & n47913;
  assign n47924 = ~n47915 & n47923;
  assign n47925 = ~n47921 & ~n47922;
  assign n47926 = ~n47924 & n47925;
  assign n47927 = ~n47886 & ~n47926;
  assign n47928 = ~n47920 & ~n47927;
  assign n47929 = P4_DATAO_REG_21_ & n44104;
  assign n47930 = ~n47598 & n47599;
  assign n47931 = ~n47598 & n47628;
  assign n47932 = ~n47636 & ~n47930;
  assign n47933 = ~n47931 & n47932;
  assign n47934 = ~n47928 & ~n47929;
  assign n47935 = ~n47933 & n47934;
  assign n47936 = n47928 & n47929;
  assign n47937 = ~n47934 & ~n47936;
  assign n47938 = n47933 & n47937;
  assign n47939 = ~n47935 & ~n47938;
  assign n47940 = n47929 & ~n47933;
  assign n47941 = n47928 & n47940;
  assign n47942 = n47939 & ~n47941;
  assign n47943 = n47882 & ~n47942;
  assign n47944 = ~n47882 & n47942;
  assign n47945 = ~n47943 & ~n47944;
  assign n47946 = n47881 & ~n47945;
  assign n47947 = ~n47882 & n47941;
  assign n47948 = n47882 & ~n47941;
  assign n47949 = n47939 & n47948;
  assign n47950 = ~n47882 & ~n47939;
  assign n47951 = ~n47947 & ~n47949;
  assign n47952 = ~n47950 & n47951;
  assign n47953 = ~n47881 & ~n47952;
  assign n47954 = ~n47946 & ~n47953;
  assign n47955 = P4_DATAO_REG_19_ & n44356;
  assign n47956 = ~n47592 & ~n47660;
  assign n47957 = ~n47659 & ~n47956;
  assign n47958 = ~n47954 & ~n47955;
  assign n47959 = ~n47957 & n47958;
  assign n47960 = n47954 & n47955;
  assign n47961 = ~n47958 & ~n47960;
  assign n47962 = n47957 & n47961;
  assign n47963 = ~n47959 & ~n47962;
  assign n47964 = n47955 & ~n47957;
  assign n47965 = n47954 & n47964;
  assign n47966 = n47963 & ~n47965;
  assign n47967 = n47878 & ~n47966;
  assign n47968 = ~n47878 & n47966;
  assign n47969 = ~n47967 & ~n47968;
  assign n47970 = n47877 & ~n47969;
  assign n47971 = ~n47878 & n47965;
  assign n47972 = n47878 & ~n47965;
  assign n47973 = n47963 & n47972;
  assign n47974 = ~n47878 & ~n47963;
  assign n47975 = ~n47971 & ~n47973;
  assign n47976 = ~n47974 & n47975;
  assign n47977 = ~n47877 & ~n47976;
  assign n47978 = ~n47970 & ~n47977;
  assign n47979 = P4_DATAO_REG_17_ & n44704;
  assign n47980 = ~n47582 & ~n47679;
  assign n47981 = ~n47678 & ~n47980;
  assign n47982 = ~n47978 & ~n47979;
  assign n47983 = ~n47981 & n47982;
  assign n47984 = n47978 & n47979;
  assign n47985 = ~n47982 & ~n47984;
  assign n47986 = n47981 & n47985;
  assign n47987 = ~n47983 & ~n47986;
  assign n47988 = n47979 & ~n47981;
  assign n47989 = n47978 & n47988;
  assign n47990 = n47987 & ~n47989;
  assign n47991 = n47873 & ~n47990;
  assign n47992 = ~n47873 & n47990;
  assign n47993 = ~n47991 & ~n47992;
  assign n47994 = n47872 & ~n47993;
  assign n47995 = ~n47873 & n47989;
  assign n47996 = n47873 & ~n47989;
  assign n47997 = n47987 & n47996;
  assign n47998 = ~n47873 & ~n47987;
  assign n47999 = ~n47995 & ~n47997;
  assign n48000 = ~n47998 & n47999;
  assign n48001 = ~n47872 & ~n48000;
  assign n48002 = ~n47994 & ~n48001;
  assign n48003 = P4_DATAO_REG_15_ & n44392;
  assign n48004 = n47868 & ~n48002;
  assign n48005 = n48003 & n48004;
  assign n48006 = n47868 & n48002;
  assign n48007 = ~n48003 & n48006;
  assign n48008 = ~n48005 & ~n48007;
  assign n48009 = ~n47868 & ~n48003;
  assign n48010 = ~n48002 & n48009;
  assign n48011 = ~n47868 & n48003;
  assign n48012 = n48002 & n48011;
  assign n48013 = ~n48010 & ~n48012;
  assign n48014 = n48008 & n48013;
  assign n48015 = n47866 & ~n48014;
  assign n48016 = ~n47860 & ~n47861;
  assign n48017 = ~n47711 & n48016;
  assign n48018 = ~n47705 & n48017;
  assign n48019 = ~n47864 & ~n48018;
  assign n48020 = n48014 & ~n48019;
  assign n48021 = ~n48015 & ~n48020;
  assign n48022 = P4_DATAO_REG_13_ & n44388;
  assign n48023 = n47713 & ~n47719;
  assign n48024 = ~n47720 & ~n48023;
  assign n48025 = ~n48021 & ~n48022;
  assign n48026 = ~n48024 & n48025;
  assign n48027 = n48021 & n48022;
  assign n48028 = ~n48025 & ~n48027;
  assign n48029 = n48024 & n48028;
  assign n48030 = ~n48026 & ~n48029;
  assign n48031 = n48022 & ~n48024;
  assign n48032 = n48021 & n48031;
  assign n48033 = n48030 & ~n48032;
  assign n48034 = ~n47724 & n47725;
  assign n48035 = ~n47724 & ~n47730;
  assign n48036 = P4_DATAO_REG_12_ & n44386;
  assign n48037 = ~n47737 & ~n48034;
  assign n48038 = ~n48035 & n48037;
  assign n48039 = ~n48036 & n48038;
  assign n48040 = n48036 & ~n48038;
  assign n48041 = ~n48039 & ~n48040;
  assign n48042 = n48033 & ~n48041;
  assign n48043 = ~n48033 & n48041;
  assign n48044 = ~n48042 & ~n48043;
  assign n48045 = ~n47855 & ~n47859;
  assign n48046 = ~n48044 & n48045;
  assign n48047 = n47855 & ~n47859;
  assign n48048 = n48044 & n48047;
  assign n48049 = ~n48046 & ~n48048;
  assign n48050 = n47859 & ~n48044;
  assign n48051 = n47855 & n48050;
  assign n48052 = ~n47857 & n48044;
  assign n48053 = n47858 & n48052;
  assign n48054 = ~n47855 & n48053;
  assign n48055 = ~n48051 & ~n48054;
  assign n48056 = n48049 & n48055;
  assign n48057 = n47854 & ~n48056;
  assign n48058 = ~n47854 & n48056;
  assign n48059 = ~n48057 & ~n48058;
  assign n48060 = n47853 & ~n48059;
  assign n48061 = ~n47854 & ~n48055;
  assign n48062 = ~n47854 & ~n48049;
  assign n48063 = n47854 & n48049;
  assign n48064 = n48055 & n48063;
  assign n48065 = ~n48061 & ~n48062;
  assign n48066 = ~n48064 & n48065;
  assign n48067 = ~n47853 & ~n48066;
  assign n48068 = ~n48060 & ~n48067;
  assign n48069 = P4_DATAO_REG_9_ & n44382;
  assign n48070 = ~n48068 & ~n48069;
  assign n48071 = ~n47563 & ~n47767;
  assign n48072 = ~n47562 & ~n48071;
  assign n48073 = ~n47775 & ~n48072;
  assign n48074 = n48070 & ~n48073;
  assign n48075 = n48068 & n48069;
  assign n48076 = ~n48070 & ~n48075;
  assign n48077 = n48073 & n48076;
  assign n48078 = ~n48074 & ~n48077;
  assign n48079 = n48069 & ~n48073;
  assign n48080 = n48068 & n48079;
  assign n48081 = n48078 & ~n48080;
  assign n48082 = n47849 & ~n48081;
  assign n48083 = ~n47849 & n48081;
  assign n48084 = ~n48082 & ~n48083;
  assign n48085 = n47848 & ~n48084;
  assign n48086 = ~n47849 & n48080;
  assign n48087 = n47849 & ~n48080;
  assign n48088 = n48078 & n48087;
  assign n48089 = ~n47849 & ~n48078;
  assign n48090 = ~n48086 & ~n48088;
  assign n48091 = ~n48089 & n48090;
  assign n48092 = ~n47848 & ~n48091;
  assign n48093 = ~n48085 & ~n48092;
  assign n48094 = ~n47843 & n48093;
  assign n48095 = n47843 & ~n48093;
  assign n48096 = ~n48094 & ~n48095;
  assign n48097 = P4_DATAO_REG_6_ & n44376;
  assign n48098 = ~n48096 & ~n48097;
  assign n48099 = n48096 & n48097;
  assign n48100 = ~n47803 & n47804;
  assign n48101 = ~n47803 & ~n47806;
  assign n48102 = ~n47813 & ~n48100;
  assign n48103 = ~n48101 & n48102;
  assign n48104 = ~n48098 & ~n48099;
  assign n48105 = n48103 & n48104;
  assign n48106 = ~n48103 & ~n48104;
  assign n48107 = ~n48105 & ~n48106;
  assign n48108 = P4_DATAO_REG_5_ & n44374;
  assign n48109 = ~n48107 & ~n48108;
  assign n48110 = n48107 & n48108;
  assign n48111 = ~n47548 & ~n47815;
  assign n48112 = ~n47821 & ~n48111;
  assign n48113 = ~n47825 & ~n48112;
  assign n48114 = ~n48109 & ~n48110;
  assign n48115 = n48113 & n48114;
  assign n48116 = n48109 & ~n48113;
  assign n48117 = n48108 & ~n48113;
  assign n48118 = n48107 & n48117;
  assign n48119 = ~n48115 & ~n48116;
  assign n48120 = ~n48118 & n48119;
  assign n48121 = n47835 & ~n48120;
  assign n48122 = ~n47835 & n48120;
  assign n48123 = ~n48121 & ~n48122;
  assign n48124 = n47834 & ~n48123;
  assign n48125 = n47835 & n48120;
  assign n48126 = ~n47835 & ~n48120;
  assign n48127 = ~n48125 & ~n48126;
  assign n48128 = ~n47834 & ~n48127;
  assign n48129 = ~n48124 & ~n48128;
  assign n48130 = P4_DATAO_REG_3_ & n44372;
  assign n48131 = n48129 & n48130;
  assign n48132 = ~n48129 & ~n48130;
  assign n48133 = ~n48131 & ~n48132;
  assign n48134 = P4_DATAO_REG_3_ & n46777;
  assign n48135 = P4_DATAO_REG_3_ & n44374;
  assign n48136 = ~n47048 & ~n47053;
  assign n48137 = ~n47049 & ~n48136;
  assign n48138 = n48135 & ~n48137;
  assign n48139 = n47280 & ~n47539;
  assign n48140 = ~n47280 & n47539;
  assign n48141 = ~n48139 & ~n48140;
  assign n48142 = n47544 & ~n48141;
  assign n48143 = ~n47538 & ~n47540;
  assign n48144 = ~n47544 & ~n48143;
  assign n48145 = ~n48142 & ~n48144;
  assign n48146 = n48135 & ~n48145;
  assign n48147 = ~n48137 & ~n48145;
  assign n48148 = ~n48138 & ~n48146;
  assign n48149 = ~n48147 & n48148;
  assign n48150 = n48134 & ~n48149;
  assign n48151 = n47547 & n47830;
  assign n48152 = n48134 & ~n48151;
  assign n48153 = ~n47279 & ~n47830;
  assign n48154 = ~n47546 & n48153;
  assign n48155 = n47279 & n47830;
  assign n48156 = ~n48153 & ~n48155;
  assign n48157 = n47546 & n48156;
  assign n48158 = ~n48154 & ~n48157;
  assign n48159 = n48152 & n48158;
  assign n48160 = ~n48151 & n48158;
  assign n48161 = ~n48149 & n48160;
  assign n48162 = ~n48150 & ~n48159;
  assign n48163 = ~n48161 & n48162;
  assign n48164 = ~n48133 & ~n48163;
  assign n48165 = n48133 & n48163;
  assign n48166 = ~n48164 & ~n48165;
  assign n48167 = n47278 & n48166;
  assign n48168 = ~n47278 & ~n48166;
  assign n48169 = P4_DATAO_REG_2_ & n44372;
  assign n48170 = P4_DATAO_REG_2_ & n46777;
  assign n48171 = ~n48135 & n48137;
  assign n48172 = ~n48138 & ~n48171;
  assign n48173 = n48145 & ~n48172;
  assign n48174 = ~n48145 & n48172;
  assign n48175 = ~n48173 & ~n48174;
  assign n48176 = n48170 & n48175;
  assign n48177 = ~n48170 & ~n48175;
  assign n48178 = ~n47057 & ~n47060;
  assign n48179 = ~n47063 & ~n47068;
  assign n48180 = ~n48178 & n48179;
  assign n48181 = ~n48177 & ~n48180;
  assign n48182 = ~n48176 & ~n48181;
  assign n48183 = n48169 & ~n48182;
  assign n48184 = n48134 & ~n48160;
  assign n48185 = ~n48134 & n48160;
  assign n48186 = ~n48184 & ~n48185;
  assign n48187 = n48149 & ~n48186;
  assign n48188 = ~n48134 & n48151;
  assign n48189 = ~n48134 & ~n48158;
  assign n48190 = ~n48159 & ~n48188;
  assign n48191 = ~n48189 & n48190;
  assign n48192 = ~n48149 & ~n48191;
  assign n48193 = ~n48187 & ~n48192;
  assign n48194 = n48169 & ~n48193;
  assign n48195 = ~n48182 & ~n48193;
  assign n48196 = ~n48183 & ~n48194;
  assign n48197 = ~n48195 & n48196;
  assign n48198 = ~n48168 & ~n48197;
  assign n48199 = ~n48167 & ~n48198;
  assign n48200 = n47276 & ~n48199;
  assign n48201 = ~n48129 & n48130;
  assign n48202 = n48129 & ~n48130;
  assign n48203 = ~n48163 & ~n48202;
  assign n48204 = ~n48201 & ~n48203;
  assign n48205 = P4_DATAO_REG_3_ & n47277;
  assign n48206 = P4_DATAO_REG_4_ & n44372;
  assign n48207 = ~n47834 & ~n48126;
  assign n48208 = ~n48125 & ~n48207;
  assign n48209 = ~n44374 & ~n44376;
  assign n48210 = ~n47815 & n48209;
  assign n48211 = n47821 & ~n48108;
  assign n48212 = ~n47825 & n48211;
  assign n48213 = ~n48107 & ~n48210;
  assign n48214 = ~n48212 & n48213;
  assign n48215 = ~n48117 & ~n48214;
  assign n48216 = P4_DATAO_REG_5_ & n46777;
  assign n48217 = n47836 & ~n48093;
  assign n48218 = ~n47840 & ~n48093;
  assign n48219 = ~n47841 & ~n48217;
  assign n48220 = ~n48218 & n48219;
  assign n48221 = P4_DATAO_REG_7_ & n44376;
  assign n48222 = ~n48068 & n48069;
  assign n48223 = ~n48068 & ~n48073;
  assign n48224 = ~n48079 & ~n48222;
  assign n48225 = ~n48223 & n48224;
  assign n48226 = P4_DATAO_REG_9_ & n44380;
  assign n48227 = P4_DATAO_REG_12_ & n44384;
  assign n48228 = ~n48035 & ~n48036;
  assign n48229 = ~n47737 & n48228;
  assign n48230 = ~n48034 & n48229;
  assign n48231 = n48033 & ~n48230;
  assign n48232 = ~n48040 & ~n48231;
  assign n48233 = P4_DATAO_REG_13_ & n44386;
  assign n48234 = ~n48021 & n48022;
  assign n48235 = ~n48021 & ~n48024;
  assign n48236 = ~n48031 & ~n48234;
  assign n48237 = ~n48235 & n48236;
  assign n48238 = n48233 & ~n48237;
  assign n48239 = ~n48233 & n48237;
  assign n48240 = ~n48238 & ~n48239;
  assign n48241 = ~n48002 & n48003;
  assign n48242 = ~n47868 & ~n48002;
  assign n48243 = ~n48011 & ~n48241;
  assign n48244 = ~n48242 & n48243;
  assign n48245 = P4_DATAO_REG_15_ & n44390;
  assign n48246 = ~n47978 & n47979;
  assign n48247 = ~n47978 & ~n47981;
  assign n48248 = ~n47988 & ~n48246;
  assign n48249 = ~n48247 & n48248;
  assign n48250 = P4_DATAO_REG_17_ & n44394;
  assign n48251 = ~n47928 & n47929;
  assign n48252 = ~n47928 & ~n47933;
  assign n48253 = ~n47940 & ~n48251;
  assign n48254 = ~n48252 & n48253;
  assign n48255 = P4_DATAO_REG_21_ & n44102;
  assign n48256 = P4_DATAO_REG_22_ & n44104;
  assign n48257 = ~n47886 & n47887;
  assign n48258 = ~n47886 & n47916;
  assign n48259 = ~n47924 & ~n48257;
  assign n48260 = ~n48258 & n48259;
  assign n48261 = ~n48256 & ~n48260;
  assign n48262 = ~n47904 & n47905;
  assign n48263 = ~n47904 & ~n47907;
  assign n48264 = ~n47914 & ~n48262;
  assign n48265 = ~n48263 & n48264;
  assign n48266 = P4_DATAO_REG_23_ & n44143;
  assign n48267 = P4_DATAO_REG_25_ & n44108;
  assign n48268 = P4_DATAO_REG_26_ & n44110;
  assign n48269 = P4_DATAO_REG_27_ & n44112;
  assign n48270 = n48268 & ~n48269;
  assign n48271 = ~n48268 & n48269;
  assign n48272 = ~n48270 & ~n48271;
  assign n48273 = n48267 & ~n48272;
  assign n48274 = ~n48267 & n48272;
  assign n48275 = P4_DATAO_REG_25_ & P4_DATAO_REG_26_;
  assign n48276 = n44119 & n48275;
  assign n48277 = ~n48273 & ~n48274;
  assign n48278 = ~n48276 & n48277;
  assign n48279 = n48267 & ~n48270;
  assign n48280 = ~n48267 & n48270;
  assign n48281 = ~n48279 & ~n48280;
  assign n48282 = n48276 & n48281;
  assign n48283 = ~n48278 & ~n48282;
  assign n48284 = P4_DATAO_REG_24_ & n44106;
  assign n48285 = ~n47895 & n47897;
  assign n48286 = ~n47894 & ~n48285;
  assign n48287 = ~n48283 & ~n48284;
  assign n48288 = ~n48286 & n48287;
  assign n48289 = n48283 & n48284;
  assign n48290 = ~n48287 & ~n48289;
  assign n48291 = n48286 & n48290;
  assign n48292 = ~n48288 & ~n48291;
  assign n48293 = n48284 & ~n48286;
  assign n48294 = n48283 & n48293;
  assign n48295 = n48292 & ~n48294;
  assign n48296 = n48266 & ~n48295;
  assign n48297 = ~n48266 & n48295;
  assign n48298 = ~n48296 & ~n48297;
  assign n48299 = n48265 & ~n48298;
  assign n48300 = ~n48266 & n48294;
  assign n48301 = ~n48266 & ~n48292;
  assign n48302 = n48266 & n48292;
  assign n48303 = ~n48294 & n48302;
  assign n48304 = ~n48300 & ~n48301;
  assign n48305 = ~n48303 & n48304;
  assign n48306 = ~n48265 & ~n48305;
  assign n48307 = ~n48299 & ~n48306;
  assign n48308 = n48261 & ~n48307;
  assign n48309 = n48256 & ~n48260;
  assign n48310 = n48307 & n48309;
  assign n48311 = ~n48308 & ~n48310;
  assign n48312 = n48260 & ~n48307;
  assign n48313 = n48256 & n48312;
  assign n48314 = n48260 & n48307;
  assign n48315 = ~n48256 & n48314;
  assign n48316 = ~n48313 & ~n48315;
  assign n48317 = n48311 & n48316;
  assign n48318 = n48255 & ~n48317;
  assign n48319 = ~n48255 & n48317;
  assign n48320 = ~n48318 & ~n48319;
  assign n48321 = n48254 & ~n48320;
  assign n48322 = ~n48255 & ~n48311;
  assign n48323 = n48255 & n48311;
  assign n48324 = n48316 & n48323;
  assign n48325 = ~n48255 & ~n48316;
  assign n48326 = ~n48322 & ~n48324;
  assign n48327 = ~n48325 & n48326;
  assign n48328 = ~n48254 & ~n48327;
  assign n48329 = ~n48321 & ~n48328;
  assign n48330 = P4_DATAO_REG_20_ & n44356;
  assign n48331 = ~n47882 & ~n47942;
  assign n48332 = ~n47881 & ~n48331;
  assign n48333 = ~n47949 & ~n48332;
  assign n48334 = ~n48329 & ~n48330;
  assign n48335 = ~n48333 & n48334;
  assign n48336 = n48329 & n48330;
  assign n48337 = ~n48334 & ~n48336;
  assign n48338 = n48333 & n48337;
  assign n48339 = ~n48335 & ~n48338;
  assign n48340 = n48330 & ~n48333;
  assign n48341 = n48329 & n48340;
  assign n48342 = n48339 & ~n48341;
  assign n48343 = ~n47954 & n47955;
  assign n48344 = ~n47954 & ~n47957;
  assign n48345 = P4_DATAO_REG_19_ & n44623;
  assign n48346 = ~n47964 & ~n48343;
  assign n48347 = ~n48344 & n48346;
  assign n48348 = ~n48345 & n48347;
  assign n48349 = n48345 & ~n48347;
  assign n48350 = ~n48348 & ~n48349;
  assign n48351 = n48342 & ~n48350;
  assign n48352 = ~n48342 & n48350;
  assign n48353 = ~n48351 & ~n48352;
  assign n48354 = P4_DATAO_REG_18_ & n44704;
  assign n48355 = ~n48353 & ~n48354;
  assign n48356 = ~n47878 & ~n47966;
  assign n48357 = ~n47877 & ~n48356;
  assign n48358 = ~n47973 & ~n48357;
  assign n48359 = n48355 & ~n48358;
  assign n48360 = n48353 & n48354;
  assign n48361 = ~n48355 & ~n48360;
  assign n48362 = n48358 & n48361;
  assign n48363 = ~n48359 & ~n48362;
  assign n48364 = n48354 & ~n48358;
  assign n48365 = n48353 & n48364;
  assign n48366 = n48363 & ~n48365;
  assign n48367 = n48250 & ~n48366;
  assign n48368 = ~n48250 & n48366;
  assign n48369 = ~n48367 & ~n48368;
  assign n48370 = n48249 & ~n48369;
  assign n48371 = n48250 & ~n48365;
  assign n48372 = n48363 & n48371;
  assign n48373 = ~n48250 & ~n48366;
  assign n48374 = ~n48372 & ~n48373;
  assign n48375 = ~n48249 & ~n48374;
  assign n48376 = ~n48370 & ~n48375;
  assign n48377 = P4_DATAO_REG_16_ & n44392;
  assign n48378 = ~n48376 & ~n48377;
  assign n48379 = ~n47873 & ~n47990;
  assign n48380 = ~n47872 & ~n48379;
  assign n48381 = ~n47997 & ~n48380;
  assign n48382 = n48378 & ~n48381;
  assign n48383 = ~n48376 & n48377;
  assign n48384 = n48376 & ~n48377;
  assign n48385 = ~n48383 & ~n48384;
  assign n48386 = n48381 & ~n48385;
  assign n48387 = ~n48382 & ~n48386;
  assign n48388 = n48377 & ~n48381;
  assign n48389 = n48376 & n48388;
  assign n48390 = n48387 & ~n48389;
  assign n48391 = n48245 & ~n48390;
  assign n48392 = ~n48245 & n48390;
  assign n48393 = ~n48391 & ~n48392;
  assign n48394 = n48244 & ~n48393;
  assign n48395 = n48245 & ~n48389;
  assign n48396 = n48387 & n48395;
  assign n48397 = ~n48245 & ~n48390;
  assign n48398 = ~n48396 & ~n48397;
  assign n48399 = ~n48244 & ~n48398;
  assign n48400 = ~n48394 & ~n48399;
  assign n48401 = ~n47865 & n48014;
  assign n48402 = ~n47864 & ~n48401;
  assign n48403 = P4_DATAO_REG_14_ & n44388;
  assign n48404 = ~n48400 & ~n48402;
  assign n48405 = ~n48403 & n48404;
  assign n48406 = ~n48400 & n48402;
  assign n48407 = n48403 & n48406;
  assign n48408 = ~n48402 & n48403;
  assign n48409 = n48402 & ~n48403;
  assign n48410 = ~n48408 & ~n48409;
  assign n48411 = n48400 & ~n48410;
  assign n48412 = ~n48405 & ~n48407;
  assign n48413 = ~n48411 & n48412;
  assign n48414 = n48240 & ~n48413;
  assign n48415 = ~n48240 & n48413;
  assign n48416 = ~n48414 & ~n48415;
  assign n48417 = ~n48227 & ~n48232;
  assign n48418 = ~n48416 & n48417;
  assign n48419 = n48227 & ~n48232;
  assign n48420 = ~n48227 & n48232;
  assign n48421 = ~n48419 & ~n48420;
  assign n48422 = n48416 & ~n48421;
  assign n48423 = ~n48418 & ~n48422;
  assign n48424 = n48227 & n48232;
  assign n48425 = ~n48416 & n48424;
  assign n48426 = n48423 & ~n48425;
  assign n48427 = n47855 & ~n48044;
  assign n48428 = ~n47859 & ~n48044;
  assign n48429 = P4_DATAO_REG_11_ & n45602;
  assign n48430 = ~n48047 & ~n48427;
  assign n48431 = ~n48428 & n48430;
  assign n48432 = ~n48429 & n48431;
  assign n48433 = n48429 & ~n48431;
  assign n48434 = ~n48432 & ~n48433;
  assign n48435 = n48426 & ~n48434;
  assign n48436 = ~n48426 & n48434;
  assign n48437 = ~n48435 & ~n48436;
  assign n48438 = P4_DATAO_REG_10_ & n44382;
  assign n48439 = ~n47853 & n48065;
  assign n48440 = ~n48064 & ~n48439;
  assign n48441 = ~n48437 & ~n48438;
  assign n48442 = ~n48440 & n48441;
  assign n48443 = n48437 & n48438;
  assign n48444 = ~n48441 & ~n48443;
  assign n48445 = n48440 & n48444;
  assign n48446 = ~n48442 & ~n48445;
  assign n48447 = ~n48440 & n48443;
  assign n48448 = n48446 & ~n48447;
  assign n48449 = n48226 & ~n48448;
  assign n48450 = ~n48226 & n48448;
  assign n48451 = ~n48449 & ~n48450;
  assign n48452 = n48225 & ~n48451;
  assign n48453 = ~n48226 & n48447;
  assign n48454 = ~n48226 & ~n48446;
  assign n48455 = n48226 & ~n48447;
  assign n48456 = n48446 & n48455;
  assign n48457 = ~n48453 & ~n48454;
  assign n48458 = ~n48456 & n48457;
  assign n48459 = ~n48225 & ~n48458;
  assign n48460 = ~n48452 & ~n48459;
  assign n48461 = P4_DATAO_REG_8_ & n44378;
  assign n48462 = ~n47849 & ~n48081;
  assign n48463 = ~n47848 & ~n48462;
  assign n48464 = ~n48088 & ~n48463;
  assign n48465 = ~n48460 & ~n48461;
  assign n48466 = ~n48464 & n48465;
  assign n48467 = n48460 & n48461;
  assign n48468 = ~n48465 & ~n48467;
  assign n48469 = n48464 & n48468;
  assign n48470 = ~n48466 & ~n48469;
  assign n48471 = n48461 & ~n48464;
  assign n48472 = n48460 & n48471;
  assign n48473 = n48470 & ~n48472;
  assign n48474 = n48221 & ~n48473;
  assign n48475 = ~n48221 & n48473;
  assign n48476 = ~n48474 & ~n48475;
  assign n48477 = n48220 & ~n48476;
  assign n48478 = ~n48221 & ~n48473;
  assign n48479 = n48221 & ~n48472;
  assign n48480 = n48470 & n48479;
  assign n48481 = ~n48478 & ~n48480;
  assign n48482 = ~n48220 & ~n48481;
  assign n48483 = ~n48477 & ~n48482;
  assign n48484 = P4_DATAO_REG_6_ & n44374;
  assign n48485 = ~n48098 & ~n48103;
  assign n48486 = ~n48099 & ~n48485;
  assign n48487 = ~n48483 & ~n48484;
  assign n48488 = ~n48486 & n48487;
  assign n48489 = n48483 & n48484;
  assign n48490 = ~n48487 & ~n48489;
  assign n48491 = n48486 & n48490;
  assign n48492 = ~n48488 & ~n48491;
  assign n48493 = n48484 & ~n48486;
  assign n48494 = n48483 & n48493;
  assign n48495 = n48492 & ~n48494;
  assign n48496 = n48216 & ~n48495;
  assign n48497 = ~n48216 & n48495;
  assign n48498 = ~n48496 & ~n48497;
  assign n48499 = n48215 & ~n48498;
  assign n48500 = n48216 & n48492;
  assign n48501 = ~n48494 & n48500;
  assign n48502 = ~n48216 & ~n48495;
  assign n48503 = ~n48501 & ~n48502;
  assign n48504 = ~n48215 & ~n48503;
  assign n48505 = ~n48499 & ~n48504;
  assign n48506 = ~n48206 & ~n48208;
  assign n48507 = ~n48505 & n48506;
  assign n48508 = n48206 & ~n48208;
  assign n48509 = n48505 & n48508;
  assign n48510 = ~n48507 & ~n48509;
  assign n48511 = n48208 & ~n48505;
  assign n48512 = n48206 & n48511;
  assign n48513 = n48208 & n48505;
  assign n48514 = ~n48206 & n48513;
  assign n48515 = ~n48512 & ~n48514;
  assign n48516 = n48510 & n48515;
  assign n48517 = n48205 & ~n48516;
  assign n48518 = ~n48205 & n48516;
  assign n48519 = ~n48517 & ~n48518;
  assign n48520 = n48204 & ~n48519;
  assign n48521 = ~n48205 & ~n48515;
  assign n48522 = ~n48205 & ~n48510;
  assign n48523 = n48205 & n48510;
  assign n48524 = n48515 & n48523;
  assign n48525 = ~n48521 & ~n48522;
  assign n48526 = ~n48524 & n48525;
  assign n48527 = ~n48204 & ~n48526;
  assign n48528 = ~n48520 & ~n48527;
  assign n48529 = n47276 & ~n48528;
  assign n48530 = ~n48199 & ~n48528;
  assign n48531 = ~n48200 & ~n48529;
  assign n48532 = ~n48530 & n48531;
  assign n48533 = n47274 & ~n48532;
  assign n48534 = P4_DATAO_REG_3_ & n47275;
  assign n48535 = ~n48205 & ~n48516;
  assign n48536 = ~n48204 & ~n48535;
  assign n48537 = ~n48524 & ~n48536;
  assign n48538 = n48534 & ~n48537;
  assign n48539 = n48206 & ~n48505;
  assign n48540 = ~n48208 & ~n48505;
  assign n48541 = ~n48508 & ~n48539;
  assign n48542 = ~n48540 & n48541;
  assign n48543 = P4_DATAO_REG_4_ & n47277;
  assign n48544 = ~n48483 & n48484;
  assign n48545 = ~n48483 & ~n48486;
  assign n48546 = ~n48493 & ~n48544;
  assign n48547 = ~n48545 & n48546;
  assign n48548 = P4_DATAO_REG_6_ & n46777;
  assign n48549 = P4_DATAO_REG_7_ & n44374;
  assign n48550 = ~n48220 & n48221;
  assign n48551 = ~n48220 & n48473;
  assign n48552 = ~n48480 & ~n48550;
  assign n48553 = ~n48551 & n48552;
  assign n48554 = ~n48549 & ~n48553;
  assign n48555 = ~n48460 & n48461;
  assign n48556 = ~n48460 & ~n48464;
  assign n48557 = ~n48471 & ~n48555;
  assign n48558 = ~n48556 & n48557;
  assign n48559 = P4_DATAO_REG_8_ & n44376;
  assign n48560 = ~n48428 & ~n48429;
  assign n48561 = ~n48047 & n48560;
  assign n48562 = ~n48427 & n48561;
  assign n48563 = n48426 & ~n48562;
  assign n48564 = ~n48433 & ~n48563;
  assign n48565 = P4_DATAO_REG_11_ & n44382;
  assign n48566 = n48564 & n48565;
  assign n48567 = P4_DATAO_REG_12_ & n45602;
  assign n48568 = n48227 & ~n48416;
  assign n48569 = ~n48232 & ~n48416;
  assign n48570 = ~n48419 & ~n48568;
  assign n48571 = ~n48569 & n48570;
  assign n48572 = n48567 & ~n48571;
  assign n48573 = ~n48567 & n48571;
  assign n48574 = ~n48572 & ~n48573;
  assign n48575 = ~n48400 & n48403;
  assign n48576 = ~n48408 & ~n48575;
  assign n48577 = ~n48404 & n48576;
  assign n48578 = P4_DATAO_REG_14_ & n44386;
  assign n48579 = ~n48376 & ~n48381;
  assign n48580 = ~n48383 & ~n48388;
  assign n48581 = ~n48579 & n48580;
  assign n48582 = P4_DATAO_REG_16_ & n44390;
  assign n48583 = ~n48353 & n48354;
  assign n48584 = ~n48353 & ~n48358;
  assign n48585 = ~n48364 & ~n48583;
  assign n48586 = ~n48584 & n48585;
  assign n48587 = P4_DATAO_REG_18_ & n44394;
  assign n48588 = ~n48329 & n48330;
  assign n48589 = ~n48329 & ~n48333;
  assign n48590 = ~n48340 & ~n48588;
  assign n48591 = ~n48589 & n48590;
  assign n48592 = P4_DATAO_REG_20_ & n44623;
  assign n48593 = P4_DATAO_REG_21_ & n44356;
  assign n48594 = ~n48254 & ~n48322;
  assign n48595 = ~n48325 & n48594;
  assign n48596 = ~n48324 & ~n48595;
  assign n48597 = ~n48593 & ~n48596;
  assign n48598 = n48256 & ~n48307;
  assign n48599 = ~n48260 & ~n48307;
  assign n48600 = ~n48309 & ~n48598;
  assign n48601 = ~n48599 & n48600;
  assign n48602 = P4_DATAO_REG_22_ & n44102;
  assign n48603 = P4_DATAO_REG_23_ & n44104;
  assign n48604 = ~n48283 & n48284;
  assign n48605 = ~n48283 & ~n48286;
  assign n48606 = ~n48293 & ~n48604;
  assign n48607 = ~n48605 & n48606;
  assign n48608 = P4_DATAO_REG_24_ & n44143;
  assign n48609 = P4_DATAO_REG_25_ & n44106;
  assign n48610 = ~n48274 & n48276;
  assign n48611 = ~n48273 & ~n48610;
  assign n48612 = ~n48609 & ~n48611;
  assign n48613 = P4_DATAO_REG_26_ & n44108;
  assign n48614 = P4_DATAO_REG_27_ & n44110;
  assign n48615 = P4_DATAO_REG_28_ & n44112;
  assign n48616 = n48614 & ~n48615;
  assign n48617 = ~n48614 & n48615;
  assign n48618 = ~n48616 & ~n48617;
  assign n48619 = n48613 & ~n48618;
  assign n48620 = ~n48613 & n48618;
  assign n48621 = P4_DATAO_REG_26_ & P4_DATAO_REG_27_;
  assign n48622 = n44119 & n48621;
  assign n48623 = ~n48619 & ~n48620;
  assign n48624 = ~n48622 & n48623;
  assign n48625 = ~n48613 & ~n48616;
  assign n48626 = ~n48619 & ~n48625;
  assign n48627 = n48622 & ~n48626;
  assign n48628 = ~n48624 & ~n48627;
  assign n48629 = n48612 & ~n48628;
  assign n48630 = n48609 & ~n48611;
  assign n48631 = n48628 & n48630;
  assign n48632 = n48611 & ~n48628;
  assign n48633 = n48609 & n48632;
  assign n48634 = n48611 & n48628;
  assign n48635 = ~n48609 & n48634;
  assign n48636 = ~n48629 & ~n48631;
  assign n48637 = ~n48633 & n48636;
  assign n48638 = ~n48635 & n48637;
  assign n48639 = n48608 & ~n48638;
  assign n48640 = ~n48608 & n48638;
  assign n48641 = ~n48639 & ~n48640;
  assign n48642 = n48607 & ~n48641;
  assign n48643 = n48608 & n48638;
  assign n48644 = ~n48608 & ~n48638;
  assign n48645 = ~n48643 & ~n48644;
  assign n48646 = ~n48607 & ~n48645;
  assign n48647 = ~n48642 & ~n48646;
  assign n48648 = n48603 & ~n48647;
  assign n48649 = ~n48266 & ~n48295;
  assign n48650 = ~n48265 & ~n48649;
  assign n48651 = ~n48303 & ~n48650;
  assign n48652 = n48648 & n48651;
  assign n48653 = ~n48603 & ~n48647;
  assign n48654 = ~n48651 & n48653;
  assign n48655 = ~n48652 & ~n48654;
  assign n48656 = n48603 & ~n48651;
  assign n48657 = ~n48303 & ~n48603;
  assign n48658 = ~n48650 & n48657;
  assign n48659 = ~n48656 & ~n48658;
  assign n48660 = n48647 & ~n48659;
  assign n48661 = n48655 & ~n48660;
  assign n48662 = n48602 & ~n48661;
  assign n48663 = ~n48602 & n48661;
  assign n48664 = ~n48662 & ~n48663;
  assign n48665 = n48601 & ~n48664;
  assign n48666 = n48602 & ~n48660;
  assign n48667 = n48655 & n48666;
  assign n48668 = ~n48602 & ~n48661;
  assign n48669 = ~n48667 & ~n48668;
  assign n48670 = ~n48601 & ~n48669;
  assign n48671 = ~n48665 & ~n48670;
  assign n48672 = n48597 & ~n48671;
  assign n48673 = n48593 & n48595;
  assign n48674 = ~n48593 & n48596;
  assign n48675 = n48324 & n48593;
  assign n48676 = ~n48673 & ~n48674;
  assign n48677 = ~n48675 & n48676;
  assign n48678 = n48671 & ~n48677;
  assign n48679 = ~n48672 & ~n48678;
  assign n48680 = n48593 & n48596;
  assign n48681 = ~n48671 & n48680;
  assign n48682 = n48679 & ~n48681;
  assign n48683 = n48592 & ~n48682;
  assign n48684 = ~n48592 & n48682;
  assign n48685 = ~n48683 & ~n48684;
  assign n48686 = n48591 & ~n48685;
  assign n48687 = ~n48592 & n48681;
  assign n48688 = n48592 & ~n48681;
  assign n48689 = n48679 & n48688;
  assign n48690 = ~n48592 & ~n48679;
  assign n48691 = ~n48687 & ~n48689;
  assign n48692 = ~n48690 & n48691;
  assign n48693 = ~n48591 & ~n48692;
  assign n48694 = ~n48686 & ~n48693;
  assign n48695 = P4_DATAO_REG_19_ & n44704;
  assign n48696 = n48342 & ~n48348;
  assign n48697 = ~n48349 & ~n48696;
  assign n48698 = ~n48694 & ~n48695;
  assign n48699 = ~n48697 & n48698;
  assign n48700 = n48694 & n48695;
  assign n48701 = ~n48698 & ~n48700;
  assign n48702 = n48697 & n48701;
  assign n48703 = ~n48699 & ~n48702;
  assign n48704 = n48695 & ~n48697;
  assign n48705 = n48694 & n48704;
  assign n48706 = n48703 & ~n48705;
  assign n48707 = n48587 & ~n48706;
  assign n48708 = ~n48587 & n48706;
  assign n48709 = ~n48707 & ~n48708;
  assign n48710 = n48586 & ~n48709;
  assign n48711 = ~n48587 & n48705;
  assign n48712 = n48587 & ~n48705;
  assign n48713 = n48703 & n48712;
  assign n48714 = ~n48587 & ~n48703;
  assign n48715 = ~n48711 & ~n48713;
  assign n48716 = ~n48714 & n48715;
  assign n48717 = ~n48586 & ~n48716;
  assign n48718 = ~n48710 & ~n48717;
  assign n48719 = P4_DATAO_REG_17_ & n44392;
  assign n48720 = ~n48249 & ~n48373;
  assign n48721 = ~n48372 & ~n48720;
  assign n48722 = ~n48718 & ~n48719;
  assign n48723 = ~n48721 & n48722;
  assign n48724 = n48718 & n48719;
  assign n48725 = ~n48722 & ~n48724;
  assign n48726 = n48721 & n48725;
  assign n48727 = ~n48723 & ~n48726;
  assign n48728 = n48719 & ~n48721;
  assign n48729 = n48718 & n48728;
  assign n48730 = n48727 & ~n48729;
  assign n48731 = n48582 & ~n48730;
  assign n48732 = ~n48582 & n48730;
  assign n48733 = ~n48731 & ~n48732;
  assign n48734 = n48581 & ~n48733;
  assign n48735 = ~n48582 & n48729;
  assign n48736 = n48582 & ~n48729;
  assign n48737 = n48727 & n48736;
  assign n48738 = ~n48582 & ~n48727;
  assign n48739 = ~n48735 & ~n48737;
  assign n48740 = ~n48738 & n48739;
  assign n48741 = ~n48581 & ~n48740;
  assign n48742 = ~n48734 & ~n48741;
  assign n48743 = P4_DATAO_REG_15_ & n44388;
  assign n48744 = ~n48244 & ~n48397;
  assign n48745 = ~n48396 & ~n48744;
  assign n48746 = ~n48742 & ~n48743;
  assign n48747 = ~n48745 & n48746;
  assign n48748 = n48742 & n48743;
  assign n48749 = ~n48746 & ~n48748;
  assign n48750 = n48745 & n48749;
  assign n48751 = ~n48747 & ~n48750;
  assign n48752 = n48743 & ~n48745;
  assign n48753 = n48742 & n48752;
  assign n48754 = n48751 & ~n48753;
  assign n48755 = n48578 & ~n48754;
  assign n48756 = ~n48578 & n48754;
  assign n48757 = ~n48755 & ~n48756;
  assign n48758 = n48577 & ~n48757;
  assign n48759 = ~n48578 & n48753;
  assign n48760 = n48578 & ~n48753;
  assign n48761 = n48751 & n48760;
  assign n48762 = ~n48578 & ~n48751;
  assign n48763 = ~n48759 & ~n48761;
  assign n48764 = ~n48762 & n48763;
  assign n48765 = ~n48577 & ~n48764;
  assign n48766 = ~n48758 & ~n48765;
  assign n48767 = P4_DATAO_REG_13_ & n44384;
  assign n48768 = ~n48239 & n48413;
  assign n48769 = ~n48238 & ~n48768;
  assign n48770 = ~n48766 & ~n48767;
  assign n48771 = ~n48769 & n48770;
  assign n48772 = n48766 & n48767;
  assign n48773 = ~n48770 & ~n48772;
  assign n48774 = n48769 & n48773;
  assign n48775 = ~n48771 & ~n48774;
  assign n48776 = n48767 & ~n48769;
  assign n48777 = n48766 & n48776;
  assign n48778 = n48775 & ~n48777;
  assign n48779 = n48574 & ~n48778;
  assign n48780 = ~n48567 & ~n48569;
  assign n48781 = ~n48568 & n48780;
  assign n48782 = ~n48419 & n48781;
  assign n48783 = ~n48572 & ~n48782;
  assign n48784 = n48778 & ~n48783;
  assign n48785 = ~n48779 & ~n48784;
  assign n48786 = n48566 & ~n48785;
  assign n48787 = ~n48564 & n48565;
  assign n48788 = n48564 & ~n48565;
  assign n48789 = ~n48787 & ~n48788;
  assign n48790 = n48785 & ~n48789;
  assign n48791 = ~n48786 & ~n48790;
  assign n48792 = ~n48564 & ~n48565;
  assign n48793 = ~n48785 & n48792;
  assign n48794 = n48791 & ~n48793;
  assign n48795 = n48438 & ~n48440;
  assign n48796 = ~n48437 & n48438;
  assign n48797 = ~n48437 & ~n48440;
  assign n48798 = P4_DATAO_REG_10_ & n44380;
  assign n48799 = ~n48795 & ~n48796;
  assign n48800 = ~n48797 & n48799;
  assign n48801 = ~n48798 & n48800;
  assign n48802 = n48798 & ~n48800;
  assign n48803 = ~n48801 & ~n48802;
  assign n48804 = n48794 & ~n48803;
  assign n48805 = ~n48794 & n48803;
  assign n48806 = ~n48804 & ~n48805;
  assign n48807 = P4_DATAO_REG_9_ & n44378;
  assign n48808 = ~n48226 & ~n48448;
  assign n48809 = ~n48225 & ~n48808;
  assign n48810 = ~n48456 & ~n48809;
  assign n48811 = ~n48806 & ~n48807;
  assign n48812 = ~n48810 & n48811;
  assign n48813 = n48806 & n48807;
  assign n48814 = ~n48811 & ~n48813;
  assign n48815 = n48810 & n48814;
  assign n48816 = ~n48812 & ~n48815;
  assign n48817 = ~n48810 & n48813;
  assign n48818 = n48816 & ~n48817;
  assign n48819 = n48559 & ~n48818;
  assign n48820 = ~n48559 & n48818;
  assign n48821 = ~n48819 & ~n48820;
  assign n48822 = n48558 & ~n48821;
  assign n48823 = ~n48559 & n48817;
  assign n48824 = ~n48559 & ~n48816;
  assign n48825 = n48559 & ~n48817;
  assign n48826 = n48816 & n48825;
  assign n48827 = ~n48823 & ~n48824;
  assign n48828 = ~n48826 & n48827;
  assign n48829 = ~n48558 & ~n48828;
  assign n48830 = ~n48822 & ~n48829;
  assign n48831 = n48554 & ~n48830;
  assign n48832 = n48549 & ~n48553;
  assign n48833 = n48830 & n48832;
  assign n48834 = ~n48831 & ~n48833;
  assign n48835 = n48553 & ~n48830;
  assign n48836 = n48549 & n48835;
  assign n48837 = ~n48551 & n48830;
  assign n48838 = n48552 & n48837;
  assign n48839 = ~n48549 & n48838;
  assign n48840 = ~n48836 & ~n48839;
  assign n48841 = n48834 & n48840;
  assign n48842 = n48548 & ~n48841;
  assign n48843 = ~n48548 & n48841;
  assign n48844 = ~n48842 & ~n48843;
  assign n48845 = n48547 & ~n48844;
  assign n48846 = ~n48548 & ~n48840;
  assign n48847 = ~n48548 & ~n48834;
  assign n48848 = n48548 & n48834;
  assign n48849 = n48840 & n48848;
  assign n48850 = ~n48846 & ~n48847;
  assign n48851 = ~n48849 & n48850;
  assign n48852 = ~n48547 & ~n48851;
  assign n48853 = ~n48845 & ~n48852;
  assign n48854 = P4_DATAO_REG_5_ & n44372;
  assign n48855 = ~n48215 & n48216;
  assign n48856 = ~n48215 & n48495;
  assign n48857 = ~n48501 & ~n48855;
  assign n48858 = ~n48856 & n48857;
  assign n48859 = ~n48853 & ~n48854;
  assign n48860 = ~n48858 & n48859;
  assign n48861 = n48853 & n48854;
  assign n48862 = ~n48859 & ~n48861;
  assign n48863 = n48858 & n48862;
  assign n48864 = ~n48860 & ~n48863;
  assign n48865 = n48854 & ~n48858;
  assign n48866 = n48853 & n48865;
  assign n48867 = n48864 & ~n48866;
  assign n48868 = n48543 & ~n48867;
  assign n48869 = ~n48543 & n48867;
  assign n48870 = ~n48868 & ~n48869;
  assign n48871 = n48542 & ~n48870;
  assign n48872 = n48543 & ~n48866;
  assign n48873 = n48864 & n48872;
  assign n48874 = ~n48543 & ~n48867;
  assign n48875 = ~n48873 & ~n48874;
  assign n48876 = ~n48542 & ~n48875;
  assign n48877 = ~n48871 & ~n48876;
  assign n48878 = n48538 & n48877;
  assign n48879 = n47274 & ~n48878;
  assign n48880 = ~n48534 & ~n48877;
  assign n48881 = ~n48537 & n48880;
  assign n48882 = n48534 & ~n48877;
  assign n48883 = ~n48534 & n48877;
  assign n48884 = ~n48882 & ~n48883;
  assign n48885 = n48537 & ~n48884;
  assign n48886 = ~n48881 & ~n48885;
  assign n48887 = n48879 & n48886;
  assign n48888 = ~n48532 & ~n48878;
  assign n48889 = n48886 & n48888;
  assign n48890 = ~n48533 & ~n48887;
  assign n48891 = ~n48889 & n48890;
  assign n48892 = n47272 & ~n48891;
  assign n48893 = ~n48537 & ~n48877;
  assign n48894 = ~n48538 & ~n48882;
  assign n48895 = ~n48893 & n48894;
  assign n48896 = P4_DATAO_REG_3_ & n47273;
  assign n48897 = ~n48853 & n48854;
  assign n48898 = ~n48853 & ~n48858;
  assign n48899 = ~n48865 & ~n48897;
  assign n48900 = ~n48898 & n48899;
  assign n48901 = P4_DATAO_REG_5_ & n47277;
  assign n48902 = P4_DATAO_REG_6_ & n44372;
  assign n48903 = ~n48548 & ~n48841;
  assign n48904 = ~n48547 & ~n48903;
  assign n48905 = ~n48849 & ~n48904;
  assign n48906 = ~n48902 & ~n48905;
  assign n48907 = n48549 & ~n48830;
  assign n48908 = ~n48553 & ~n48830;
  assign n48909 = ~n48832 & ~n48907;
  assign n48910 = ~n48908 & n48909;
  assign n48911 = P4_DATAO_REG_7_ & n46777;
  assign n48912 = n48807 & ~n48810;
  assign n48913 = ~n48806 & n48807;
  assign n48914 = ~n48806 & ~n48810;
  assign n48915 = ~n48912 & ~n48913;
  assign n48916 = ~n48914 & n48915;
  assign n48917 = P4_DATAO_REG_9_ & n44376;
  assign n48918 = P4_DATAO_REG_10_ & n44378;
  assign n48919 = ~n48797 & ~n48798;
  assign n48920 = ~n48795 & n48919;
  assign n48921 = ~n48796 & n48920;
  assign n48922 = n48794 & ~n48921;
  assign n48923 = ~n48802 & ~n48922;
  assign n48924 = ~n48918 & ~n48923;
  assign n48925 = P4_DATAO_REG_11_ & n44380;
  assign n48926 = n48565 & ~n48785;
  assign n48927 = ~n48564 & ~n48785;
  assign n48928 = ~n48787 & ~n48926;
  assign n48929 = ~n48927 & n48928;
  assign n48930 = n48925 & ~n48929;
  assign n48931 = ~n48925 & n48929;
  assign n48932 = ~n48766 & n48767;
  assign n48933 = ~n48766 & ~n48769;
  assign n48934 = ~n48776 & ~n48932;
  assign n48935 = ~n48933 & n48934;
  assign n48936 = P4_DATAO_REG_13_ & n45602;
  assign n48937 = ~n48742 & n48743;
  assign n48938 = ~n48742 & ~n48745;
  assign n48939 = ~n48752 & ~n48937;
  assign n48940 = ~n48938 & n48939;
  assign n48941 = P4_DATAO_REG_15_ & n44386;
  assign n48942 = ~n48718 & n48719;
  assign n48943 = ~n48718 & ~n48721;
  assign n48944 = ~n48728 & ~n48942;
  assign n48945 = ~n48943 & n48944;
  assign n48946 = P4_DATAO_REG_17_ & n44390;
  assign n48947 = P4_DATAO_REG_19_ & n44394;
  assign n48948 = ~n48694 & n48695;
  assign n48949 = ~n48694 & ~n48697;
  assign n48950 = ~n48704 & ~n48948;
  assign n48951 = ~n48949 & n48950;
  assign n48952 = n48947 & ~n48951;
  assign n48953 = ~n48947 & n48951;
  assign n48954 = ~n48952 & ~n48953;
  assign n48955 = P4_DATAO_REG_20_ & n44704;
  assign n48956 = ~n48592 & ~n48682;
  assign n48957 = ~n48591 & ~n48956;
  assign n48958 = ~n48689 & ~n48957;
  assign n48959 = ~n48955 & ~n48958;
  assign n48960 = n48593 & ~n48671;
  assign n48961 = n48593 & ~n48596;
  assign n48962 = ~n48596 & ~n48671;
  assign n48963 = ~n48960 & ~n48961;
  assign n48964 = ~n48962 & n48963;
  assign n48965 = P4_DATAO_REG_21_ & n44623;
  assign n48966 = ~n48647 & ~n48651;
  assign n48967 = ~n48648 & ~n48656;
  assign n48968 = ~n48966 & n48967;
  assign n48969 = P4_DATAO_REG_23_ & n44102;
  assign n48970 = n48609 & ~n48628;
  assign n48971 = ~n48611 & ~n48628;
  assign n48972 = ~n48630 & ~n48970;
  assign n48973 = ~n48971 & n48972;
  assign n48974 = P4_DATAO_REG_25_ & n44143;
  assign n48975 = P4_DATAO_REG_27_ & n44108;
  assign n48976 = P4_DATAO_REG_28_ & n44110;
  assign n48977 = P4_DATAO_REG_29_ & n44112;
  assign n48978 = n48976 & ~n48977;
  assign n48979 = ~n48976 & n48977;
  assign n48980 = ~n48978 & ~n48979;
  assign n48981 = n48975 & ~n48980;
  assign n48982 = ~n48975 & n48980;
  assign n48983 = P4_DATAO_REG_27_ & P4_DATAO_REG_28_;
  assign n48984 = n44119 & n48983;
  assign n48985 = ~n48981 & ~n48982;
  assign n48986 = ~n48984 & n48985;
  assign n48987 = n48975 & ~n48978;
  assign n48988 = ~n48975 & n48978;
  assign n48989 = ~n48987 & ~n48988;
  assign n48990 = n48984 & n48989;
  assign n48991 = ~n48986 & ~n48990;
  assign n48992 = P4_DATAO_REG_26_ & n44106;
  assign n48993 = ~n48620 & n48622;
  assign n48994 = ~n48619 & ~n48993;
  assign n48995 = ~n48991 & ~n48992;
  assign n48996 = ~n48994 & n48995;
  assign n48997 = n48991 & n48992;
  assign n48998 = ~n48995 & ~n48997;
  assign n48999 = n48994 & n48998;
  assign n49000 = ~n48996 & ~n48999;
  assign n49001 = n48992 & ~n48994;
  assign n49002 = n48991 & n49001;
  assign n49003 = n49000 & ~n49002;
  assign n49004 = n48974 & ~n49003;
  assign n49005 = ~n48974 & n49003;
  assign n49006 = ~n49004 & ~n49005;
  assign n49007 = n48973 & ~n49006;
  assign n49008 = ~n48974 & n49002;
  assign n49009 = ~n48974 & ~n49000;
  assign n49010 = n48974 & n49000;
  assign n49011 = ~n49002 & n49010;
  assign n49012 = ~n49008 & ~n49009;
  assign n49013 = ~n49011 & n49012;
  assign n49014 = ~n48973 & ~n49013;
  assign n49015 = ~n49007 & ~n49014;
  assign n49016 = P4_DATAO_REG_24_ & n44104;
  assign n49017 = ~n48607 & ~n48644;
  assign n49018 = ~n48643 & ~n49017;
  assign n49019 = ~n49015 & ~n49016;
  assign n49020 = ~n49018 & n49019;
  assign n49021 = n49015 & n49016;
  assign n49022 = ~n49019 & ~n49021;
  assign n49023 = n49018 & n49022;
  assign n49024 = ~n49020 & ~n49023;
  assign n49025 = n49016 & ~n49018;
  assign n49026 = n49015 & n49025;
  assign n49027 = n49024 & ~n49026;
  assign n49028 = n48969 & ~n49027;
  assign n49029 = ~n48969 & n49027;
  assign n49030 = ~n49028 & ~n49029;
  assign n49031 = n48968 & ~n49030;
  assign n49032 = ~n48969 & n49026;
  assign n49033 = n48969 & ~n49026;
  assign n49034 = n49024 & n49033;
  assign n49035 = ~n48969 & ~n49024;
  assign n49036 = ~n49032 & ~n49034;
  assign n49037 = ~n49035 & n49036;
  assign n49038 = ~n48968 & ~n49037;
  assign n49039 = ~n49031 & ~n49038;
  assign n49040 = P4_DATAO_REG_22_ & n44356;
  assign n49041 = ~n48601 & ~n48668;
  assign n49042 = ~n48667 & ~n49041;
  assign n49043 = ~n49039 & ~n49040;
  assign n49044 = ~n49042 & n49043;
  assign n49045 = ~n49039 & n49040;
  assign n49046 = n49039 & ~n49040;
  assign n49047 = ~n49045 & ~n49046;
  assign n49048 = n49042 & ~n49047;
  assign n49049 = ~n49044 & ~n49048;
  assign n49050 = n49040 & ~n49042;
  assign n49051 = n49039 & n49050;
  assign n49052 = n49049 & ~n49051;
  assign n49053 = n48965 & ~n49052;
  assign n49054 = ~n48965 & n49052;
  assign n49055 = ~n49053 & ~n49054;
  assign n49056 = n48964 & ~n49055;
  assign n49057 = n48965 & ~n49051;
  assign n49058 = n49049 & n49057;
  assign n49059 = ~n48965 & ~n49052;
  assign n49060 = ~n49058 & ~n49059;
  assign n49061 = ~n48964 & ~n49060;
  assign n49062 = ~n49056 & ~n49061;
  assign n49063 = n48959 & ~n49062;
  assign n49064 = n48955 & ~n48958;
  assign n49065 = n49062 & n49064;
  assign n49066 = n48958 & ~n49062;
  assign n49067 = n48955 & n49066;
  assign n49068 = n48958 & n49062;
  assign n49069 = ~n48955 & n49068;
  assign n49070 = ~n49063 & ~n49065;
  assign n49071 = ~n49067 & n49070;
  assign n49072 = ~n49069 & n49071;
  assign n49073 = n48954 & ~n49072;
  assign n49074 = ~n48947 & ~n48949;
  assign n49075 = ~n48704 & n49074;
  assign n49076 = ~n48948 & n49075;
  assign n49077 = ~n48952 & ~n49076;
  assign n49078 = n49072 & ~n49077;
  assign n49079 = ~n49073 & ~n49078;
  assign n49080 = P4_DATAO_REG_18_ & n44392;
  assign n49081 = ~n48587 & ~n48706;
  assign n49082 = ~n48586 & ~n49081;
  assign n49083 = ~n48713 & ~n49082;
  assign n49084 = ~n49079 & ~n49080;
  assign n49085 = ~n49083 & n49084;
  assign n49086 = n49079 & n49080;
  assign n49087 = ~n49084 & ~n49086;
  assign n49088 = n49083 & n49087;
  assign n49089 = ~n49085 & ~n49088;
  assign n49090 = n49080 & ~n49083;
  assign n49091 = n49079 & n49090;
  assign n49092 = n49089 & ~n49091;
  assign n49093 = n48946 & ~n49092;
  assign n49094 = ~n48946 & n49092;
  assign n49095 = ~n49093 & ~n49094;
  assign n49096 = n48945 & ~n49095;
  assign n49097 = ~n48946 & n49091;
  assign n49098 = n48946 & ~n49091;
  assign n49099 = n49089 & n49098;
  assign n49100 = ~n48946 & ~n49089;
  assign n49101 = ~n49097 & ~n49099;
  assign n49102 = ~n49100 & n49101;
  assign n49103 = ~n48945 & ~n49102;
  assign n49104 = ~n49096 & ~n49103;
  assign n49105 = P4_DATAO_REG_16_ & n44388;
  assign n49106 = ~n48582 & ~n48730;
  assign n49107 = ~n48581 & ~n49106;
  assign n49108 = ~n48737 & ~n49107;
  assign n49109 = ~n49104 & ~n49105;
  assign n49110 = ~n49108 & n49109;
  assign n49111 = n49104 & n49105;
  assign n49112 = ~n49109 & ~n49111;
  assign n49113 = n49108 & n49112;
  assign n49114 = ~n49110 & ~n49113;
  assign n49115 = n49105 & ~n49108;
  assign n49116 = n49104 & n49115;
  assign n49117 = n49114 & ~n49116;
  assign n49118 = n48941 & ~n49117;
  assign n49119 = ~n48941 & n49117;
  assign n49120 = ~n49118 & ~n49119;
  assign n49121 = n48940 & ~n49120;
  assign n49122 = ~n48941 & n49116;
  assign n49123 = n48941 & ~n49116;
  assign n49124 = n49114 & n49123;
  assign n49125 = ~n48941 & ~n49114;
  assign n49126 = ~n49122 & ~n49124;
  assign n49127 = ~n49125 & n49126;
  assign n49128 = ~n48940 & ~n49127;
  assign n49129 = ~n49121 & ~n49128;
  assign n49130 = P4_DATAO_REG_14_ & n44384;
  assign n49131 = ~n48578 & ~n48754;
  assign n49132 = ~n48577 & ~n49131;
  assign n49133 = ~n48761 & ~n49132;
  assign n49134 = ~n49129 & ~n49130;
  assign n49135 = ~n49133 & n49134;
  assign n49136 = n49129 & n49130;
  assign n49137 = ~n49134 & ~n49136;
  assign n49138 = n49133 & n49137;
  assign n49139 = ~n49135 & ~n49138;
  assign n49140 = n49130 & ~n49133;
  assign n49141 = n49129 & n49140;
  assign n49142 = n49139 & ~n49141;
  assign n49143 = n48936 & ~n49142;
  assign n49144 = ~n48936 & n49142;
  assign n49145 = ~n49143 & ~n49144;
  assign n49146 = n48935 & ~n49145;
  assign n49147 = ~n48936 & n49141;
  assign n49148 = n48936 & ~n49141;
  assign n49149 = n49139 & n49148;
  assign n49150 = ~n48936 & ~n49139;
  assign n49151 = ~n49147 & ~n49149;
  assign n49152 = ~n49150 & n49151;
  assign n49153 = ~n48935 & ~n49152;
  assign n49154 = ~n49146 & ~n49153;
  assign n49155 = ~n48573 & n48778;
  assign n49156 = ~n48572 & ~n49155;
  assign n49157 = P4_DATAO_REG_12_ & n44382;
  assign n49158 = ~n49154 & ~n49156;
  assign n49159 = ~n49157 & n49158;
  assign n49160 = ~n49154 & n49156;
  assign n49161 = n49157 & n49160;
  assign n49162 = ~n49156 & n49157;
  assign n49163 = n49156 & ~n49157;
  assign n49164 = ~n49162 & ~n49163;
  assign n49165 = n49154 & ~n49164;
  assign n49166 = ~n49159 & ~n49161;
  assign n49167 = ~n49165 & n49166;
  assign n49168 = ~n48930 & ~n48931;
  assign n49169 = ~n49167 & n49168;
  assign n49170 = ~n48925 & ~n48927;
  assign n49171 = ~n48926 & n49170;
  assign n49172 = ~n48787 & n49171;
  assign n49173 = ~n48930 & ~n49172;
  assign n49174 = n49167 & ~n49173;
  assign n49175 = ~n49169 & ~n49174;
  assign n49176 = n48924 & ~n49175;
  assign n49177 = n48918 & ~n48923;
  assign n49178 = ~n48918 & n48923;
  assign n49179 = ~n49177 & ~n49178;
  assign n49180 = n49175 & ~n49179;
  assign n49181 = ~n49176 & ~n49180;
  assign n49182 = n48918 & n48923;
  assign n49183 = ~n49175 & n49182;
  assign n49184 = n49181 & ~n49183;
  assign n49185 = n48917 & ~n49184;
  assign n49186 = ~n48917 & n49184;
  assign n49187 = ~n49185 & ~n49186;
  assign n49188 = n48916 & ~n49187;
  assign n49189 = ~n48917 & ~n49175;
  assign n49190 = n49182 & n49189;
  assign n49191 = n48917 & ~n49183;
  assign n49192 = n49181 & n49191;
  assign n49193 = ~n48917 & ~n49181;
  assign n49194 = ~n49190 & ~n49192;
  assign n49195 = ~n49193 & n49194;
  assign n49196 = ~n48916 & ~n49195;
  assign n49197 = ~n49188 & ~n49196;
  assign n49198 = P4_DATAO_REG_8_ & n44374;
  assign n49199 = ~n48559 & ~n48818;
  assign n49200 = ~n48558 & ~n49199;
  assign n49201 = ~n48826 & ~n49200;
  assign n49202 = ~n49197 & ~n49198;
  assign n49203 = ~n49201 & n49202;
  assign n49204 = n49197 & n49198;
  assign n49205 = ~n49202 & ~n49204;
  assign n49206 = n49201 & n49205;
  assign n49207 = ~n49203 & ~n49206;
  assign n49208 = n49198 & ~n49201;
  assign n49209 = n49197 & n49208;
  assign n49210 = n49207 & ~n49209;
  assign n49211 = n48911 & ~n49210;
  assign n49212 = ~n48911 & n49210;
  assign n49213 = ~n49211 & ~n49212;
  assign n49214 = n48910 & ~n49213;
  assign n49215 = ~n48911 & n49209;
  assign n49216 = n48911 & ~n49209;
  assign n49217 = n49207 & n49216;
  assign n49218 = ~n48911 & ~n49207;
  assign n49219 = ~n49215 & ~n49217;
  assign n49220 = ~n49218 & n49219;
  assign n49221 = ~n48910 & ~n49220;
  assign n49222 = ~n49214 & ~n49221;
  assign n49223 = n48906 & ~n49222;
  assign n49224 = n48902 & n48904;
  assign n49225 = ~n48902 & n48905;
  assign n49226 = n48849 & n48902;
  assign n49227 = ~n49224 & ~n49225;
  assign n49228 = ~n49226 & n49227;
  assign n49229 = n49222 & ~n49228;
  assign n49230 = ~n49223 & ~n49229;
  assign n49231 = n48902 & n48905;
  assign n49232 = ~n49222 & n49231;
  assign n49233 = n49230 & ~n49232;
  assign n49234 = n48901 & ~n49233;
  assign n49235 = ~n48901 & n49233;
  assign n49236 = ~n49234 & ~n49235;
  assign n49237 = n48900 & ~n49236;
  assign n49238 = ~n48901 & ~n49222;
  assign n49239 = n49231 & n49238;
  assign n49240 = n48901 & ~n49232;
  assign n49241 = n49230 & n49240;
  assign n49242 = ~n48901 & ~n49230;
  assign n49243 = ~n49239 & ~n49241;
  assign n49244 = ~n49242 & n49243;
  assign n49245 = ~n48900 & ~n49244;
  assign n49246 = ~n49237 & ~n49245;
  assign n49247 = P4_DATAO_REG_4_ & n47275;
  assign n49248 = ~n48542 & ~n48874;
  assign n49249 = ~n48873 & ~n49248;
  assign n49250 = ~n49246 & ~n49247;
  assign n49251 = ~n49249 & n49250;
  assign n49252 = n49246 & n49247;
  assign n49253 = ~n49250 & ~n49252;
  assign n49254 = n49249 & n49253;
  assign n49255 = ~n49251 & ~n49254;
  assign n49256 = n49247 & ~n49249;
  assign n49257 = n49246 & n49256;
  assign n49258 = n49255 & ~n49257;
  assign n49259 = n48896 & ~n49258;
  assign n49260 = ~n48896 & n49258;
  assign n49261 = ~n49259 & ~n49260;
  assign n49262 = n48895 & ~n49261;
  assign n49263 = ~n48896 & n49257;
  assign n49264 = n48896 & ~n49257;
  assign n49265 = n49255 & n49264;
  assign n49266 = ~n48896 & ~n49255;
  assign n49267 = ~n49263 & ~n49265;
  assign n49268 = ~n49266 & n49267;
  assign n49269 = ~n48895 & ~n49268;
  assign n49270 = ~n49262 & ~n49269;
  assign n49271 = n48892 & n49270;
  assign n49272 = n47270 & ~n49271;
  assign n49273 = ~n47272 & ~n49270;
  assign n49274 = ~n48891 & n49273;
  assign n49275 = n47272 & n49270;
  assign n49276 = ~n49273 & ~n49275;
  assign n49277 = n48891 & n49276;
  assign n49278 = ~n49274 & ~n49277;
  assign n49279 = n49272 & n49278;
  assign n49280 = ~n49271 & n49278;
  assign n49281 = ~n47270 & ~n49280;
  assign n49282 = P4_DATAO_REG_1_ & n47271;
  assign n49283 = P4_DATAO_REG_1_ & n47275;
  assign n49284 = P4_DATAO_REG_1_ & n47277;
  assign n49285 = ~n48176 & ~n48177;
  assign n49286 = ~n48180 & ~n49285;
  assign n49287 = n48180 & n49285;
  assign n49288 = ~n49286 & ~n49287;
  assign n49289 = ~n44372 & ~n46777;
  assign n49290 = ~n47070 & n49289;
  assign n49291 = P4_DATAO_REG_1_ & n44372;
  assign n49292 = ~n47075 & ~n49291;
  assign n49293 = n46776 & n49292;
  assign n49294 = ~n49288 & ~n49290;
  assign n49295 = ~n49293 & n49294;
  assign n49296 = ~n46778 & ~n47070;
  assign n49297 = ~n46776 & ~n49296;
  assign n49298 = ~n47075 & ~n49297;
  assign n49299 = n49291 & ~n49298;
  assign n49300 = ~n49295 & ~n49299;
  assign n49301 = n49284 & ~n49300;
  assign n49302 = ~n48169 & n48182;
  assign n49303 = ~n48183 & ~n49302;
  assign n49304 = n48193 & ~n49303;
  assign n49305 = ~n48193 & n49303;
  assign n49306 = ~n49304 & ~n49305;
  assign n49307 = ~n49284 & n49300;
  assign n49308 = n49306 & ~n49307;
  assign n49309 = ~n49301 & ~n49308;
  assign n49310 = n49283 & ~n49309;
  assign n49311 = ~n48167 & ~n48168;
  assign n49312 = n48197 & n49311;
  assign n49313 = ~n48197 & ~n49311;
  assign n49314 = ~n49312 & ~n49313;
  assign n49315 = n49283 & ~n49314;
  assign n49316 = ~n49309 & ~n49314;
  assign n49317 = ~n49310 & ~n49315;
  assign n49318 = ~n49316 & n49317;
  assign n49319 = n47276 & ~n48167;
  assign n49320 = ~n48198 & n49319;
  assign n49321 = ~n48528 & n49320;
  assign n49322 = n48200 & n48528;
  assign n49323 = ~n49321 & ~n49322;
  assign n49324 = ~n47276 & ~n48199;
  assign n49325 = ~n48528 & n49324;
  assign n49326 = ~n47276 & ~n48167;
  assign n49327 = ~n48198 & n49326;
  assign n49328 = n48528 & n49327;
  assign n49329 = ~n49325 & ~n49328;
  assign n49330 = n49323 & n49329;
  assign n49331 = P4_DATAO_REG_1_ & n47273;
  assign n49332 = n49330 & n49331;
  assign n49333 = ~n49282 & n49318;
  assign n49334 = ~n49332 & n49333;
  assign n49335 = ~n47271 & ~n47273;
  assign n49336 = ~n49330 & n49335;
  assign n49337 = ~n49334 & ~n49336;
  assign n49338 = ~n48878 & n48886;
  assign n49339 = n47274 & ~n49338;
  assign n49340 = ~n47274 & n49338;
  assign n49341 = ~n49339 & ~n49340;
  assign n49342 = n48532 & ~n49341;
  assign n49343 = ~n47274 & ~n49338;
  assign n49344 = ~n48887 & ~n49343;
  assign n49345 = ~n48532 & ~n49344;
  assign n49346 = ~n49342 & ~n49345;
  assign n49347 = n49337 & ~n49346;
  assign n49348 = ~n49323 & ~n49331;
  assign n49349 = ~n49329 & ~n49331;
  assign n49350 = ~n49318 & ~n49348;
  assign n49351 = ~n49349 & n49350;
  assign n49352 = ~n49332 & ~n49351;
  assign n49353 = n49282 & ~n49352;
  assign n49354 = ~n49347 & ~n49353;
  assign n49355 = ~n49281 & ~n49354;
  assign n49356 = ~n49279 & ~n49355;
  assign n49357 = n47268 & ~n49356;
  assign n49358 = n47272 & ~n49270;
  assign n49359 = ~n48891 & ~n49270;
  assign n49360 = ~n48892 & ~n49358;
  assign n49361 = ~n49359 & n49360;
  assign n49362 = P4_DATAO_REG_2_ & n47269;
  assign n49363 = ~n49246 & n49247;
  assign n49364 = ~n49246 & ~n49249;
  assign n49365 = ~n49256 & ~n49363;
  assign n49366 = ~n49364 & n49365;
  assign n49367 = P4_DATAO_REG_4_ & n47273;
  assign n49368 = P4_DATAO_REG_5_ & n47275;
  assign n49369 = ~n49239 & ~n49242;
  assign n49370 = ~n48900 & n49369;
  assign n49371 = ~n49241 & ~n49370;
  assign n49372 = ~n49368 & ~n49371;
  assign n49373 = P4_DATAO_REG_6_ & n47277;
  assign n49374 = n48902 & ~n49222;
  assign n49375 = n48902 & ~n48905;
  assign n49376 = ~n48905 & ~n49222;
  assign n49377 = ~n49374 & ~n49375;
  assign n49378 = ~n49376 & n49377;
  assign n49379 = n49373 & ~n49378;
  assign n49380 = ~n49373 & n49378;
  assign n49381 = ~n49379 & ~n49380;
  assign n49382 = P4_DATAO_REG_7_ & n44372;
  assign n49383 = ~n48911 & ~n49210;
  assign n49384 = ~n48910 & ~n49383;
  assign n49385 = ~n49217 & ~n49384;
  assign n49386 = ~n49382 & ~n49385;
  assign n49387 = P4_DATAO_REG_8_ & n46777;
  assign n49388 = ~n49197 & n49198;
  assign n49389 = ~n49197 & ~n49201;
  assign n49390 = ~n49208 & ~n49388;
  assign n49391 = ~n49389 & n49390;
  assign n49392 = n49387 & ~n49391;
  assign n49393 = ~n49387 & n49391;
  assign n49394 = ~n49392 & ~n49393;
  assign n49395 = ~n48917 & ~n49184;
  assign n49396 = ~n48916 & ~n49395;
  assign n49397 = ~n49192 & ~n49396;
  assign n49398 = P4_DATAO_REG_9_ & n44374;
  assign n49399 = n49397 & n49398;
  assign n49400 = n48918 & ~n49175;
  assign n49401 = ~n48923 & ~n49175;
  assign n49402 = ~n49177 & ~n49400;
  assign n49403 = ~n49401 & n49402;
  assign n49404 = P4_DATAO_REG_10_ & n44376;
  assign n49405 = ~n49154 & n49157;
  assign n49406 = ~n49162 & ~n49405;
  assign n49407 = ~n49158 & n49406;
  assign n49408 = P4_DATAO_REG_12_ & n44380;
  assign n49409 = ~n49129 & n49130;
  assign n49410 = ~n49129 & ~n49133;
  assign n49411 = ~n49140 & ~n49409;
  assign n49412 = ~n49410 & n49411;
  assign n49413 = P4_DATAO_REG_14_ & n45602;
  assign n49414 = ~n49104 & n49105;
  assign n49415 = ~n49104 & ~n49108;
  assign n49416 = ~n49115 & ~n49414;
  assign n49417 = ~n49415 & n49416;
  assign n49418 = P4_DATAO_REG_16_ & n44386;
  assign n49419 = ~n49079 & n49080;
  assign n49420 = ~n49079 & ~n49083;
  assign n49421 = ~n49090 & ~n49419;
  assign n49422 = ~n49420 & n49421;
  assign n49423 = P4_DATAO_REG_18_ & n44390;
  assign n49424 = n48955 & ~n49062;
  assign n49425 = ~n48958 & ~n49062;
  assign n49426 = ~n49064 & ~n49424;
  assign n49427 = ~n49425 & n49426;
  assign n49428 = P4_DATAO_REG_20_ & n44394;
  assign n49429 = ~n49039 & ~n49042;
  assign n49430 = ~n49045 & ~n49050;
  assign n49431 = ~n49429 & n49430;
  assign n49432 = P4_DATAO_REG_22_ & n44623;
  assign n49433 = ~n49015 & n49016;
  assign n49434 = ~n49015 & ~n49018;
  assign n49435 = ~n49025 & ~n49433;
  assign n49436 = ~n49434 & n49435;
  assign n49437 = P4_DATAO_REG_24_ & n44102;
  assign n49438 = ~n48991 & n48992;
  assign n49439 = ~n48991 & ~n48994;
  assign n49440 = ~n49001 & ~n49438;
  assign n49441 = ~n49439 & n49440;
  assign n49442 = P4_DATAO_REG_26_ & n44143;
  assign n49443 = P4_DATAO_REG_28_ & n44108;
  assign n49444 = P4_DATAO_REG_29_ & n44110;
  assign n49445 = P4_DATAO_REG_30_ & n44112;
  assign n49446 = n49444 & ~n49445;
  assign n49447 = ~n49444 & n49445;
  assign n49448 = ~n49446 & ~n49447;
  assign n49449 = n49443 & ~n49448;
  assign n49450 = ~n49443 & n49448;
  assign n49451 = P4_DATAO_REG_28_ & P4_DATAO_REG_29_;
  assign n49452 = n44119 & n49451;
  assign n49453 = ~n49449 & ~n49450;
  assign n49454 = ~n49452 & n49453;
  assign n49455 = ~n49443 & ~n49446;
  assign n49456 = n49443 & ~n49445;
  assign n49457 = ~n49455 & ~n49456;
  assign n49458 = n49452 & ~n49457;
  assign n49459 = ~n49454 & ~n49458;
  assign n49460 = P4_DATAO_REG_27_ & n44106;
  assign n49461 = ~n48982 & n48984;
  assign n49462 = ~n48981 & ~n49461;
  assign n49463 = ~n49459 & ~n49460;
  assign n49464 = ~n49462 & n49463;
  assign n49465 = n49459 & n49460;
  assign n49466 = ~n49463 & ~n49465;
  assign n49467 = n49462 & n49466;
  assign n49468 = ~n49464 & ~n49467;
  assign n49469 = n49460 & ~n49462;
  assign n49470 = n49459 & n49469;
  assign n49471 = n49468 & ~n49470;
  assign n49472 = n49442 & ~n49471;
  assign n49473 = ~n49442 & n49471;
  assign n49474 = ~n49472 & ~n49473;
  assign n49475 = n49441 & ~n49474;
  assign n49476 = ~n49442 & n49470;
  assign n49477 = ~n49442 & ~n49468;
  assign n49478 = n49442 & n49468;
  assign n49479 = ~n49470 & n49478;
  assign n49480 = ~n49476 & ~n49477;
  assign n49481 = ~n49479 & n49480;
  assign n49482 = ~n49441 & ~n49481;
  assign n49483 = ~n49475 & ~n49482;
  assign n49484 = P4_DATAO_REG_25_ & n44104;
  assign n49485 = ~n48974 & ~n49003;
  assign n49486 = ~n48973 & ~n49485;
  assign n49487 = ~n49011 & ~n49486;
  assign n49488 = ~n49483 & ~n49484;
  assign n49489 = ~n49487 & n49488;
  assign n49490 = n49483 & n49484;
  assign n49491 = ~n49488 & ~n49490;
  assign n49492 = n49487 & n49491;
  assign n49493 = ~n49489 & ~n49492;
  assign n49494 = n49484 & ~n49487;
  assign n49495 = n49483 & n49494;
  assign n49496 = n49493 & ~n49495;
  assign n49497 = n49437 & ~n49496;
  assign n49498 = ~n49437 & n49496;
  assign n49499 = ~n49497 & ~n49498;
  assign n49500 = n49436 & ~n49499;
  assign n49501 = ~n49437 & n49495;
  assign n49502 = n49437 & ~n49495;
  assign n49503 = n49493 & n49502;
  assign n49504 = ~n49437 & ~n49493;
  assign n49505 = ~n49501 & ~n49503;
  assign n49506 = ~n49504 & n49505;
  assign n49507 = ~n49436 & ~n49506;
  assign n49508 = ~n49500 & ~n49507;
  assign n49509 = P4_DATAO_REG_23_ & n44356;
  assign n49510 = ~n48969 & ~n49027;
  assign n49511 = ~n48968 & ~n49510;
  assign n49512 = ~n49034 & ~n49511;
  assign n49513 = ~n49508 & ~n49509;
  assign n49514 = ~n49512 & n49513;
  assign n49515 = n49508 & n49509;
  assign n49516 = ~n49513 & ~n49515;
  assign n49517 = n49512 & n49516;
  assign n49518 = ~n49514 & ~n49517;
  assign n49519 = n49509 & ~n49512;
  assign n49520 = n49508 & n49519;
  assign n49521 = n49518 & ~n49520;
  assign n49522 = n49432 & ~n49521;
  assign n49523 = ~n49432 & n49521;
  assign n49524 = ~n49522 & ~n49523;
  assign n49525 = n49431 & ~n49524;
  assign n49526 = ~n49432 & n49520;
  assign n49527 = n49432 & ~n49520;
  assign n49528 = n49518 & n49527;
  assign n49529 = ~n49432 & ~n49518;
  assign n49530 = ~n49526 & ~n49528;
  assign n49531 = ~n49529 & n49530;
  assign n49532 = ~n49431 & ~n49531;
  assign n49533 = ~n49525 & ~n49532;
  assign n49534 = P4_DATAO_REG_21_ & n44704;
  assign n49535 = ~n48964 & ~n49059;
  assign n49536 = ~n49058 & ~n49535;
  assign n49537 = ~n49533 & ~n49534;
  assign n49538 = ~n49536 & n49537;
  assign n49539 = n49533 & n49534;
  assign n49540 = ~n49537 & ~n49539;
  assign n49541 = n49536 & n49540;
  assign n49542 = ~n49538 & ~n49541;
  assign n49543 = n49534 & ~n49536;
  assign n49544 = n49533 & n49543;
  assign n49545 = n49542 & ~n49544;
  assign n49546 = n49428 & ~n49545;
  assign n49547 = ~n49428 & n49545;
  assign n49548 = ~n49546 & ~n49547;
  assign n49549 = n49427 & ~n49548;
  assign n49550 = ~n49428 & n49544;
  assign n49551 = ~n49428 & ~n49542;
  assign n49552 = n49428 & ~n49544;
  assign n49553 = n49542 & n49552;
  assign n49554 = ~n49550 & ~n49551;
  assign n49555 = ~n49553 & n49554;
  assign n49556 = ~n49427 & ~n49555;
  assign n49557 = ~n49549 & ~n49556;
  assign n49558 = P4_DATAO_REG_19_ & n44392;
  assign n49559 = ~n48953 & n49072;
  assign n49560 = ~n48952 & ~n49559;
  assign n49561 = ~n49557 & ~n49558;
  assign n49562 = ~n49560 & n49561;
  assign n49563 = n49557 & n49558;
  assign n49564 = ~n49561 & ~n49563;
  assign n49565 = n49560 & n49564;
  assign n49566 = ~n49562 & ~n49565;
  assign n49567 = n49558 & ~n49560;
  assign n49568 = n49557 & n49567;
  assign n49569 = n49566 & ~n49568;
  assign n49570 = n49423 & ~n49569;
  assign n49571 = ~n49423 & n49569;
  assign n49572 = ~n49570 & ~n49571;
  assign n49573 = n49422 & ~n49572;
  assign n49574 = ~n49423 & n49568;
  assign n49575 = ~n49423 & ~n49566;
  assign n49576 = n49423 & ~n49568;
  assign n49577 = n49566 & n49576;
  assign n49578 = ~n49574 & ~n49575;
  assign n49579 = ~n49577 & n49578;
  assign n49580 = ~n49422 & ~n49579;
  assign n49581 = ~n49573 & ~n49580;
  assign n49582 = P4_DATAO_REG_17_ & n44388;
  assign n49583 = ~n48946 & ~n49092;
  assign n49584 = ~n48945 & ~n49583;
  assign n49585 = ~n49099 & ~n49584;
  assign n49586 = ~n49581 & ~n49582;
  assign n49587 = ~n49585 & n49586;
  assign n49588 = n49581 & n49582;
  assign n49589 = ~n49586 & ~n49588;
  assign n49590 = n49585 & n49589;
  assign n49591 = ~n49587 & ~n49590;
  assign n49592 = n49582 & ~n49585;
  assign n49593 = n49581 & n49592;
  assign n49594 = n49591 & ~n49593;
  assign n49595 = n49418 & ~n49594;
  assign n49596 = ~n49418 & n49594;
  assign n49597 = ~n49595 & ~n49596;
  assign n49598 = n49417 & ~n49597;
  assign n49599 = ~n49418 & n49593;
  assign n49600 = n49418 & ~n49593;
  assign n49601 = n49591 & n49600;
  assign n49602 = ~n49418 & ~n49591;
  assign n49603 = ~n49599 & ~n49601;
  assign n49604 = ~n49602 & n49603;
  assign n49605 = ~n49417 & ~n49604;
  assign n49606 = ~n49598 & ~n49605;
  assign n49607 = P4_DATAO_REG_15_ & n44384;
  assign n49608 = ~n48941 & ~n49117;
  assign n49609 = ~n48940 & ~n49608;
  assign n49610 = ~n49124 & ~n49609;
  assign n49611 = ~n49606 & ~n49607;
  assign n49612 = ~n49610 & n49611;
  assign n49613 = n49606 & n49607;
  assign n49614 = ~n49611 & ~n49613;
  assign n49615 = n49610 & n49614;
  assign n49616 = ~n49612 & ~n49615;
  assign n49617 = n49607 & ~n49610;
  assign n49618 = n49606 & n49617;
  assign n49619 = n49616 & ~n49618;
  assign n49620 = n49413 & ~n49619;
  assign n49621 = ~n49413 & n49619;
  assign n49622 = ~n49620 & ~n49621;
  assign n49623 = n49412 & ~n49622;
  assign n49624 = ~n49413 & n49618;
  assign n49625 = n49413 & ~n49618;
  assign n49626 = n49616 & n49625;
  assign n49627 = ~n49413 & ~n49616;
  assign n49628 = ~n49624 & ~n49626;
  assign n49629 = ~n49627 & n49628;
  assign n49630 = ~n49412 & ~n49629;
  assign n49631 = ~n49623 & ~n49630;
  assign n49632 = P4_DATAO_REG_13_ & n44382;
  assign n49633 = ~n48936 & ~n49142;
  assign n49634 = ~n48935 & ~n49633;
  assign n49635 = ~n49149 & ~n49634;
  assign n49636 = ~n49631 & ~n49632;
  assign n49637 = ~n49635 & n49636;
  assign n49638 = n49631 & n49632;
  assign n49639 = ~n49636 & ~n49638;
  assign n49640 = n49635 & n49639;
  assign n49641 = ~n49637 & ~n49640;
  assign n49642 = n49632 & ~n49635;
  assign n49643 = n49631 & n49642;
  assign n49644 = n49641 & ~n49643;
  assign n49645 = n49408 & ~n49644;
  assign n49646 = ~n49408 & n49644;
  assign n49647 = ~n49645 & ~n49646;
  assign n49648 = n49407 & ~n49647;
  assign n49649 = ~n49408 & n49643;
  assign n49650 = n49408 & ~n49643;
  assign n49651 = n49641 & n49650;
  assign n49652 = ~n49408 & ~n49641;
  assign n49653 = ~n49649 & ~n49651;
  assign n49654 = ~n49652 & n49653;
  assign n49655 = ~n49407 & ~n49654;
  assign n49656 = ~n49648 & ~n49655;
  assign n49657 = P4_DATAO_REG_11_ & n44378;
  assign n49658 = ~n48931 & n49167;
  assign n49659 = ~n48930 & ~n49658;
  assign n49660 = ~n49656 & ~n49657;
  assign n49661 = ~n49659 & n49660;
  assign n49662 = n49656 & n49657;
  assign n49663 = ~n49660 & ~n49662;
  assign n49664 = n49659 & n49663;
  assign n49665 = ~n49661 & ~n49664;
  assign n49666 = n49657 & ~n49659;
  assign n49667 = n49656 & n49666;
  assign n49668 = n49665 & ~n49667;
  assign n49669 = n49404 & ~n49668;
  assign n49670 = ~n49404 & n49668;
  assign n49671 = ~n49669 & ~n49670;
  assign n49672 = n49403 & ~n49671;
  assign n49673 = ~n49404 & n49667;
  assign n49674 = n49404 & ~n49667;
  assign n49675 = n49665 & n49674;
  assign n49676 = ~n49404 & ~n49665;
  assign n49677 = ~n49673 & ~n49675;
  assign n49678 = ~n49676 & n49677;
  assign n49679 = ~n49403 & ~n49678;
  assign n49680 = ~n49672 & ~n49679;
  assign n49681 = n49399 & ~n49680;
  assign n49682 = ~n49397 & n49398;
  assign n49683 = n49397 & ~n49398;
  assign n49684 = ~n49682 & ~n49683;
  assign n49685 = n49680 & ~n49684;
  assign n49686 = ~n49681 & ~n49685;
  assign n49687 = ~n49397 & ~n49398;
  assign n49688 = ~n49680 & n49687;
  assign n49689 = n49686 & ~n49688;
  assign n49690 = n49394 & ~n49689;
  assign n49691 = ~n49394 & n49689;
  assign n49692 = ~n49690 & ~n49691;
  assign n49693 = n49386 & ~n49692;
  assign n49694 = n49382 & ~n49385;
  assign n49695 = n49692 & n49694;
  assign n49696 = n49385 & ~n49692;
  assign n49697 = n49382 & n49696;
  assign n49698 = n49385 & n49692;
  assign n49699 = ~n49382 & n49698;
  assign n49700 = ~n49693 & ~n49695;
  assign n49701 = ~n49697 & n49700;
  assign n49702 = ~n49699 & n49701;
  assign n49703 = n49381 & ~n49702;
  assign n49704 = ~n49381 & n49702;
  assign n49705 = ~n49703 & ~n49704;
  assign n49706 = n49372 & ~n49705;
  assign n49707 = n49368 & ~n49371;
  assign n49708 = ~n49241 & ~n49368;
  assign n49709 = ~n49370 & n49708;
  assign n49710 = ~n49707 & ~n49709;
  assign n49711 = n49705 & ~n49710;
  assign n49712 = ~n49706 & ~n49711;
  assign n49713 = n49368 & n49371;
  assign n49714 = ~n49705 & n49713;
  assign n49715 = n49712 & ~n49714;
  assign n49716 = n49367 & ~n49715;
  assign n49717 = ~n49367 & n49715;
  assign n49718 = ~n49716 & ~n49717;
  assign n49719 = n49366 & ~n49718;
  assign n49720 = ~n49367 & ~n49705;
  assign n49721 = n49713 & n49720;
  assign n49722 = ~n49367 & ~n49712;
  assign n49723 = n49367 & ~n49714;
  assign n49724 = n49712 & n49723;
  assign n49725 = ~n49721 & ~n49722;
  assign n49726 = ~n49724 & n49725;
  assign n49727 = ~n49366 & ~n49726;
  assign n49728 = ~n49719 & ~n49727;
  assign n49729 = P4_DATAO_REG_3_ & n47271;
  assign n49730 = ~n48896 & ~n49258;
  assign n49731 = ~n48895 & ~n49730;
  assign n49732 = ~n49265 & ~n49731;
  assign n49733 = ~n49728 & ~n49729;
  assign n49734 = ~n49732 & n49733;
  assign n49735 = n49728 & n49729;
  assign n49736 = ~n49733 & ~n49735;
  assign n49737 = n49732 & n49736;
  assign n49738 = ~n49734 & ~n49737;
  assign n49739 = n49729 & ~n49732;
  assign n49740 = n49728 & n49739;
  assign n49741 = n49738 & ~n49740;
  assign n49742 = n49362 & ~n49741;
  assign n49743 = ~n49362 & n49741;
  assign n49744 = ~n49742 & ~n49743;
  assign n49745 = n49361 & ~n49744;
  assign n49746 = ~n49362 & n49740;
  assign n49747 = n49362 & ~n49740;
  assign n49748 = n49738 & n49747;
  assign n49749 = ~n49362 & ~n49738;
  assign n49750 = ~n49746 & ~n49748;
  assign n49751 = ~n49749 & n49750;
  assign n49752 = ~n49361 & ~n49751;
  assign n49753 = ~n49745 & ~n49752;
  assign n49754 = n47268 & ~n49753;
  assign n49755 = ~n49356 & ~n49753;
  assign n49756 = ~n49357 & ~n49754;
  assign n49757 = ~n49755 & n49756;
  assign n49758 = ~n49362 & ~n49741;
  assign n49759 = ~n49361 & ~n49758;
  assign n49760 = ~n49748 & ~n49759;
  assign n49761 = SEL & DIN_30_;
  assign n49762 = P4_DATAO_REG_1_ & n49761;
  assign n49763 = P4_DATAO_REG_2_ & n47267;
  assign n49764 = n49762 & ~n49763;
  assign n49765 = ~n49762 & n49763;
  assign n49766 = ~n49764 & ~n49765;
  assign n49767 = ~n49728 & n49729;
  assign n49768 = ~n49728 & ~n49732;
  assign n49769 = ~n49739 & ~n49767;
  assign n49770 = ~n49768 & n49769;
  assign n49771 = n49368 & ~n49705;
  assign n49772 = ~n49371 & ~n49705;
  assign n49773 = ~n49707 & ~n49771;
  assign n49774 = ~n49772 & n49773;
  assign n49775 = P4_DATAO_REG_4_ & n47271;
  assign n49776 = ~n49380 & n49702;
  assign n49777 = ~n49379 & ~n49776;
  assign n49778 = n49382 & ~n49692;
  assign n49779 = ~n49385 & ~n49692;
  assign n49780 = ~n49694 & ~n49778;
  assign n49781 = ~n49779 & n49780;
  assign n49782 = ~n49393 & n49689;
  assign n49783 = ~n49392 & ~n49782;
  assign n49784 = ~n49404 & ~n49668;
  assign n49785 = ~n49403 & ~n49784;
  assign n49786 = ~n49675 & ~n49785;
  assign n49787 = P4_DATAO_REG_11_ & n44376;
  assign n49788 = ~n49656 & n49657;
  assign n49789 = ~n49656 & ~n49659;
  assign n49790 = ~n49666 & ~n49788;
  assign n49791 = ~n49789 & n49790;
  assign n49792 = ~n49408 & ~n49644;
  assign n49793 = ~n49407 & ~n49792;
  assign n49794 = ~n49651 & ~n49793;
  assign n49795 = ~n49631 & n49632;
  assign n49796 = ~n49631 & ~n49635;
  assign n49797 = ~n49642 & ~n49795;
  assign n49798 = ~n49796 & n49797;
  assign n49799 = ~n49413 & ~n49619;
  assign n49800 = ~n49412 & ~n49799;
  assign n49801 = ~n49626 & ~n49800;
  assign n49802 = ~n49606 & n49607;
  assign n49803 = ~n49606 & ~n49610;
  assign n49804 = ~n49617 & ~n49802;
  assign n49805 = ~n49803 & n49804;
  assign n49806 = ~n49418 & ~n49594;
  assign n49807 = ~n49417 & ~n49806;
  assign n49808 = ~n49601 & ~n49807;
  assign n49809 = P4_DATAO_REG_15_ & n45602;
  assign n49810 = P4_DATAO_REG_16_ & n44384;
  assign n49811 = n49809 & ~n49810;
  assign n49812 = ~n49809 & n49810;
  assign n49813 = ~n49811 & ~n49812;
  assign n49814 = ~n49581 & n49582;
  assign n49815 = ~n49581 & ~n49585;
  assign n49816 = ~n49592 & ~n49814;
  assign n49817 = ~n49815 & n49816;
  assign n49818 = ~n49557 & n49558;
  assign n49819 = ~n49557 & ~n49560;
  assign n49820 = ~n49567 & ~n49818;
  assign n49821 = ~n49819 & n49820;
  assign n49822 = ~n49428 & ~n49545;
  assign n49823 = ~n49427 & ~n49822;
  assign n49824 = ~n49553 & ~n49823;
  assign n49825 = ~n49432 & ~n49521;
  assign n49826 = ~n49431 & ~n49825;
  assign n49827 = ~n49528 & ~n49826;
  assign n49828 = ~n49508 & n49509;
  assign n49829 = ~n49508 & ~n49512;
  assign n49830 = ~n49519 & ~n49828;
  assign n49831 = ~n49829 & n49830;
  assign n49832 = P4_DATAO_REG_22_ & n44704;
  assign n49833 = P4_DATAO_REG_23_ & n44623;
  assign n49834 = n49832 & ~n49833;
  assign n49835 = ~n49832 & n49833;
  assign n49836 = ~n49834 & ~n49835;
  assign n49837 = P4_DATAO_REG_25_ & n44102;
  assign n49838 = P4_DATAO_REG_24_ & n44356;
  assign n49839 = n49837 & ~n49838;
  assign n49840 = ~n49837 & n49838;
  assign n49841 = ~n49839 & ~n49840;
  assign n49842 = P4_DATAO_REG_29_ & n44119;
  assign n49843 = n44108 & n49842;
  assign n49844 = P4_DATAO_REG_29_ & n44108;
  assign n49845 = P4_DATAO_REG_30_ & n44110;
  assign n49846 = ~n44112 & ~n49845;
  assign n49847 = P4_DATAO_REG_31_ & n49846;
  assign n49848 = ~P4_DATAO_REG_31_ & n49845;
  assign n49849 = P4_DATAO_REG_30_ & n44119;
  assign n49850 = ~n49847 & ~n49848;
  assign n49851 = ~n49849 & n49850;
  assign n49852 = n49844 & ~n49851;
  assign n49853 = ~n49844 & n49851;
  assign n49854 = ~n49852 & ~n49853;
  assign n49855 = ~n49842 & n49854;
  assign n49856 = ~n49843 & ~n49855;
  assign n49857 = ~n49450 & n49452;
  assign n49858 = ~n49449 & ~n49857;
  assign n49859 = P4_DATAO_REG_28_ & n44106;
  assign n49860 = n49858 & ~n49859;
  assign n49861 = ~n49858 & n49859;
  assign n49862 = ~n49860 & ~n49861;
  assign n49863 = ~n49856 & n49862;
  assign n49864 = n49856 & ~n49862;
  assign n49865 = ~n49863 & ~n49864;
  assign n49866 = ~n49459 & n49460;
  assign n49867 = ~n49459 & ~n49462;
  assign n49868 = ~n49469 & ~n49866;
  assign n49869 = ~n49867 & n49868;
  assign n49870 = P4_DATAO_REG_26_ & n44104;
  assign n49871 = P4_DATAO_REG_27_ & n44143;
  assign n49872 = n49870 & ~n49871;
  assign n49873 = ~n49870 & n49871;
  assign n49874 = ~n49872 & ~n49873;
  assign n49875 = n49869 & n49874;
  assign n49876 = ~n49869 & ~n49874;
  assign n49877 = ~n49875 & ~n49876;
  assign n49878 = ~n49865 & n49877;
  assign n49879 = n49865 & ~n49877;
  assign n49880 = ~n49878 & ~n49879;
  assign n49881 = ~n49442 & ~n49471;
  assign n49882 = ~n49441 & ~n49881;
  assign n49883 = ~n49479 & ~n49882;
  assign n49884 = ~n49880 & ~n49883;
  assign n49885 = n49880 & n49883;
  assign n49886 = ~n49884 & ~n49885;
  assign n49887 = ~n49841 & n49886;
  assign n49888 = n49841 & ~n49886;
  assign n49889 = ~n49887 & ~n49888;
  assign n49890 = ~n49483 & n49484;
  assign n49891 = ~n49483 & ~n49487;
  assign n49892 = ~n49494 & ~n49890;
  assign n49893 = ~n49891 & n49892;
  assign n49894 = ~n49889 & ~n49893;
  assign n49895 = n49889 & n49893;
  assign n49896 = ~n49894 & ~n49895;
  assign n49897 = ~n49437 & ~n49496;
  assign n49898 = ~n49436 & ~n49897;
  assign n49899 = ~n49503 & ~n49898;
  assign n49900 = ~n49896 & ~n49899;
  assign n49901 = n49896 & n49899;
  assign n49902 = ~n49900 & ~n49901;
  assign n49903 = ~n49836 & n49902;
  assign n49904 = n49836 & ~n49902;
  assign n49905 = ~n49903 & ~n49904;
  assign n49906 = n49831 & n49905;
  assign n49907 = ~n49831 & ~n49905;
  assign n49908 = ~n49906 & ~n49907;
  assign n49909 = n49827 & n49908;
  assign n49910 = ~n49827 & ~n49908;
  assign n49911 = ~n49909 & ~n49910;
  assign n49912 = ~n49533 & n49534;
  assign n49913 = ~n49533 & ~n49536;
  assign n49914 = ~n49543 & ~n49912;
  assign n49915 = ~n49913 & n49914;
  assign n49916 = ~n49911 & ~n49915;
  assign n49917 = n49911 & n49915;
  assign n49918 = ~n49916 & ~n49917;
  assign n49919 = n49824 & n49918;
  assign n49920 = ~n49824 & ~n49918;
  assign n49921 = ~n49919 & ~n49920;
  assign n49922 = P4_DATAO_REG_19_ & n44390;
  assign n49923 = P4_DATAO_REG_21_ & n44394;
  assign n49924 = P4_DATAO_REG_20_ & n44392;
  assign n49925 = n49923 & ~n49924;
  assign n49926 = ~n49923 & n49924;
  assign n49927 = ~n49925 & ~n49926;
  assign n49928 = n49922 & n49927;
  assign n49929 = ~n49922 & ~n49927;
  assign n49930 = ~n49928 & ~n49929;
  assign n49931 = ~n49921 & n49930;
  assign n49932 = n49921 & ~n49930;
  assign n49933 = ~n49931 & ~n49932;
  assign n49934 = P4_DATAO_REG_18_ & n44388;
  assign n49935 = ~n49933 & ~n49934;
  assign n49936 = n49933 & n49934;
  assign n49937 = ~n49935 & ~n49936;
  assign n49938 = n49821 & n49937;
  assign n49939 = ~n49821 & ~n49937;
  assign n49940 = ~n49938 & ~n49939;
  assign n49941 = P4_DATAO_REG_17_ & n44386;
  assign n49942 = ~n49940 & ~n49941;
  assign n49943 = n49940 & n49941;
  assign n49944 = ~n49942 & ~n49943;
  assign n49945 = ~n49423 & ~n49569;
  assign n49946 = ~n49422 & ~n49945;
  assign n49947 = ~n49577 & ~n49946;
  assign n49948 = ~n49944 & ~n49947;
  assign n49949 = n49944 & n49947;
  assign n49950 = ~n49948 & ~n49949;
  assign n49951 = n49817 & n49950;
  assign n49952 = ~n49817 & ~n49950;
  assign n49953 = ~n49951 & ~n49952;
  assign n49954 = ~n49813 & n49953;
  assign n49955 = n49813 & ~n49953;
  assign n49956 = ~n49954 & ~n49955;
  assign n49957 = n49808 & n49956;
  assign n49958 = ~n49808 & ~n49956;
  assign n49959 = ~n49957 & ~n49958;
  assign n49960 = n49805 & n49959;
  assign n49961 = ~n49805 & ~n49959;
  assign n49962 = ~n49960 & ~n49961;
  assign n49963 = P4_DATAO_REG_14_ & n44382;
  assign n49964 = ~n49962 & ~n49963;
  assign n49965 = n49962 & n49963;
  assign n49966 = ~n49964 & ~n49965;
  assign n49967 = n49801 & n49966;
  assign n49968 = ~n49801 & ~n49966;
  assign n49969 = ~n49967 & ~n49968;
  assign n49970 = n49798 & n49969;
  assign n49971 = ~n49798 & ~n49969;
  assign n49972 = ~n49970 & ~n49971;
  assign n49973 = P4_DATAO_REG_13_ & n44380;
  assign n49974 = P4_DATAO_REG_12_ & n44378;
  assign n49975 = n49973 & ~n49974;
  assign n49976 = ~n49973 & n49974;
  assign n49977 = ~n49975 & ~n49976;
  assign n49978 = ~n49972 & n49977;
  assign n49979 = n49972 & ~n49977;
  assign n49980 = ~n49978 & ~n49979;
  assign n49981 = n49794 & n49980;
  assign n49982 = ~n49794 & ~n49980;
  assign n49983 = ~n49981 & ~n49982;
  assign n49984 = n49791 & n49983;
  assign n49985 = ~n49791 & ~n49983;
  assign n49986 = ~n49984 & ~n49985;
  assign n49987 = n49787 & n49986;
  assign n49988 = ~n49787 & ~n49986;
  assign n49989 = ~n49987 & ~n49988;
  assign n49990 = n49786 & n49989;
  assign n49991 = ~n49786 & ~n49989;
  assign n49992 = ~n49990 & ~n49991;
  assign n49993 = P4_DATAO_REG_10_ & n44374;
  assign n49994 = P4_DATAO_REG_9_ & n46777;
  assign n49995 = n49993 & ~n49994;
  assign n49996 = ~n49993 & n49994;
  assign n49997 = ~n49995 & ~n49996;
  assign n49998 = P4_DATAO_REG_8_ & n44372;
  assign n49999 = ~n49997 & ~n49998;
  assign n50000 = n49997 & n49998;
  assign n50001 = ~n49999 & ~n50000;
  assign n50002 = ~n49992 & n50001;
  assign n50003 = n49992 & ~n50001;
  assign n50004 = ~n50002 & ~n50003;
  assign n50005 = n49398 & ~n49680;
  assign n50006 = ~n49397 & ~n49680;
  assign n50007 = ~n49682 & ~n50005;
  assign n50008 = ~n50006 & n50007;
  assign n50009 = ~n50004 & ~n50008;
  assign n50010 = n50004 & n50008;
  assign n50011 = ~n50009 & ~n50010;
  assign n50012 = n49783 & n50011;
  assign n50013 = ~n49783 & ~n50011;
  assign n50014 = ~n50012 & ~n50013;
  assign n50015 = P4_DATAO_REG_7_ & n47277;
  assign n50016 = ~n50014 & ~n50015;
  assign n50017 = n50014 & n50015;
  assign n50018 = ~n50016 & ~n50017;
  assign n50019 = n49781 & n50018;
  assign n50020 = ~n49781 & ~n50018;
  assign n50021 = ~n50019 & ~n50020;
  assign n50022 = n49777 & n50021;
  assign n50023 = ~n49777 & ~n50021;
  assign n50024 = ~n50022 & ~n50023;
  assign n50025 = P4_DATAO_REG_6_ & n47275;
  assign n50026 = P4_DATAO_REG_5_ & n47273;
  assign n50027 = n50025 & ~n50026;
  assign n50028 = ~n50025 & n50026;
  assign n50029 = ~n50027 & ~n50028;
  assign n50030 = ~n50024 & n50029;
  assign n50031 = n50024 & ~n50029;
  assign n50032 = ~n50030 & ~n50031;
  assign n50033 = n49775 & n50032;
  assign n50034 = ~n49775 & ~n50032;
  assign n50035 = ~n50033 & ~n50034;
  assign n50036 = n49774 & n50035;
  assign n50037 = ~n49774 & ~n50035;
  assign n50038 = ~n50036 & ~n50037;
  assign n50039 = P4_DATAO_REG_3_ & n47269;
  assign n50040 = ~n50038 & ~n50039;
  assign n50041 = n50038 & n50039;
  assign n50042 = ~n50040 & ~n50041;
  assign n50043 = ~n49367 & ~n49715;
  assign n50044 = ~n49366 & ~n50043;
  assign n50045 = ~n49724 & ~n50044;
  assign n50046 = ~n50042 & ~n50045;
  assign n50047 = n50042 & n50045;
  assign n50048 = ~n50046 & ~n50047;
  assign n50049 = n49770 & n50048;
  assign n50050 = ~n49770 & ~n50048;
  assign n50051 = ~n50049 & ~n50050;
  assign n50052 = ~n49766 & n50051;
  assign n50053 = n49766 & ~n50051;
  assign n50054 = ~n50052 & ~n50053;
  assign n50055 = n49760 & n50054;
  assign n50056 = ~n49760 & ~n50054;
  assign n50057 = ~n50055 & ~n50056;
  assign n50058 = n49757 & n50057;
  assign n50059 = ~n49757 & ~n50057;
  assign n50060 = ~n50058 & ~n50059;
  assign n50061 = SEL & DIN_31_;
  assign n50062 = ~P4_DATAO_REG_0_ & n50061;
  assign n50063 = P4_DATAO_REG_0_ & n49761;
  assign n50064 = n47270 & ~n49280;
  assign n50065 = ~n47270 & n49280;
  assign n50066 = ~n50064 & ~n50065;
  assign n50067 = n49354 & ~n50066;
  assign n50068 = ~n47270 & n49271;
  assign n50069 = ~n47270 & ~n49278;
  assign n50070 = ~n49279 & ~n50068;
  assign n50071 = ~n50069 & n50070;
  assign n50072 = ~n49354 & ~n50071;
  assign n50073 = ~n50067 & ~n50072;
  assign n50074 = P4_DATAO_REG_0_ & n47267;
  assign n50075 = n50073 & ~n50074;
  assign n50076 = ~n49282 & ~n49332;
  assign n50077 = ~n49351 & n50076;
  assign n50078 = ~n49353 & ~n50077;
  assign n50079 = n49346 & ~n50078;
  assign n50080 = ~n49282 & n49352;
  assign n50081 = ~n49353 & ~n50080;
  assign n50082 = ~n49346 & n50081;
  assign n50083 = ~n50079 & ~n50082;
  assign n50084 = P4_DATAO_REG_0_ & n47271;
  assign n50085 = P4_DATAO_REG_0_ & n47273;
  assign n50086 = P4_DATAO_REG_0_ & n47275;
  assign n50087 = ~n49301 & ~n49307;
  assign n50088 = n49306 & ~n50087;
  assign n50089 = ~n49306 & n50087;
  assign n50090 = ~n50088 & ~n50089;
  assign n50091 = n50086 & ~n50090;
  assign n50092 = ~n50086 & n50090;
  assign n50093 = P4_DATAO_REG_0_ & n47277;
  assign n50094 = n44373 & ~n47253;
  assign n50095 = ~n47078 & ~n47253;
  assign n50096 = ~n47079 & ~n50094;
  assign n50097 = ~n50095 & n50096;
  assign n50098 = n50093 & ~n50097;
  assign n50099 = ~n49288 & ~n49291;
  assign n50100 = n49288 & n49291;
  assign n50101 = ~n50099 & ~n50100;
  assign n50102 = n49298 & n50101;
  assign n50103 = ~n49298 & n50099;
  assign n50104 = n49288 & n49299;
  assign n50105 = ~n50102 & ~n50103;
  assign n50106 = ~n50104 & n50105;
  assign n50107 = ~n50097 & n50106;
  assign n50108 = n50093 & n50106;
  assign n50109 = ~n50098 & ~n50107;
  assign n50110 = ~n50108 & n50109;
  assign n50111 = ~n50092 & ~n50110;
  assign n50112 = ~n50091 & ~n50111;
  assign n50113 = n50085 & ~n50112;
  assign n50114 = ~n49283 & n49314;
  assign n50115 = ~n49315 & ~n50114;
  assign n50116 = n49309 & ~n50115;
  assign n50117 = ~n49283 & ~n49314;
  assign n50118 = ~n49309 & n50117;
  assign n50119 = n49310 & n49314;
  assign n50120 = ~n50116 & ~n50118;
  assign n50121 = ~n50119 & n50120;
  assign n50122 = ~n50085 & ~n50091;
  assign n50123 = ~n50111 & n50122;
  assign n50124 = n50121 & ~n50123;
  assign n50125 = ~n50113 & ~n50124;
  assign n50126 = n50084 & ~n50125;
  assign n50127 = n49330 & ~n49331;
  assign n50128 = n49318 & n50127;
  assign n50129 = ~n49318 & n49332;
  assign n50130 = ~n50128 & ~n50129;
  assign n50131 = n49318 & ~n49331;
  assign n50132 = ~n49318 & n49331;
  assign n50133 = ~n50131 & ~n50132;
  assign n50134 = ~n49330 & n50133;
  assign n50135 = n50130 & ~n50134;
  assign n50136 = n50084 & ~n50135;
  assign n50137 = ~n50125 & ~n50135;
  assign n50138 = ~n50126 & ~n50136;
  assign n50139 = ~n50137 & n50138;
  assign n50140 = n50083 & ~n50139;
  assign n50141 = P4_DATAO_REG_0_ & n47269;
  assign n50142 = n50083 & n50141;
  assign n50143 = ~n50139 & n50141;
  assign n50144 = ~n50140 & ~n50142;
  assign n50145 = ~n50143 & n50144;
  assign n50146 = ~n50075 & ~n50145;
  assign n50147 = ~n50073 & n50074;
  assign n50148 = ~n50146 & ~n50147;
  assign n50149 = n50063 & ~n50148;
  assign n50150 = ~n50063 & ~n50074;
  assign n50151 = n50073 & n50150;
  assign n50152 = n49357 & n49753;
  assign n50153 = ~n50140 & ~n50143;
  assign n50154 = ~n50063 & n50153;
  assign n50155 = ~n50142 & n50154;
  assign n50156 = ~n50147 & n50155;
  assign n50157 = ~n50151 & ~n50152;
  assign n50158 = ~n50156 & n50157;
  assign n50159 = ~n47268 & ~n49753;
  assign n50160 = ~n49356 & n50159;
  assign n50161 = n47268 & n49753;
  assign n50162 = ~n50159 & ~n50161;
  assign n50163 = n49356 & n50162;
  assign n50164 = ~n50160 & ~n50163;
  assign n50165 = n50158 & n50164;
  assign n50166 = ~n50062 & ~n50149;
  assign n50167 = ~n50165 & n50166;
  assign n50168 = ~n50060 & ~n50167;
  assign n50169 = n50060 & n50167;
  assign n50170 = P4_DATAO_REG_31_ & ~n50061;
  assign n50171 = ~P4_DATAO_REG_31_ & n50061;
  assign n50172 = ~n50170 & ~n50171;
  assign n50173 = ~n50168 & ~n50169;
  assign n50174 = n50172 & n50173;
  assign n50175 = ~n50063 & ~n50147;
  assign n50176 = ~n50146 & n50175;
  assign n50177 = ~n50152 & n50164;
  assign n50178 = ~n50176 & n50177;
  assign n50179 = n50166 & ~n50178;
  assign n50180 = ~n50060 & ~n50179;
  assign n50181 = n50060 & n50179;
  assign n50182 = ~n50180 & ~n50181;
  assign n50183 = ~n50172 & ~n50182;
  assign n50184 = ~n50174 & ~n50183;
  assign n50185 = ~n12460 & ~n50184;
  assign n50186 = ~n47266 & ~n50185;
  assign n50187 = n47260 & ~n50186;
  assign n50188 = n47265 & ~n50187;
  assign n50189 = ~n44086 & n47265;
  assign n8106 = ~n50188 & ~n50189;
  assign n50191 = P1_P1_INSTQUEUE_REG_15__6_ & ~n44092;
  assign n50192 = P1_BUF1_REG_6_ & n12460;
  assign n50193 = n44103 & ~n44280;
  assign n50194 = ~n44103 & n44280;
  assign n50195 = ~n50193 & ~n50194;
  assign n50196 = n44221 & ~n50195;
  assign n50197 = ~n44103 & ~n44280;
  assign n50198 = ~n44221 & n50197;
  assign n50199 = n44222 & n44280;
  assign n50200 = ~n50196 & ~n50198;
  assign n50201 = ~n50199 & n50200;
  assign n50202 = ~n12460 & ~n50201;
  assign n50203 = ~n50192 & ~n50202;
  assign n50204 = n44042 & ~n50203;
  assign n50205 = n44100 & n50204;
  assign n50206 = ~n43432 & n44094;
  assign n50207 = n44037 & n50206;
  assign n50208 = P1_BUF1_REG_22_ & n12460;
  assign n50209 = n47081 & ~n47250;
  assign n50210 = ~n47081 & n47250;
  assign n50211 = ~n50209 & ~n50210;
  assign n50212 = n47241 & ~n50211;
  assign n50213 = ~n47081 & ~n47250;
  assign n50214 = ~n47241 & n50213;
  assign n50215 = n47242 & n47250;
  assign n50216 = ~n50212 & ~n50214;
  assign n50217 = ~n50215 & n50216;
  assign n50218 = ~n12460 & ~n50217;
  assign n50219 = ~n50208 & ~n50218;
  assign n50220 = n47260 & ~n50219;
  assign n50221 = n44088 & n50220;
  assign n50222 = P1_BUF1_REG_30_ & n12460;
  assign n50223 = n50063 & ~n50177;
  assign n50224 = ~n50063 & n50177;
  assign n50225 = ~n50223 & ~n50224;
  assign n50226 = n50148 & ~n50225;
  assign n50227 = ~n50063 & ~n50177;
  assign n50228 = ~n50148 & n50227;
  assign n50229 = n50149 & n50177;
  assign n50230 = ~n50226 & ~n50228;
  assign n50231 = ~n50229 & n50230;
  assign n50232 = ~n12460 & ~n50231;
  assign n50233 = ~n50222 & ~n50232;
  assign n50234 = n47260 & ~n50233;
  assign n50235 = n44086 & n50234;
  assign n50236 = ~n50191 & ~n50205;
  assign n50237 = ~n50207 & n50236;
  assign n50238 = ~n50221 & n50237;
  assign n8111 = n50235 | ~n50238;
  assign n50240 = P1_P1_INSTQUEUE_REG_15__5_ & ~n44092;
  assign n50241 = P1_BUF1_REG_5_ & n12460;
  assign n50242 = ~n44105 & ~n44183;
  assign n50243 = n44105 & n44183;
  assign n50244 = ~n50242 & ~n50243;
  assign n50245 = n44219 & ~n50244;
  assign n50246 = ~n44184 & ~n44185;
  assign n50247 = ~n44219 & ~n50246;
  assign n50248 = ~n50245 & ~n50247;
  assign n50249 = ~n12460 & ~n50248;
  assign n50250 = ~n50241 & ~n50249;
  assign n50251 = n44042 & ~n50250;
  assign n50252 = n44100 & n50251;
  assign n50253 = ~n43401 & n44094;
  assign n50254 = n44037 & n50253;
  assign n50255 = P1_BUF1_REG_21_ & n12460;
  assign n50256 = ~n47082 & ~n47086;
  assign n50257 = n47082 & n47086;
  assign n50258 = ~n50256 & ~n50257;
  assign n50259 = n47239 & ~n50258;
  assign n50260 = ~n47239 & n50258;
  assign n50261 = ~n50259 & ~n50260;
  assign n50262 = ~n12460 & ~n50261;
  assign n50263 = ~n50255 & ~n50262;
  assign n50264 = n47260 & ~n50263;
  assign n50265 = n44088 & n50264;
  assign n50266 = P1_BUF1_REG_29_ & n12460;
  assign n50267 = ~n50073 & ~n50074;
  assign n50268 = n50073 & n50074;
  assign n50269 = ~n50267 & ~n50268;
  assign n50270 = n50145 & ~n50269;
  assign n50271 = ~n50075 & ~n50147;
  assign n50272 = ~n50145 & ~n50271;
  assign n50273 = ~n50270 & ~n50272;
  assign n50274 = ~n12460 & ~n50273;
  assign n50275 = ~n50266 & ~n50274;
  assign n50276 = n47260 & ~n50275;
  assign n50277 = n44086 & n50276;
  assign n50278 = ~n50240 & ~n50252;
  assign n50279 = ~n50254 & n50278;
  assign n50280 = ~n50265 & n50279;
  assign n8116 = n50277 | ~n50280;
  assign n50282 = P1_P1_INSTQUEUE_REG_15__4_ & ~n44092;
  assign n50283 = P1_BUF1_REG_4_ & n12460;
  assign n50284 = n44186 & ~n44216;
  assign n50285 = ~n44186 & n44216;
  assign n50286 = ~n50284 & ~n50285;
  assign n50287 = n44207 & ~n50286;
  assign n50288 = ~n44186 & ~n44216;
  assign n50289 = ~n44207 & n50288;
  assign n50290 = n44208 & n44216;
  assign n50291 = ~n50287 & ~n50289;
  assign n50292 = ~n50290 & n50291;
  assign n50293 = ~n12460 & ~n50292;
  assign n50294 = ~n50283 & ~n50293;
  assign n50295 = n44042 & ~n50294;
  assign n50296 = n44100 & n50295;
  assign n50297 = ~n43464 & n44094;
  assign n50298 = n44037 & n50297;
  assign n50299 = P1_BUF1_REG_20_ & n12460;
  assign n50300 = ~n47089 & ~n47236;
  assign n50301 = n47089 & n47236;
  assign n50302 = ~n50300 & ~n50301;
  assign n50303 = n47229 & n50302;
  assign n50304 = ~n47229 & n50300;
  assign n50305 = n47230 & n47236;
  assign n50306 = ~n50303 & ~n50304;
  assign n50307 = ~n50305 & n50306;
  assign n50308 = ~n12460 & ~n50307;
  assign n50309 = ~n50299 & ~n50308;
  assign n50310 = n47260 & ~n50309;
  assign n50311 = n44088 & n50310;
  assign n50312 = P1_BUF1_REG_28_ & n12460;
  assign n50313 = n50139 & ~n50141;
  assign n50314 = ~n50143 & ~n50313;
  assign n50315 = ~n50083 & n50314;
  assign n50316 = n50083 & n50313;
  assign n50317 = ~n50139 & n50142;
  assign n50318 = ~n50315 & ~n50316;
  assign n50319 = ~n50317 & n50318;
  assign n50320 = ~n12460 & ~n50319;
  assign n50321 = ~n50312 & ~n50320;
  assign n50322 = n47260 & ~n50321;
  assign n50323 = n44086 & n50322;
  assign n50324 = ~n50282 & ~n50296;
  assign n50325 = ~n50298 & n50324;
  assign n50326 = ~n50311 & n50325;
  assign n8121 = n50323 | ~n50326;
  assign n50328 = P1_P1_INSTQUEUE_REG_15__3_ & ~n44092;
  assign n50329 = P1_BUF1_REG_3_ & n12460;
  assign n50330 = ~n44187 & ~n44191;
  assign n50331 = n44187 & n44191;
  assign n50332 = ~n50330 & ~n50331;
  assign n50333 = n44205 & ~n50332;
  assign n50334 = ~n44192 & ~n44193;
  assign n50335 = ~n44205 & ~n50334;
  assign n50336 = ~n50333 & ~n50335;
  assign n50337 = ~n12460 & ~n50336;
  assign n50338 = ~n50329 & ~n50337;
  assign n50339 = n44042 & ~n50338;
  assign n50340 = n44100 & n50339;
  assign n50341 = ~n43526 & n44094;
  assign n50342 = n44037 & n50341;
  assign n50343 = P1_BUF1_REG_19_ & n12460;
  assign n50344 = ~n47090 & ~n47094;
  assign n50345 = n47090 & n47094;
  assign n50346 = ~n50344 & ~n50345;
  assign n50347 = n47227 & ~n50346;
  assign n50348 = ~n47095 & ~n47096;
  assign n50349 = ~n47227 & ~n50348;
  assign n50350 = ~n50347 & ~n50349;
  assign n50351 = ~n12460 & ~n50350;
  assign n50352 = ~n50343 & ~n50351;
  assign n50353 = n47260 & ~n50352;
  assign n50354 = n44088 & n50353;
  assign n50355 = P1_BUF1_REG_27_ & n12460;
  assign n50356 = ~n50084 & n50135;
  assign n50357 = ~n50136 & ~n50356;
  assign n50358 = n50125 & n50357;
  assign n50359 = ~n50125 & ~n50357;
  assign n50360 = ~n50358 & ~n50359;
  assign n50361 = ~n12460 & ~n50360;
  assign n50362 = ~n50355 & ~n50361;
  assign n50363 = n47260 & ~n50362;
  assign n50364 = n44086 & n50363;
  assign n50365 = ~n50328 & ~n50340;
  assign n50366 = ~n50342 & n50365;
  assign n50367 = ~n50354 & n50366;
  assign n8126 = n50364 | ~n50367;
  assign n50369 = P1_P1_INSTQUEUE_REG_15__2_ & ~n44092;
  assign n50370 = P1_BUF1_REG_2_ & n12460;
  assign n50371 = n44197 & ~n44203;
  assign n50372 = ~n44197 & n44203;
  assign n50373 = ~n50371 & ~n50372;
  assign n50374 = ~n44196 & n50373;
  assign n50375 = n44196 & n50372;
  assign n50376 = n44198 & ~n44203;
  assign n50377 = ~n50374 & ~n50375;
  assign n50378 = ~n50376 & n50377;
  assign n50379 = ~n12460 & ~n50378;
  assign n50380 = ~n50370 & ~n50379;
  assign n50381 = n44042 & ~n50380;
  assign n50382 = n44100 & n50381;
  assign n50383 = ~n43557 & n44094;
  assign n50384 = n44037 & n50383;
  assign n50385 = P1_BUF1_REG_18_ & n12460;
  assign n50386 = n47097 & ~n47224;
  assign n50387 = ~n47097 & n47224;
  assign n50388 = ~n50386 & ~n50387;
  assign n50389 = n47215 & ~n50388;
  assign n50390 = ~n47097 & ~n47224;
  assign n50391 = ~n47215 & n50390;
  assign n50392 = n47216 & n47224;
  assign n50393 = ~n50389 & ~n50391;
  assign n50394 = ~n50392 & n50393;
  assign n50395 = ~n12460 & ~n50394;
  assign n50396 = ~n50385 & ~n50395;
  assign n50397 = n47260 & ~n50396;
  assign n50398 = n44088 & n50397;
  assign n50399 = P1_BUF1_REG_26_ & n12460;
  assign n50400 = n50085 & ~n50121;
  assign n50401 = ~n50085 & n50121;
  assign n50402 = ~n50400 & ~n50401;
  assign n50403 = n50112 & ~n50402;
  assign n50404 = ~n50085 & ~n50121;
  assign n50405 = ~n50112 & n50404;
  assign n50406 = n50113 & n50121;
  assign n50407 = ~n50403 & ~n50405;
  assign n50408 = ~n50406 & n50407;
  assign n50409 = ~n12460 & ~n50408;
  assign n50410 = ~n50399 & ~n50409;
  assign n50411 = n47260 & ~n50410;
  assign n50412 = n44086 & n50411;
  assign n50413 = ~n50369 & ~n50382;
  assign n50414 = ~n50384 & n50413;
  assign n50415 = ~n50398 & n50414;
  assign n8131 = n50412 | ~n50415;
  assign n50417 = P1_P1_INSTQUEUE_REG_15__1_ & ~n44092;
  assign n50418 = P1_BUF1_REG_1_ & n12460;
  assign n50419 = P4_DATAO_REG_1_ & n44112;
  assign n50420 = P4_DATAO_REG_0_ & n44110;
  assign n50421 = n50419 & ~n50420;
  assign n50422 = ~n50419 & n50420;
  assign n50423 = ~n50421 & ~n50422;
  assign n50424 = ~n12460 & ~n50423;
  assign n50425 = ~n50418 & ~n50424;
  assign n50426 = n44042 & ~n50425;
  assign n50427 = n44100 & n50426;
  assign n50428 = ~n43592 & n44094;
  assign n50429 = n44037 & n50428;
  assign n50430 = P1_BUF1_REG_17_ & n12460;
  assign n50431 = ~n47205 & ~n47213;
  assign n50432 = n47212 & n50431;
  assign n50433 = ~n47212 & ~n50431;
  assign n50434 = ~n50432 & ~n50433;
  assign n50435 = ~n12460 & ~n50434;
  assign n50436 = ~n50430 & ~n50435;
  assign n50437 = n47260 & ~n50436;
  assign n50438 = n44088 & n50437;
  assign n50439 = P1_BUF1_REG_25_ & n12460;
  assign n50440 = ~n50086 & ~n50090;
  assign n50441 = n50086 & n50090;
  assign n50442 = ~n50440 & ~n50441;
  assign n50443 = n50110 & ~n50442;
  assign n50444 = ~n50091 & ~n50092;
  assign n50445 = ~n50110 & ~n50444;
  assign n50446 = ~n50443 & ~n50445;
  assign n50447 = ~n12460 & ~n50446;
  assign n50448 = ~n50439 & ~n50447;
  assign n50449 = n47260 & ~n50448;
  assign n50450 = n44086 & n50449;
  assign n50451 = ~n50417 & ~n50427;
  assign n50452 = ~n50429 & n50451;
  assign n50453 = ~n50438 & n50452;
  assign n8136 = n50450 | ~n50453;
  assign n50455 = P1_P1_INSTQUEUE_REG_15__0_ & ~n44092;
  assign n50456 = P1_BUF1_REG_0_ & n12460;
  assign n50457 = ~n12460 & n44195;
  assign n50458 = ~n50456 & ~n50457;
  assign n50459 = n44042 & ~n50458;
  assign n50460 = n44100 & n50459;
  assign n50461 = ~n43623 & n44094;
  assign n50462 = n44037 & n50461;
  assign n50463 = P1_BUF1_REG_16_ & n12460;
  assign n50464 = n47107 & ~n47202;
  assign n50465 = ~n47107 & n47202;
  assign n50466 = ~n50464 & ~n50465;
  assign n50467 = ~n47106 & n50466;
  assign n50468 = n47106 & n50465;
  assign n50469 = n47108 & ~n47202;
  assign n50470 = ~n50467 & ~n50468;
  assign n50471 = ~n50469 & n50470;
  assign n50472 = ~n12460 & ~n50471;
  assign n50473 = ~n50463 & ~n50472;
  assign n50474 = n47260 & ~n50473;
  assign n50475 = n44088 & n50474;
  assign n50476 = P1_BUF1_REG_24_ & n12460;
  assign n50477 = n50093 & ~n50106;
  assign n50478 = ~n50093 & n50106;
  assign n50479 = ~n50477 & ~n50478;
  assign n50480 = n50097 & ~n50479;
  assign n50481 = ~n50093 & ~n50106;
  assign n50482 = ~n50097 & n50481;
  assign n50483 = n50098 & n50106;
  assign n50484 = ~n50480 & ~n50482;
  assign n50485 = ~n50483 & n50484;
  assign n50486 = ~n12460 & ~n50485;
  assign n50487 = ~n50476 & ~n50486;
  assign n50488 = n47260 & ~n50487;
  assign n50489 = n44086 & n50488;
  assign n50490 = ~n50455 & ~n50460;
  assign n50491 = ~n50462 & n50490;
  assign n50492 = ~n50475 & n50491;
  assign n8141 = n50489 | ~n50492;
  assign n50494 = P1_P1_INSTQUEUEWR_ADDR_REG_3_ & P1_P1_INSTQUEUEWR_ADDR_REG_1_;
  assign n50495 = P1_P1_INSTQUEUEWR_ADDR_REG_2_ & ~P1_P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n50496 = n50494 & n50495;
  assign n50497 = P1_P1_STATE2_REG_3_ & ~n50496;
  assign n50498 = n44042 & ~n50497;
  assign n50499 = n44050 & n44060;
  assign n50500 = ~n50496 & ~n50499;
  assign n50501 = P1_P1_INSTQUEUEWR_ADDR_REG_0_ & ~n44065;
  assign n50502 = n44085 & n50501;
  assign n50503 = n44063 & n44087;
  assign n50504 = ~n50502 & ~n50503;
  assign n50505 = n44059 & ~n50504;
  assign n50506 = n50500 & ~n50505;
  assign n50507 = n50498 & ~n50506;
  assign n50508 = P1_P1_INSTQUEUE_REG_14__7_ & ~n50507;
  assign n50509 = n44095 & n50496;
  assign n50510 = n44097 & n50504;
  assign n50511 = n44059 & ~n50510;
  assign n50512 = ~n50500 & ~n50511;
  assign n50513 = n44369 & n50512;
  assign n50514 = n47261 & n50503;
  assign n50515 = ~n50508 & ~n50509;
  assign n50516 = ~n50513 & n50515;
  assign n50517 = ~n50514 & n50516;
  assign n50518 = ~n50187 & n50517;
  assign n50519 = ~n50502 & n50517;
  assign n8146 = ~n50518 & ~n50519;
  assign n50521 = P1_P1_INSTQUEUE_REG_14__6_ & ~n50507;
  assign n50522 = n50204 & n50512;
  assign n50523 = n50206 & n50496;
  assign n50524 = n50220 & n50503;
  assign n50525 = n50234 & n50502;
  assign n50526 = ~n50521 & ~n50522;
  assign n50527 = ~n50523 & n50526;
  assign n50528 = ~n50524 & n50527;
  assign n8151 = n50525 | ~n50528;
  assign n50530 = P1_P1_INSTQUEUE_REG_14__5_ & ~n50507;
  assign n50531 = n50251 & n50512;
  assign n50532 = n50253 & n50496;
  assign n50533 = n50264 & n50503;
  assign n50534 = n50276 & n50502;
  assign n50535 = ~n50530 & ~n50531;
  assign n50536 = ~n50532 & n50535;
  assign n50537 = ~n50533 & n50536;
  assign n8156 = n50534 | ~n50537;
  assign n50539 = P1_P1_INSTQUEUE_REG_14__4_ & ~n50507;
  assign n50540 = n50295 & n50512;
  assign n50541 = n50297 & n50496;
  assign n50542 = n50310 & n50503;
  assign n50543 = n50322 & n50502;
  assign n50544 = ~n50539 & ~n50540;
  assign n50545 = ~n50541 & n50544;
  assign n50546 = ~n50542 & n50545;
  assign n8161 = n50543 | ~n50546;
  assign n50548 = P1_P1_INSTQUEUE_REG_14__3_ & ~n50507;
  assign n50549 = n50339 & n50512;
  assign n50550 = n50341 & n50496;
  assign n50551 = n50353 & n50503;
  assign n50552 = n50363 & n50502;
  assign n50553 = ~n50548 & ~n50549;
  assign n50554 = ~n50550 & n50553;
  assign n50555 = ~n50551 & n50554;
  assign n8166 = n50552 | ~n50555;
  assign n50557 = P1_P1_INSTQUEUE_REG_14__2_ & ~n50507;
  assign n50558 = n50381 & n50512;
  assign n50559 = n50383 & n50496;
  assign n50560 = n50397 & n50503;
  assign n50561 = n50411 & n50502;
  assign n50562 = ~n50557 & ~n50558;
  assign n50563 = ~n50559 & n50562;
  assign n50564 = ~n50560 & n50563;
  assign n8171 = n50561 | ~n50564;
  assign n50566 = P1_P1_INSTQUEUE_REG_14__1_ & ~n50507;
  assign n50567 = n50426 & n50512;
  assign n50568 = n50428 & n50496;
  assign n50569 = n50437 & n50503;
  assign n50570 = n50449 & n50502;
  assign n50571 = ~n50566 & ~n50567;
  assign n50572 = ~n50568 & n50571;
  assign n50573 = ~n50569 & n50572;
  assign n8176 = n50570 | ~n50573;
  assign n50575 = P1_P1_INSTQUEUE_REG_14__0_ & ~n50507;
  assign n50576 = n50459 & n50512;
  assign n50577 = n50461 & n50496;
  assign n50578 = n50474 & n50503;
  assign n50579 = n50488 & n50502;
  assign n50580 = ~n50575 & ~n50576;
  assign n50581 = ~n50577 & n50580;
  assign n50582 = ~n50578 & n50581;
  assign n8181 = n50579 | ~n50582;
  assign n50584 = P1_P1_INSTQUEUEWR_ADDR_REG_3_ & P1_P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n50585 = n44051 & n50584;
  assign n50586 = P1_P1_STATE2_REG_3_ & ~n50585;
  assign n50587 = n44042 & ~n50586;
  assign n50588 = n44050 & n44061;
  assign n50589 = ~n50585 & ~n50588;
  assign n50590 = ~P1_P1_INSTQUEUEWR_ADDR_REG_0_ & n44065;
  assign n50591 = n44085 & n50590;
  assign n50592 = n44064 & n44087;
  assign n50593 = ~n50591 & ~n50592;
  assign n50594 = n44059 & ~n50593;
  assign n50595 = n50589 & ~n50594;
  assign n50596 = n50587 & ~n50595;
  assign n50597 = P1_P1_INSTQUEUE_REG_13__7_ & ~n50596;
  assign n50598 = n44095 & n50585;
  assign n50599 = n44097 & n50593;
  assign n50600 = n44059 & ~n50599;
  assign n50601 = ~n50589 & ~n50600;
  assign n50602 = n44369 & n50601;
  assign n50603 = n47261 & n50592;
  assign n50604 = ~n50597 & ~n50598;
  assign n50605 = ~n50602 & n50604;
  assign n50606 = ~n50603 & n50605;
  assign n50607 = ~n50187 & n50606;
  assign n50608 = ~n50591 & n50606;
  assign n8186 = ~n50607 & ~n50608;
  assign n50610 = P1_P1_INSTQUEUE_REG_13__6_ & ~n50596;
  assign n50611 = n50204 & n50601;
  assign n50612 = n50206 & n50585;
  assign n50613 = n50220 & n50592;
  assign n50614 = n50234 & n50591;
  assign n50615 = ~n50610 & ~n50611;
  assign n50616 = ~n50612 & n50615;
  assign n50617 = ~n50613 & n50616;
  assign n8191 = n50614 | ~n50617;
  assign n50619 = P1_P1_INSTQUEUE_REG_13__5_ & ~n50596;
  assign n50620 = n50251 & n50601;
  assign n50621 = n50253 & n50585;
  assign n50622 = n50264 & n50592;
  assign n50623 = n50276 & n50591;
  assign n50624 = ~n50619 & ~n50620;
  assign n50625 = ~n50621 & n50624;
  assign n50626 = ~n50622 & n50625;
  assign n8196 = n50623 | ~n50626;
  assign n50628 = P1_P1_INSTQUEUE_REG_13__4_ & ~n50596;
  assign n50629 = n50295 & n50601;
  assign n50630 = n50297 & n50585;
  assign n50631 = n50310 & n50592;
  assign n50632 = n50322 & n50591;
  assign n50633 = ~n50628 & ~n50629;
  assign n50634 = ~n50630 & n50633;
  assign n50635 = ~n50631 & n50634;
  assign n8201 = n50632 | ~n50635;
  assign n50637 = P1_P1_INSTQUEUE_REG_13__3_ & ~n50596;
  assign n50638 = n50339 & n50601;
  assign n50639 = n50341 & n50585;
  assign n50640 = n50353 & n50592;
  assign n50641 = n50363 & n50591;
  assign n50642 = ~n50637 & ~n50638;
  assign n50643 = ~n50639 & n50642;
  assign n50644 = ~n50640 & n50643;
  assign n8206 = n50641 | ~n50644;
  assign n50646 = P1_P1_INSTQUEUE_REG_13__2_ & ~n50596;
  assign n50647 = n50381 & n50601;
  assign n50648 = n50383 & n50585;
  assign n50649 = n50397 & n50592;
  assign n50650 = n50411 & n50591;
  assign n50651 = ~n50646 & ~n50647;
  assign n50652 = ~n50648 & n50651;
  assign n50653 = ~n50649 & n50652;
  assign n8211 = n50650 | ~n50653;
  assign n50655 = P1_P1_INSTQUEUE_REG_13__1_ & ~n50596;
  assign n50656 = n50426 & n50601;
  assign n50657 = n50428 & n50585;
  assign n50658 = n50437 & n50592;
  assign n50659 = n50449 & n50591;
  assign n50660 = ~n50655 & ~n50656;
  assign n50661 = ~n50657 & n50660;
  assign n50662 = ~n50658 & n50661;
  assign n8216 = n50659 | ~n50662;
  assign n50664 = P1_P1_INSTQUEUE_REG_13__0_ & ~n50596;
  assign n50665 = n50459 & n50601;
  assign n50666 = n50461 & n50585;
  assign n50667 = n50474 & n50592;
  assign n50668 = n50488 & n50591;
  assign n50669 = ~n50664 & ~n50665;
  assign n50670 = ~n50666 & n50669;
  assign n50671 = ~n50667 & n50670;
  assign n8221 = n50668 | ~n50671;
  assign n50673 = P1_P1_INSTQUEUEWR_ADDR_REG_3_ & ~P1_P1_INSTQUEUEWR_ADDR_REG_1_;
  assign n50674 = n50495 & n50673;
  assign n50675 = P1_P1_STATE2_REG_3_ & ~n50674;
  assign n50676 = n44042 & ~n50675;
  assign n50677 = P1_P1_INSTQUEUEWR_ADDR_REG_0_ & n44065;
  assign n50678 = n44085 & n50677;
  assign n50679 = ~P1_P1_INSTQUEUEWR_ADDR_REG_0_ & n44062;
  assign n50680 = n44087 & n50679;
  assign n50681 = ~n50678 & ~n50680;
  assign n50682 = n44059 & ~n50681;
  assign n50683 = n44050 & n44053;
  assign n50684 = ~n50682 & ~n50683;
  assign n50685 = n50676 & ~n50684;
  assign n50686 = P1_P1_INSTQUEUE_REG_12__7_ & ~n50685;
  assign n50687 = n44095 & n50674;
  assign n50688 = n44097 & n50681;
  assign n50689 = n44059 & ~n50688;
  assign n50690 = n50683 & ~n50689;
  assign n50691 = n44369 & n50690;
  assign n50692 = n47261 & n50680;
  assign n50693 = ~n50686 & ~n50687;
  assign n50694 = ~n50691 & n50693;
  assign n50695 = ~n50692 & n50694;
  assign n50696 = ~n50187 & n50695;
  assign n50697 = ~n50678 & n50695;
  assign n8226 = ~n50696 & ~n50697;
  assign n50699 = P1_P1_INSTQUEUE_REG_12__6_ & ~n50685;
  assign n50700 = n50204 & n50690;
  assign n50701 = n50206 & n50674;
  assign n50702 = n50220 & n50680;
  assign n50703 = n50234 & n50678;
  assign n50704 = ~n50699 & ~n50700;
  assign n50705 = ~n50701 & n50704;
  assign n50706 = ~n50702 & n50705;
  assign n8231 = n50703 | ~n50706;
  assign n50708 = P1_P1_INSTQUEUE_REG_12__5_ & ~n50685;
  assign n50709 = n50251 & n50690;
  assign n50710 = n50253 & n50674;
  assign n50711 = n50264 & n50680;
  assign n50712 = n50276 & n50678;
  assign n50713 = ~n50708 & ~n50709;
  assign n50714 = ~n50710 & n50713;
  assign n50715 = ~n50711 & n50714;
  assign n8236 = n50712 | ~n50715;
  assign n50717 = P1_P1_INSTQUEUE_REG_12__4_ & ~n50685;
  assign n50718 = n50295 & n50690;
  assign n50719 = n50297 & n50674;
  assign n50720 = n50310 & n50680;
  assign n50721 = n50322 & n50678;
  assign n50722 = ~n50717 & ~n50718;
  assign n50723 = ~n50719 & n50722;
  assign n50724 = ~n50720 & n50723;
  assign n8241 = n50721 | ~n50724;
  assign n50726 = P1_P1_INSTQUEUE_REG_12__3_ & ~n50685;
  assign n50727 = n50339 & n50690;
  assign n50728 = n50341 & n50674;
  assign n50729 = n50353 & n50680;
  assign n50730 = n50363 & n50678;
  assign n50731 = ~n50726 & ~n50727;
  assign n50732 = ~n50728 & n50731;
  assign n50733 = ~n50729 & n50732;
  assign n8246 = n50730 | ~n50733;
  assign n50735 = P1_P1_INSTQUEUE_REG_12__2_ & ~n50685;
  assign n50736 = n50381 & n50690;
  assign n50737 = n50383 & n50674;
  assign n50738 = n50397 & n50680;
  assign n50739 = n50411 & n50678;
  assign n50740 = ~n50735 & ~n50736;
  assign n50741 = ~n50737 & n50740;
  assign n50742 = ~n50738 & n50741;
  assign n8251 = n50739 | ~n50742;
  assign n50744 = P1_P1_INSTQUEUE_REG_12__1_ & ~n50685;
  assign n50745 = n50426 & n50690;
  assign n50746 = n50428 & n50674;
  assign n50747 = n50437 & n50680;
  assign n50748 = n50449 & n50678;
  assign n50749 = ~n50744 & ~n50745;
  assign n50750 = ~n50746 & n50749;
  assign n50751 = ~n50747 & n50750;
  assign n8256 = n50748 | ~n50751;
  assign n50753 = P1_P1_INSTQUEUE_REG_12__0_ & ~n50685;
  assign n50754 = n50459 & n50690;
  assign n50755 = n50461 & n50674;
  assign n50756 = n50474 & n50680;
  assign n50757 = n50488 & n50678;
  assign n50758 = ~n50753 & ~n50754;
  assign n50759 = ~n50755 & n50758;
  assign n50760 = ~n50756 & n50759;
  assign n8261 = n50757 | ~n50760;
  assign n50762 = P1_P1_INSTQUEUEWR_ADDR_REG_3_ & ~P1_P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n50763 = n44035 & n50762;
  assign n50764 = P1_P1_STATE2_REG_3_ & ~n50763;
  assign n50765 = n44042 & ~n50764;
  assign n50766 = n44046 & ~n44049;
  assign n50767 = n44054 & n50766;
  assign n50768 = ~n50763 & ~n50767;
  assign n50769 = n44073 & ~n44084;
  assign n50770 = n44066 & n50769;
  assign n50771 = n44070 & n44079;
  assign n50772 = ~n50770 & ~n50771;
  assign n50773 = n44059 & ~n50772;
  assign n50774 = n50768 & ~n50773;
  assign n50775 = n50765 & ~n50774;
  assign n50776 = P1_P1_INSTQUEUE_REG_11__7_ & ~n50775;
  assign n50777 = n44095 & n50763;
  assign n50778 = n44097 & n50772;
  assign n50779 = n44059 & ~n50778;
  assign n50780 = ~n50768 & ~n50779;
  assign n50781 = n44369 & n50780;
  assign n50782 = n47261 & n50771;
  assign n50783 = ~n50776 & ~n50777;
  assign n50784 = ~n50781 & n50783;
  assign n50785 = ~n50782 & n50784;
  assign n50786 = ~n50187 & n50785;
  assign n50787 = ~n50770 & n50785;
  assign n8266 = ~n50786 & ~n50787;
  assign n50789 = P1_P1_INSTQUEUE_REG_11__6_ & ~n50775;
  assign n50790 = n50204 & n50780;
  assign n50791 = n50206 & n50763;
  assign n50792 = n50220 & n50771;
  assign n50793 = n50234 & n50770;
  assign n50794 = ~n50789 & ~n50790;
  assign n50795 = ~n50791 & n50794;
  assign n50796 = ~n50792 & n50795;
  assign n8271 = n50793 | ~n50796;
  assign n50798 = P1_P1_INSTQUEUE_REG_11__5_ & ~n50775;
  assign n50799 = n50251 & n50780;
  assign n50800 = n50253 & n50763;
  assign n50801 = n50264 & n50771;
  assign n50802 = n50276 & n50770;
  assign n50803 = ~n50798 & ~n50799;
  assign n50804 = ~n50800 & n50803;
  assign n50805 = ~n50801 & n50804;
  assign n8276 = n50802 | ~n50805;
  assign n50807 = P1_P1_INSTQUEUE_REG_11__4_ & ~n50775;
  assign n50808 = n50295 & n50780;
  assign n50809 = n50297 & n50763;
  assign n50810 = n50310 & n50771;
  assign n50811 = n50322 & n50770;
  assign n50812 = ~n50807 & ~n50808;
  assign n50813 = ~n50809 & n50812;
  assign n50814 = ~n50810 & n50813;
  assign n8281 = n50811 | ~n50814;
  assign n50816 = P1_P1_INSTQUEUE_REG_11__3_ & ~n50775;
  assign n50817 = n50339 & n50780;
  assign n50818 = n50341 & n50763;
  assign n50819 = n50353 & n50771;
  assign n50820 = n50363 & n50770;
  assign n50821 = ~n50816 & ~n50817;
  assign n50822 = ~n50818 & n50821;
  assign n50823 = ~n50819 & n50822;
  assign n8286 = n50820 | ~n50823;
  assign n50825 = P1_P1_INSTQUEUE_REG_11__2_ & ~n50775;
  assign n50826 = n50381 & n50780;
  assign n50827 = n50383 & n50763;
  assign n50828 = n50397 & n50771;
  assign n50829 = n50411 & n50770;
  assign n50830 = ~n50825 & ~n50826;
  assign n50831 = ~n50827 & n50830;
  assign n50832 = ~n50828 & n50831;
  assign n8291 = n50829 | ~n50832;
  assign n50834 = P1_P1_INSTQUEUE_REG_11__1_ & ~n50775;
  assign n50835 = n50426 & n50780;
  assign n50836 = n50428 & n50763;
  assign n50837 = n50437 & n50771;
  assign n50838 = n50449 & n50770;
  assign n50839 = ~n50834 & ~n50835;
  assign n50840 = ~n50836 & n50839;
  assign n50841 = ~n50837 & n50840;
  assign n8296 = n50838 | ~n50841;
  assign n50843 = P1_P1_INSTQUEUE_REG_11__0_ & ~n50775;
  assign n50844 = n50459 & n50780;
  assign n50845 = n50461 & n50763;
  assign n50846 = n50474 & n50771;
  assign n50847 = n50488 & n50770;
  assign n50848 = ~n50843 & ~n50844;
  assign n50849 = ~n50845 & n50848;
  assign n50850 = ~n50846 & n50849;
  assign n8301 = n50847 | ~n50850;
  assign n50852 = ~P1_P1_INSTQUEUEWR_ADDR_REG_2_ & ~P1_P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n50853 = n50494 & n50852;
  assign n50854 = P1_P1_STATE2_REG_3_ & ~n50853;
  assign n50855 = n44042 & ~n50854;
  assign n50856 = n44060 & n50766;
  assign n50857 = ~n50853 & ~n50856;
  assign n50858 = n50501 & n50769;
  assign n50859 = n44063 & n44079;
  assign n50860 = ~n50858 & ~n50859;
  assign n50861 = n44059 & ~n50860;
  assign n50862 = n50857 & ~n50861;
  assign n50863 = n50855 & ~n50862;
  assign n50864 = P1_P1_INSTQUEUE_REG_10__7_ & ~n50863;
  assign n50865 = n44095 & n50853;
  assign n50866 = n44097 & n50860;
  assign n50867 = n44059 & ~n50866;
  assign n50868 = ~n50857 & ~n50867;
  assign n50869 = n44369 & n50868;
  assign n50870 = n47261 & n50859;
  assign n50871 = ~n50864 & ~n50865;
  assign n50872 = ~n50869 & n50871;
  assign n50873 = ~n50870 & n50872;
  assign n50874 = ~n50187 & n50873;
  assign n50875 = ~n50858 & n50873;
  assign n8306 = ~n50874 & ~n50875;
  assign n50877 = P1_P1_INSTQUEUE_REG_10__6_ & ~n50863;
  assign n50878 = n50204 & n50868;
  assign n50879 = n50206 & n50853;
  assign n50880 = n50220 & n50859;
  assign n50881 = n50234 & n50858;
  assign n50882 = ~n50877 & ~n50878;
  assign n50883 = ~n50879 & n50882;
  assign n50884 = ~n50880 & n50883;
  assign n8311 = n50881 | ~n50884;
  assign n50886 = P1_P1_INSTQUEUE_REG_10__5_ & ~n50863;
  assign n50887 = n50251 & n50868;
  assign n50888 = n50253 & n50853;
  assign n50889 = n50264 & n50859;
  assign n50890 = n50276 & n50858;
  assign n50891 = ~n50886 & ~n50887;
  assign n50892 = ~n50888 & n50891;
  assign n50893 = ~n50889 & n50892;
  assign n8316 = n50890 | ~n50893;
  assign n50895 = P1_P1_INSTQUEUE_REG_10__4_ & ~n50863;
  assign n50896 = n50295 & n50868;
  assign n50897 = n50297 & n50853;
  assign n50898 = n50310 & n50859;
  assign n50899 = n50322 & n50858;
  assign n50900 = ~n50895 & ~n50896;
  assign n50901 = ~n50897 & n50900;
  assign n50902 = ~n50898 & n50901;
  assign n8321 = n50899 | ~n50902;
  assign n50904 = P1_P1_INSTQUEUE_REG_10__3_ & ~n50863;
  assign n50905 = n50339 & n50868;
  assign n50906 = n50341 & n50853;
  assign n50907 = n50353 & n50859;
  assign n50908 = n50363 & n50858;
  assign n50909 = ~n50904 & ~n50905;
  assign n50910 = ~n50906 & n50909;
  assign n50911 = ~n50907 & n50910;
  assign n8326 = n50908 | ~n50911;
  assign n50913 = P1_P1_INSTQUEUE_REG_10__2_ & ~n50863;
  assign n50914 = n50381 & n50868;
  assign n50915 = n50383 & n50853;
  assign n50916 = n50397 & n50859;
  assign n50917 = n50411 & n50858;
  assign n50918 = ~n50913 & ~n50914;
  assign n50919 = ~n50915 & n50918;
  assign n50920 = ~n50916 & n50919;
  assign n8331 = n50917 | ~n50920;
  assign n50922 = P1_P1_INSTQUEUE_REG_10__1_ & ~n50863;
  assign n50923 = n50426 & n50868;
  assign n50924 = n50428 & n50853;
  assign n50925 = n50437 & n50859;
  assign n50926 = n50449 & n50858;
  assign n50927 = ~n50922 & ~n50923;
  assign n50928 = ~n50924 & n50927;
  assign n50929 = ~n50925 & n50928;
  assign n8336 = n50926 | ~n50929;
  assign n50931 = P1_P1_INSTQUEUE_REG_10__0_ & ~n50863;
  assign n50932 = n50459 & n50868;
  assign n50933 = n50461 & n50853;
  assign n50934 = n50474 & n50859;
  assign n50935 = n50488 & n50858;
  assign n50936 = ~n50931 & ~n50932;
  assign n50937 = ~n50933 & n50936;
  assign n50938 = ~n50934 & n50937;
  assign n8341 = n50935 | ~n50938;
  assign n50940 = n44051 & n50762;
  assign n50941 = P1_P1_STATE2_REG_3_ & ~n50940;
  assign n50942 = n44042 & ~n50941;
  assign n50943 = n44061 & n50766;
  assign n50944 = ~n50940 & ~n50943;
  assign n50945 = n50590 & n50769;
  assign n50946 = n44064 & n44079;
  assign n50947 = ~n50945 & ~n50946;
  assign n50948 = n44059 & ~n50947;
  assign n50949 = n50944 & ~n50948;
  assign n50950 = n50942 & ~n50949;
  assign n50951 = P1_P1_INSTQUEUE_REG_9__7_ & ~n50950;
  assign n50952 = n44095 & n50940;
  assign n50953 = n44097 & n50947;
  assign n50954 = n44059 & ~n50953;
  assign n50955 = ~n50944 & ~n50954;
  assign n50956 = n44369 & n50955;
  assign n50957 = n47261 & n50946;
  assign n50958 = ~n50951 & ~n50952;
  assign n50959 = ~n50956 & n50958;
  assign n50960 = ~n50957 & n50959;
  assign n50961 = ~n50187 & n50960;
  assign n50962 = ~n50945 & n50960;
  assign n8346 = ~n50961 & ~n50962;
  assign n50964 = P1_P1_INSTQUEUE_REG_9__6_ & ~n50950;
  assign n50965 = n50204 & n50955;
  assign n50966 = n50206 & n50940;
  assign n50967 = n50220 & n50946;
  assign n50968 = n50234 & n50945;
  assign n50969 = ~n50964 & ~n50965;
  assign n50970 = ~n50966 & n50969;
  assign n50971 = ~n50967 & n50970;
  assign n8351 = n50968 | ~n50971;
  assign n50973 = P1_P1_INSTQUEUE_REG_9__5_ & ~n50950;
  assign n50974 = n50251 & n50955;
  assign n50975 = n50253 & n50940;
  assign n50976 = n50264 & n50946;
  assign n50977 = n50276 & n50945;
  assign n50978 = ~n50973 & ~n50974;
  assign n50979 = ~n50975 & n50978;
  assign n50980 = ~n50976 & n50979;
  assign n8356 = n50977 | ~n50980;
  assign n50982 = P1_P1_INSTQUEUE_REG_9__4_ & ~n50950;
  assign n50983 = n50295 & n50955;
  assign n50984 = n50297 & n50940;
  assign n50985 = n50310 & n50946;
  assign n50986 = n50322 & n50945;
  assign n50987 = ~n50982 & ~n50983;
  assign n50988 = ~n50984 & n50987;
  assign n50989 = ~n50985 & n50988;
  assign n8361 = n50986 | ~n50989;
  assign n50991 = P1_P1_INSTQUEUE_REG_9__3_ & ~n50950;
  assign n50992 = n50339 & n50955;
  assign n50993 = n50341 & n50940;
  assign n50994 = n50353 & n50946;
  assign n50995 = n50363 & n50945;
  assign n50996 = ~n50991 & ~n50992;
  assign n50997 = ~n50993 & n50996;
  assign n50998 = ~n50994 & n50997;
  assign n8366 = n50995 | ~n50998;
  assign n51000 = P1_P1_INSTQUEUE_REG_9__2_ & ~n50950;
  assign n51001 = n50381 & n50955;
  assign n51002 = n50383 & n50940;
  assign n51003 = n50397 & n50946;
  assign n51004 = n50411 & n50945;
  assign n51005 = ~n51000 & ~n51001;
  assign n51006 = ~n51002 & n51005;
  assign n51007 = ~n51003 & n51006;
  assign n8371 = n51004 | ~n51007;
  assign n51009 = P1_P1_INSTQUEUE_REG_9__1_ & ~n50950;
  assign n51010 = n50426 & n50955;
  assign n51011 = n50428 & n50940;
  assign n51012 = n50437 & n50946;
  assign n51013 = n50449 & n50945;
  assign n51014 = ~n51009 & ~n51010;
  assign n51015 = ~n51011 & n51014;
  assign n51016 = ~n51012 & n51015;
  assign n8376 = n51013 | ~n51016;
  assign n51018 = P1_P1_INSTQUEUE_REG_9__0_ & ~n50950;
  assign n51019 = n50459 & n50955;
  assign n51020 = n50461 & n50940;
  assign n51021 = n50474 & n50946;
  assign n51022 = n50488 & n50945;
  assign n51023 = ~n51018 & ~n51019;
  assign n51024 = ~n51020 & n51023;
  assign n51025 = ~n51021 & n51024;
  assign n8381 = n51022 | ~n51025;
  assign n51027 = n50673 & n50852;
  assign n51028 = P1_P1_STATE2_REG_3_ & ~n51027;
  assign n51029 = n44042 & ~n51028;
  assign n51030 = n50677 & n50769;
  assign n51031 = n44079 & n50679;
  assign n51032 = ~n51030 & ~n51031;
  assign n51033 = n44059 & ~n51032;
  assign n51034 = n44053 & n50766;
  assign n51035 = ~n51033 & ~n51034;
  assign n51036 = n51029 & ~n51035;
  assign n51037 = P1_P1_INSTQUEUE_REG_8__7_ & ~n51036;
  assign n51038 = n44095 & n51027;
  assign n51039 = n44097 & n51032;
  assign n51040 = n44059 & ~n51039;
  assign n51041 = n51034 & ~n51040;
  assign n51042 = n44369 & n51041;
  assign n51043 = n47261 & n51031;
  assign n51044 = ~n51037 & ~n51038;
  assign n51045 = ~n51042 & n51044;
  assign n51046 = ~n51043 & n51045;
  assign n51047 = ~n50187 & n51046;
  assign n51048 = ~n51030 & n51046;
  assign n8386 = ~n51047 & ~n51048;
  assign n51050 = P1_P1_INSTQUEUE_REG_8__6_ & ~n51036;
  assign n51051 = n50204 & n51041;
  assign n51052 = n50206 & n51027;
  assign n51053 = n50220 & n51031;
  assign n51054 = n50234 & n51030;
  assign n51055 = ~n51050 & ~n51051;
  assign n51056 = ~n51052 & n51055;
  assign n51057 = ~n51053 & n51056;
  assign n8391 = n51054 | ~n51057;
  assign n51059 = P1_P1_INSTQUEUE_REG_8__5_ & ~n51036;
  assign n51060 = n50251 & n51041;
  assign n51061 = n50253 & n51027;
  assign n51062 = n50264 & n51031;
  assign n51063 = n50276 & n51030;
  assign n51064 = ~n51059 & ~n51060;
  assign n51065 = ~n51061 & n51064;
  assign n51066 = ~n51062 & n51065;
  assign n8396 = n51063 | ~n51066;
  assign n51068 = P1_P1_INSTQUEUE_REG_8__4_ & ~n51036;
  assign n51069 = n50295 & n51041;
  assign n51070 = n50297 & n51027;
  assign n51071 = n50310 & n51031;
  assign n51072 = n50322 & n51030;
  assign n51073 = ~n51068 & ~n51069;
  assign n51074 = ~n51070 & n51073;
  assign n51075 = ~n51071 & n51074;
  assign n8401 = n51072 | ~n51075;
  assign n51077 = P1_P1_INSTQUEUE_REG_8__3_ & ~n51036;
  assign n51078 = n50339 & n51041;
  assign n51079 = n50341 & n51027;
  assign n51080 = n50353 & n51031;
  assign n51081 = n50363 & n51030;
  assign n51082 = ~n51077 & ~n51078;
  assign n51083 = ~n51079 & n51082;
  assign n51084 = ~n51080 & n51083;
  assign n8406 = n51081 | ~n51084;
  assign n51086 = P1_P1_INSTQUEUE_REG_8__2_ & ~n51036;
  assign n51087 = n50381 & n51041;
  assign n51088 = n50383 & n51027;
  assign n51089 = n50397 & n51031;
  assign n51090 = n50411 & n51030;
  assign n51091 = ~n51086 & ~n51087;
  assign n51092 = ~n51088 & n51091;
  assign n51093 = ~n51089 & n51092;
  assign n8411 = n51090 | ~n51093;
  assign n51095 = P1_P1_INSTQUEUE_REG_8__1_ & ~n51036;
  assign n51096 = n50426 & n51041;
  assign n51097 = n50428 & n51027;
  assign n51098 = n50437 & n51031;
  assign n51099 = n50449 & n51030;
  assign n51100 = ~n51095 & ~n51096;
  assign n51101 = ~n51097 & n51100;
  assign n51102 = ~n51098 & n51101;
  assign n8416 = n51099 | ~n51102;
  assign n51104 = P1_P1_INSTQUEUE_REG_8__0_ & ~n51036;
  assign n51105 = n50459 & n51041;
  assign n51106 = n50461 & n51027;
  assign n51107 = n50474 & n51031;
  assign n51108 = n50488 & n51030;
  assign n51109 = ~n51104 & ~n51105;
  assign n51110 = ~n51106 & n51109;
  assign n51111 = ~n51107 & n51110;
  assign n8421 = n51108 | ~n51111;
  assign n51113 = P1_P1_STATE2_REG_3_ & ~n44047;
  assign n51114 = n44042 & ~n51113;
  assign n51115 = ~n44047 & ~n44075;
  assign n51116 = ~n44073 & n44084;
  assign n51117 = n44066 & n51116;
  assign n51118 = ~n44083 & ~n51117;
  assign n51119 = n44059 & ~n51118;
  assign n51120 = n51115 & ~n51119;
  assign n51121 = n51114 & ~n51120;
  assign n51122 = P1_P1_INSTQUEUE_REG_7__7_ & ~n51121;
  assign n51123 = n44047 & n44095;
  assign n51124 = n44097 & n51118;
  assign n51125 = n44059 & ~n51124;
  assign n51126 = ~n51115 & ~n51125;
  assign n51127 = n44369 & n51126;
  assign n51128 = n44083 & n47261;
  assign n51129 = ~n51122 & ~n51123;
  assign n51130 = ~n51127 & n51129;
  assign n51131 = ~n51128 & n51130;
  assign n51132 = ~n50187 & n51131;
  assign n51133 = ~n51117 & n51131;
  assign n8426 = ~n51132 & ~n51133;
  assign n51135 = P1_P1_INSTQUEUE_REG_7__6_ & ~n51121;
  assign n51136 = n50204 & n51126;
  assign n51137 = n44047 & n50206;
  assign n51138 = n44083 & n50220;
  assign n51139 = n50234 & n51117;
  assign n51140 = ~n51135 & ~n51136;
  assign n51141 = ~n51137 & n51140;
  assign n51142 = ~n51138 & n51141;
  assign n8431 = n51139 | ~n51142;
  assign n51144 = P1_P1_INSTQUEUE_REG_7__5_ & ~n51121;
  assign n51145 = n50251 & n51126;
  assign n51146 = n44047 & n50253;
  assign n51147 = n44083 & n50264;
  assign n51148 = n50276 & n51117;
  assign n51149 = ~n51144 & ~n51145;
  assign n51150 = ~n51146 & n51149;
  assign n51151 = ~n51147 & n51150;
  assign n8436 = n51148 | ~n51151;
  assign n51153 = P1_P1_INSTQUEUE_REG_7__4_ & ~n51121;
  assign n51154 = n50295 & n51126;
  assign n51155 = n44047 & n50297;
  assign n51156 = n44083 & n50310;
  assign n51157 = n50322 & n51117;
  assign n51158 = ~n51153 & ~n51154;
  assign n51159 = ~n51155 & n51158;
  assign n51160 = ~n51156 & n51159;
  assign n8441 = n51157 | ~n51160;
  assign n51162 = P1_P1_INSTQUEUE_REG_7__3_ & ~n51121;
  assign n51163 = n50339 & n51126;
  assign n51164 = n44047 & n50341;
  assign n51165 = n44083 & n50353;
  assign n51166 = n50363 & n51117;
  assign n51167 = ~n51162 & ~n51163;
  assign n51168 = ~n51164 & n51167;
  assign n51169 = ~n51165 & n51168;
  assign n8446 = n51166 | ~n51169;
  assign n51171 = P1_P1_INSTQUEUE_REG_7__2_ & ~n51121;
  assign n51172 = n50381 & n51126;
  assign n51173 = n44047 & n50383;
  assign n51174 = n44083 & n50397;
  assign n51175 = n50411 & n51117;
  assign n51176 = ~n51171 & ~n51172;
  assign n51177 = ~n51173 & n51176;
  assign n51178 = ~n51174 & n51177;
  assign n8451 = n51175 | ~n51178;
  assign n51180 = P1_P1_INSTQUEUE_REG_7__1_ & ~n51121;
  assign n51181 = n50426 & n51126;
  assign n51182 = n44047 & n50428;
  assign n51183 = n44083 & n50437;
  assign n51184 = n50449 & n51117;
  assign n51185 = ~n51180 & ~n51181;
  assign n51186 = ~n51182 & n51185;
  assign n51187 = ~n51183 & n51186;
  assign n8456 = n51184 | ~n51187;
  assign n51189 = P1_P1_INSTQUEUE_REG_7__0_ & ~n51121;
  assign n51190 = n50459 & n51126;
  assign n51191 = n44047 & n50461;
  assign n51192 = n44083 & n50474;
  assign n51193 = n50488 & n51117;
  assign n51194 = ~n51189 & ~n51190;
  assign n51195 = ~n51191 & n51194;
  assign n51196 = ~n51192 & n51195;
  assign n8461 = n51193 | ~n51196;
  assign n51198 = ~P1_P1_INSTQUEUEWR_ADDR_REG_3_ & P1_P1_INSTQUEUEWR_ADDR_REG_1_;
  assign n51199 = n50495 & n51198;
  assign n51200 = P1_P1_STATE2_REG_3_ & ~n51199;
  assign n51201 = n44042 & ~n51200;
  assign n51202 = n44060 & n44074;
  assign n51203 = ~n51199 & ~n51202;
  assign n51204 = n50501 & n51116;
  assign n51205 = n44063 & n44082;
  assign n51206 = ~n51204 & ~n51205;
  assign n51207 = n44059 & ~n51206;
  assign n51208 = n51203 & ~n51207;
  assign n51209 = n51201 & ~n51208;
  assign n51210 = P1_P1_INSTQUEUE_REG_6__7_ & ~n51209;
  assign n51211 = n44095 & n51199;
  assign n51212 = n44097 & n51206;
  assign n51213 = n44059 & ~n51212;
  assign n51214 = ~n51203 & ~n51213;
  assign n51215 = n44369 & n51214;
  assign n51216 = n47261 & n51205;
  assign n51217 = ~n51210 & ~n51211;
  assign n51218 = ~n51215 & n51217;
  assign n51219 = ~n51216 & n51218;
  assign n51220 = ~n50187 & n51219;
  assign n51221 = ~n51204 & n51219;
  assign n8466 = ~n51220 & ~n51221;
  assign n51223 = P1_P1_INSTQUEUE_REG_6__6_ & ~n51209;
  assign n51224 = n50204 & n51214;
  assign n51225 = n50206 & n51199;
  assign n51226 = n50220 & n51205;
  assign n51227 = n50234 & n51204;
  assign n51228 = ~n51223 & ~n51224;
  assign n51229 = ~n51225 & n51228;
  assign n51230 = ~n51226 & n51229;
  assign n8471 = n51227 | ~n51230;
  assign n51232 = P1_P1_INSTQUEUE_REG_6__5_ & ~n51209;
  assign n51233 = n50251 & n51214;
  assign n51234 = n50253 & n51199;
  assign n51235 = n50264 & n51205;
  assign n51236 = n50276 & n51204;
  assign n51237 = ~n51232 & ~n51233;
  assign n51238 = ~n51234 & n51237;
  assign n51239 = ~n51235 & n51238;
  assign n8476 = n51236 | ~n51239;
  assign n51241 = P1_P1_INSTQUEUE_REG_6__4_ & ~n51209;
  assign n51242 = n50295 & n51214;
  assign n51243 = n50297 & n51199;
  assign n51244 = n50310 & n51205;
  assign n51245 = n50322 & n51204;
  assign n51246 = ~n51241 & ~n51242;
  assign n51247 = ~n51243 & n51246;
  assign n51248 = ~n51244 & n51247;
  assign n8481 = n51245 | ~n51248;
  assign n51250 = P1_P1_INSTQUEUE_REG_6__3_ & ~n51209;
  assign n51251 = n50339 & n51214;
  assign n51252 = n50341 & n51199;
  assign n51253 = n50353 & n51205;
  assign n51254 = n50363 & n51204;
  assign n51255 = ~n51250 & ~n51251;
  assign n51256 = ~n51252 & n51255;
  assign n51257 = ~n51253 & n51256;
  assign n8486 = n51254 | ~n51257;
  assign n51259 = P1_P1_INSTQUEUE_REG_6__2_ & ~n51209;
  assign n51260 = n50381 & n51214;
  assign n51261 = n50383 & n51199;
  assign n51262 = n50397 & n51205;
  assign n51263 = n50411 & n51204;
  assign n51264 = ~n51259 & ~n51260;
  assign n51265 = ~n51261 & n51264;
  assign n51266 = ~n51262 & n51265;
  assign n8491 = n51263 | ~n51266;
  assign n51268 = P1_P1_INSTQUEUE_REG_6__1_ & ~n51209;
  assign n51269 = n50426 & n51214;
  assign n51270 = n50428 & n51199;
  assign n51271 = n50437 & n51205;
  assign n51272 = n50449 & n51204;
  assign n51273 = ~n51268 & ~n51269;
  assign n51274 = ~n51270 & n51273;
  assign n51275 = ~n51271 & n51274;
  assign n8496 = n51272 | ~n51275;
  assign n51277 = P1_P1_INSTQUEUE_REG_6__0_ & ~n51209;
  assign n51278 = n50459 & n51214;
  assign n51279 = n50461 & n51199;
  assign n51280 = n50474 & n51205;
  assign n51281 = n50488 & n51204;
  assign n51282 = ~n51277 & ~n51278;
  assign n51283 = ~n51279 & n51282;
  assign n51284 = ~n51280 & n51283;
  assign n8501 = n51281 | ~n51284;
  assign n51286 = ~P1_P1_INSTQUEUEWR_ADDR_REG_3_ & P1_P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n51287 = n44051 & n51286;
  assign n51288 = P1_P1_STATE2_REG_3_ & ~n51287;
  assign n51289 = n44042 & ~n51288;
  assign n51290 = n44061 & n44074;
  assign n51291 = ~n51287 & ~n51290;
  assign n51292 = n50590 & n51116;
  assign n51293 = n44064 & n44082;
  assign n51294 = ~n51292 & ~n51293;
  assign n51295 = n44059 & ~n51294;
  assign n51296 = n51291 & ~n51295;
  assign n51297 = n51289 & ~n51296;
  assign n51298 = P1_P1_INSTQUEUE_REG_5__7_ & ~n51297;
  assign n51299 = n44095 & n51287;
  assign n51300 = n44097 & n51294;
  assign n51301 = n44059 & ~n51300;
  assign n51302 = ~n51291 & ~n51301;
  assign n51303 = n44369 & n51302;
  assign n51304 = n47261 & n51293;
  assign n51305 = ~n51298 & ~n51299;
  assign n51306 = ~n51303 & n51305;
  assign n51307 = ~n51304 & n51306;
  assign n51308 = ~n50187 & n51307;
  assign n51309 = ~n51292 & n51307;
  assign n8506 = ~n51308 & ~n51309;
  assign n51311 = P1_P1_INSTQUEUE_REG_5__6_ & ~n51297;
  assign n51312 = n50204 & n51302;
  assign n51313 = n50206 & n51287;
  assign n51314 = n50220 & n51293;
  assign n51315 = n50234 & n51292;
  assign n51316 = ~n51311 & ~n51312;
  assign n51317 = ~n51313 & n51316;
  assign n51318 = ~n51314 & n51317;
  assign n8511 = n51315 | ~n51318;
  assign n51320 = P1_P1_INSTQUEUE_REG_5__5_ & ~n51297;
  assign n51321 = n50251 & n51302;
  assign n51322 = n50253 & n51287;
  assign n51323 = n50264 & n51293;
  assign n51324 = n50276 & n51292;
  assign n51325 = ~n51320 & ~n51321;
  assign n51326 = ~n51322 & n51325;
  assign n51327 = ~n51323 & n51326;
  assign n8516 = n51324 | ~n51327;
  assign n51329 = P1_P1_INSTQUEUE_REG_5__4_ & ~n51297;
  assign n51330 = n50295 & n51302;
  assign n51331 = n50297 & n51287;
  assign n51332 = n50310 & n51293;
  assign n51333 = n50322 & n51292;
  assign n51334 = ~n51329 & ~n51330;
  assign n51335 = ~n51331 & n51334;
  assign n51336 = ~n51332 & n51335;
  assign n8521 = n51333 | ~n51336;
  assign n51338 = P1_P1_INSTQUEUE_REG_5__3_ & ~n51297;
  assign n51339 = n50339 & n51302;
  assign n51340 = n50341 & n51287;
  assign n51341 = n50353 & n51293;
  assign n51342 = n50363 & n51292;
  assign n51343 = ~n51338 & ~n51339;
  assign n51344 = ~n51340 & n51343;
  assign n51345 = ~n51341 & n51344;
  assign n8526 = n51342 | ~n51345;
  assign n51347 = P1_P1_INSTQUEUE_REG_5__2_ & ~n51297;
  assign n51348 = n50381 & n51302;
  assign n51349 = n50383 & n51287;
  assign n51350 = n50397 & n51293;
  assign n51351 = n50411 & n51292;
  assign n51352 = ~n51347 & ~n51348;
  assign n51353 = ~n51349 & n51352;
  assign n51354 = ~n51350 & n51353;
  assign n8531 = n51351 | ~n51354;
  assign n51356 = P1_P1_INSTQUEUE_REG_5__1_ & ~n51297;
  assign n51357 = n50426 & n51302;
  assign n51358 = n50428 & n51287;
  assign n51359 = n50437 & n51293;
  assign n51360 = n50449 & n51292;
  assign n51361 = ~n51356 & ~n51357;
  assign n51362 = ~n51358 & n51361;
  assign n51363 = ~n51359 & n51362;
  assign n8536 = n51360 | ~n51363;
  assign n51365 = P1_P1_INSTQUEUE_REG_5__0_ & ~n51297;
  assign n51366 = n50459 & n51302;
  assign n51367 = n50461 & n51287;
  assign n51368 = n50474 & n51293;
  assign n51369 = n50488 & n51292;
  assign n51370 = ~n51365 & ~n51366;
  assign n51371 = ~n51367 & n51370;
  assign n51372 = ~n51368 & n51371;
  assign n8541 = n51369 | ~n51372;
  assign n51374 = ~P1_P1_INSTQUEUEWR_ADDR_REG_3_ & ~P1_P1_INSTQUEUEWR_ADDR_REG_1_;
  assign n51375 = n50495 & n51374;
  assign n51376 = P1_P1_STATE2_REG_3_ & ~n51375;
  assign n51377 = n44042 & ~n51376;
  assign n51378 = n50677 & n51116;
  assign n51379 = n44082 & n50679;
  assign n51380 = ~n51378 & ~n51379;
  assign n51381 = n44059 & ~n51380;
  assign n51382 = n44053 & n44074;
  assign n51383 = ~n51381 & ~n51382;
  assign n51384 = n51377 & ~n51383;
  assign n51385 = P1_P1_INSTQUEUE_REG_4__7_ & ~n51384;
  assign n51386 = n44095 & n51375;
  assign n51387 = n44059 & ~n44097;
  assign n51388 = n51382 & ~n51387;
  assign n51389 = n44369 & n51388;
  assign n51390 = n47261 & n51379;
  assign n51391 = ~n51385 & ~n51386;
  assign n51392 = ~n51389 & n51391;
  assign n51393 = ~n51390 & n51392;
  assign n51394 = ~n50187 & n51393;
  assign n51395 = ~n51378 & n51393;
  assign n8546 = ~n51394 & ~n51395;
  assign n51397 = P1_P1_INSTQUEUE_REG_4__6_ & ~n51384;
  assign n51398 = n50204 & n51388;
  assign n51399 = n50206 & n51375;
  assign n51400 = n50220 & n51379;
  assign n51401 = n50234 & n51378;
  assign n51402 = ~n51397 & ~n51398;
  assign n51403 = ~n51399 & n51402;
  assign n51404 = ~n51400 & n51403;
  assign n8551 = n51401 | ~n51404;
  assign n51406 = P1_P1_INSTQUEUE_REG_4__5_ & ~n51384;
  assign n51407 = n50251 & n51388;
  assign n51408 = n50253 & n51375;
  assign n51409 = n50264 & n51379;
  assign n51410 = n50276 & n51378;
  assign n51411 = ~n51406 & ~n51407;
  assign n51412 = ~n51408 & n51411;
  assign n51413 = ~n51409 & n51412;
  assign n8556 = n51410 | ~n51413;
  assign n51415 = P1_P1_INSTQUEUE_REG_4__4_ & ~n51384;
  assign n51416 = n50295 & n51388;
  assign n51417 = n50297 & n51375;
  assign n51418 = n50310 & n51379;
  assign n51419 = n50322 & n51378;
  assign n51420 = ~n51415 & ~n51416;
  assign n51421 = ~n51417 & n51420;
  assign n51422 = ~n51418 & n51421;
  assign n8561 = n51419 | ~n51422;
  assign n51424 = P1_P1_INSTQUEUE_REG_4__3_ & ~n51384;
  assign n51425 = n50339 & n51388;
  assign n51426 = n50341 & n51375;
  assign n51427 = n50353 & n51379;
  assign n51428 = n50363 & n51378;
  assign n51429 = ~n51424 & ~n51425;
  assign n51430 = ~n51426 & n51429;
  assign n51431 = ~n51427 & n51430;
  assign n8566 = n51428 | ~n51431;
  assign n51433 = P1_P1_INSTQUEUE_REG_4__2_ & ~n51384;
  assign n51434 = n50381 & n51388;
  assign n51435 = n50383 & n51375;
  assign n51436 = n50397 & n51379;
  assign n51437 = n50411 & n51378;
  assign n51438 = ~n51433 & ~n51434;
  assign n51439 = ~n51435 & n51438;
  assign n51440 = ~n51436 & n51439;
  assign n8571 = n51437 | ~n51440;
  assign n51442 = P1_P1_INSTQUEUE_REG_4__1_ & ~n51384;
  assign n51443 = n50426 & n51388;
  assign n51444 = n50428 & n51375;
  assign n51445 = n50437 & n51379;
  assign n51446 = n50449 & n51378;
  assign n51447 = ~n51442 & ~n51443;
  assign n51448 = ~n51444 & n51447;
  assign n51449 = ~n51445 & n51448;
  assign n8576 = n51446 | ~n51449;
  assign n51451 = P1_P1_INSTQUEUE_REG_4__0_ & ~n51384;
  assign n51452 = n50459 & n51388;
  assign n51453 = n50461 & n51375;
  assign n51454 = n50474 & n51379;
  assign n51455 = n50488 & n51378;
  assign n51456 = ~n51451 & ~n51452;
  assign n51457 = ~n51453 & n51456;
  assign n51458 = ~n51454 & n51457;
  assign n8581 = n51455 | ~n51458;
  assign n51460 = ~P1_P1_INSTQUEUEWR_ADDR_REG_3_ & ~P1_P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n51461 = n44035 & n51460;
  assign n51462 = P1_P1_STATE2_REG_3_ & ~n51461;
  assign n51463 = n44042 & ~n51462;
  assign n51464 = n44046 & n44049;
  assign n51465 = n44054 & n51464;
  assign n51466 = ~n51461 & ~n51465;
  assign n51467 = n44073 & n44084;
  assign n51468 = n44066 & n51467;
  assign n51469 = n44069 & n44078;
  assign n51470 = n44070 & n51469;
  assign n51471 = ~n51468 & ~n51470;
  assign n51472 = n44059 & ~n51471;
  assign n51473 = n51466 & ~n51472;
  assign n51474 = n51463 & ~n51473;
  assign n51475 = P1_P1_INSTQUEUE_REG_3__7_ & ~n51474;
  assign n51476 = n44095 & n51461;
  assign n51477 = ~n51387 & ~n51466;
  assign n51478 = n44369 & n51477;
  assign n51479 = n47261 & n51470;
  assign n51480 = ~n51475 & ~n51476;
  assign n51481 = ~n51478 & n51480;
  assign n51482 = ~n51479 & n51481;
  assign n51483 = ~n50187 & n51482;
  assign n51484 = ~n51468 & n51482;
  assign n8586 = ~n51483 & ~n51484;
  assign n51486 = P1_P1_INSTQUEUE_REG_3__6_ & ~n51474;
  assign n51487 = n50204 & n51477;
  assign n51488 = n50206 & n51461;
  assign n51489 = n50220 & n51470;
  assign n51490 = n50234 & n51468;
  assign n51491 = ~n51486 & ~n51487;
  assign n51492 = ~n51488 & n51491;
  assign n51493 = ~n51489 & n51492;
  assign n8591 = n51490 | ~n51493;
  assign n51495 = P1_P1_INSTQUEUE_REG_3__5_ & ~n51474;
  assign n51496 = n50251 & n51477;
  assign n51497 = n50253 & n51461;
  assign n51498 = n50264 & n51470;
  assign n51499 = n50276 & n51468;
  assign n51500 = ~n51495 & ~n51496;
  assign n51501 = ~n51497 & n51500;
  assign n51502 = ~n51498 & n51501;
  assign n8596 = n51499 | ~n51502;
  assign n51504 = P1_P1_INSTQUEUE_REG_3__4_ & ~n51474;
  assign n51505 = n50295 & n51477;
  assign n51506 = n50297 & n51461;
  assign n51507 = n50310 & n51470;
  assign n51508 = n50322 & n51468;
  assign n51509 = ~n51504 & ~n51505;
  assign n51510 = ~n51506 & n51509;
  assign n51511 = ~n51507 & n51510;
  assign n8601 = n51508 | ~n51511;
  assign n51513 = P1_P1_INSTQUEUE_REG_3__3_ & ~n51474;
  assign n51514 = n50339 & n51477;
  assign n51515 = n50341 & n51461;
  assign n51516 = n50353 & n51470;
  assign n51517 = n50363 & n51468;
  assign n51518 = ~n51513 & ~n51514;
  assign n51519 = ~n51515 & n51518;
  assign n51520 = ~n51516 & n51519;
  assign n8606 = n51517 | ~n51520;
  assign n51522 = P1_P1_INSTQUEUE_REG_3__2_ & ~n51474;
  assign n51523 = n50381 & n51477;
  assign n51524 = n50383 & n51461;
  assign n51525 = n50397 & n51470;
  assign n51526 = n50411 & n51468;
  assign n51527 = ~n51522 & ~n51523;
  assign n51528 = ~n51524 & n51527;
  assign n51529 = ~n51525 & n51528;
  assign n8611 = n51526 | ~n51529;
  assign n51531 = P1_P1_INSTQUEUE_REG_3__1_ & ~n51474;
  assign n51532 = n50426 & n51477;
  assign n51533 = n50428 & n51461;
  assign n51534 = n50437 & n51470;
  assign n51535 = n50449 & n51468;
  assign n51536 = ~n51531 & ~n51532;
  assign n51537 = ~n51533 & n51536;
  assign n51538 = ~n51534 & n51537;
  assign n8616 = n51535 | ~n51538;
  assign n51540 = P1_P1_INSTQUEUE_REG_3__0_ & ~n51474;
  assign n51541 = n50459 & n51477;
  assign n51542 = n50461 & n51461;
  assign n51543 = n50474 & n51470;
  assign n51544 = n50488 & n51468;
  assign n51545 = ~n51540 & ~n51541;
  assign n51546 = ~n51542 & n51545;
  assign n51547 = ~n51543 & n51546;
  assign n8621 = n51544 | ~n51547;
  assign n51549 = n50852 & n51198;
  assign n51550 = P1_P1_STATE2_REG_3_ & ~n51549;
  assign n51551 = n44042 & ~n51550;
  assign n51552 = n44060 & n51464;
  assign n51553 = ~n51549 & ~n51552;
  assign n51554 = n50501 & n51467;
  assign n51555 = n44063 & n51469;
  assign n51556 = ~n51554 & ~n51555;
  assign n51557 = n44059 & ~n51556;
  assign n51558 = n51553 & ~n51557;
  assign n51559 = n51551 & ~n51558;
  assign n51560 = P1_P1_INSTQUEUE_REG_2__7_ & ~n51559;
  assign n51561 = n44095 & n51549;
  assign n51562 = ~n51387 & ~n51553;
  assign n51563 = n44369 & n51562;
  assign n51564 = n47261 & n51555;
  assign n51565 = ~n51560 & ~n51561;
  assign n51566 = ~n51563 & n51565;
  assign n51567 = ~n51564 & n51566;
  assign n51568 = ~n50187 & n51567;
  assign n51569 = ~n51554 & n51567;
  assign n8626 = ~n51568 & ~n51569;
  assign n51571 = P1_P1_INSTQUEUE_REG_2__6_ & ~n51559;
  assign n51572 = n50204 & n51562;
  assign n51573 = n50206 & n51549;
  assign n51574 = n50220 & n51555;
  assign n51575 = n50234 & n51554;
  assign n51576 = ~n51571 & ~n51572;
  assign n51577 = ~n51573 & n51576;
  assign n51578 = ~n51574 & n51577;
  assign n8631 = n51575 | ~n51578;
  assign n51580 = P1_P1_INSTQUEUE_REG_2__5_ & ~n51559;
  assign n51581 = n50251 & n51562;
  assign n51582 = n50253 & n51549;
  assign n51583 = n50264 & n51555;
  assign n51584 = n50276 & n51554;
  assign n51585 = ~n51580 & ~n51581;
  assign n51586 = ~n51582 & n51585;
  assign n51587 = ~n51583 & n51586;
  assign n8636 = n51584 | ~n51587;
  assign n51589 = P1_P1_INSTQUEUE_REG_2__4_ & ~n51559;
  assign n51590 = n50295 & n51562;
  assign n51591 = n50297 & n51549;
  assign n51592 = n50310 & n51555;
  assign n51593 = n50322 & n51554;
  assign n51594 = ~n51589 & ~n51590;
  assign n51595 = ~n51591 & n51594;
  assign n51596 = ~n51592 & n51595;
  assign n8641 = n51593 | ~n51596;
  assign n51598 = P1_P1_INSTQUEUE_REG_2__3_ & ~n51559;
  assign n51599 = n50339 & n51562;
  assign n51600 = n50341 & n51549;
  assign n51601 = n50353 & n51555;
  assign n51602 = n50363 & n51554;
  assign n51603 = ~n51598 & ~n51599;
  assign n51604 = ~n51600 & n51603;
  assign n51605 = ~n51601 & n51604;
  assign n8646 = n51602 | ~n51605;
  assign n51607 = P1_P1_INSTQUEUE_REG_2__2_ & ~n51559;
  assign n51608 = n50381 & n51562;
  assign n51609 = n50383 & n51549;
  assign n51610 = n50397 & n51555;
  assign n51611 = n50411 & n51554;
  assign n51612 = ~n51607 & ~n51608;
  assign n51613 = ~n51609 & n51612;
  assign n51614 = ~n51610 & n51613;
  assign n8651 = n51611 | ~n51614;
  assign n51616 = P1_P1_INSTQUEUE_REG_2__1_ & ~n51559;
  assign n51617 = n50426 & n51562;
  assign n51618 = n50428 & n51549;
  assign n51619 = n50437 & n51555;
  assign n51620 = n50449 & n51554;
  assign n51621 = ~n51616 & ~n51617;
  assign n51622 = ~n51618 & n51621;
  assign n51623 = ~n51619 & n51622;
  assign n8656 = n51620 | ~n51623;
  assign n51625 = P1_P1_INSTQUEUE_REG_2__0_ & ~n51559;
  assign n51626 = n50459 & n51562;
  assign n51627 = n50461 & n51549;
  assign n51628 = n50474 & n51555;
  assign n51629 = n50488 & n51554;
  assign n51630 = ~n51625 & ~n51626;
  assign n51631 = ~n51627 & n51630;
  assign n51632 = ~n51628 & n51631;
  assign n8661 = n51629 | ~n51632;
  assign n51634 = n44051 & n51460;
  assign n51635 = P1_P1_STATE2_REG_3_ & ~n51634;
  assign n51636 = n44042 & ~n51635;
  assign n51637 = n44061 & n51464;
  assign n51638 = ~n51634 & ~n51637;
  assign n51639 = n50590 & n51467;
  assign n51640 = n44064 & n51469;
  assign n51641 = ~n51639 & ~n51640;
  assign n51642 = n44059 & ~n51641;
  assign n51643 = n51638 & ~n51642;
  assign n51644 = n51636 & ~n51643;
  assign n51645 = P1_P1_INSTQUEUE_REG_1__7_ & ~n51644;
  assign n51646 = n44095 & n51634;
  assign n51647 = ~n51387 & ~n51638;
  assign n51648 = n44369 & n51647;
  assign n51649 = n47261 & n51640;
  assign n51650 = ~n51645 & ~n51646;
  assign n51651 = ~n51648 & n51650;
  assign n51652 = ~n51649 & n51651;
  assign n51653 = ~n50187 & n51652;
  assign n51654 = ~n51639 & n51652;
  assign n8666 = ~n51653 & ~n51654;
  assign n51656 = P1_P1_INSTQUEUE_REG_1__6_ & ~n51644;
  assign n51657 = n50204 & n51647;
  assign n51658 = n50206 & n51634;
  assign n51659 = n50220 & n51640;
  assign n51660 = n50234 & n51639;
  assign n51661 = ~n51656 & ~n51657;
  assign n51662 = ~n51658 & n51661;
  assign n51663 = ~n51659 & n51662;
  assign n8671 = n51660 | ~n51663;
  assign n51665 = P1_P1_INSTQUEUE_REG_1__5_ & ~n51644;
  assign n51666 = n50251 & n51647;
  assign n51667 = n50253 & n51634;
  assign n51668 = n50264 & n51640;
  assign n51669 = n50276 & n51639;
  assign n51670 = ~n51665 & ~n51666;
  assign n51671 = ~n51667 & n51670;
  assign n51672 = ~n51668 & n51671;
  assign n8676 = n51669 | ~n51672;
  assign n51674 = P1_P1_INSTQUEUE_REG_1__4_ & ~n51644;
  assign n51675 = n50295 & n51647;
  assign n51676 = n50297 & n51634;
  assign n51677 = n50310 & n51640;
  assign n51678 = n50322 & n51639;
  assign n51679 = ~n51674 & ~n51675;
  assign n51680 = ~n51676 & n51679;
  assign n51681 = ~n51677 & n51680;
  assign n8681 = n51678 | ~n51681;
  assign n51683 = P1_P1_INSTQUEUE_REG_1__3_ & ~n51644;
  assign n51684 = n50339 & n51647;
  assign n51685 = n50341 & n51634;
  assign n51686 = n50353 & n51640;
  assign n51687 = n50363 & n51639;
  assign n51688 = ~n51683 & ~n51684;
  assign n51689 = ~n51685 & n51688;
  assign n51690 = ~n51686 & n51689;
  assign n8686 = n51687 | ~n51690;
  assign n51692 = P1_P1_INSTQUEUE_REG_1__2_ & ~n51644;
  assign n51693 = n50381 & n51647;
  assign n51694 = n50383 & n51634;
  assign n51695 = n50397 & n51640;
  assign n51696 = n50411 & n51639;
  assign n51697 = ~n51692 & ~n51693;
  assign n51698 = ~n51694 & n51697;
  assign n51699 = ~n51695 & n51698;
  assign n8691 = n51696 | ~n51699;
  assign n51701 = P1_P1_INSTQUEUE_REG_1__1_ & ~n51644;
  assign n51702 = n50426 & n51647;
  assign n51703 = n50428 & n51634;
  assign n51704 = n50437 & n51640;
  assign n51705 = n50449 & n51639;
  assign n51706 = ~n51701 & ~n51702;
  assign n51707 = ~n51703 & n51706;
  assign n51708 = ~n51704 & n51707;
  assign n8696 = n51705 | ~n51708;
  assign n51710 = P1_P1_INSTQUEUE_REG_1__0_ & ~n51644;
  assign n51711 = n50459 & n51647;
  assign n51712 = n50461 & n51634;
  assign n51713 = n50474 & n51640;
  assign n51714 = n50488 & n51639;
  assign n51715 = ~n51710 & ~n51711;
  assign n51716 = ~n51712 & n51715;
  assign n51717 = ~n51713 & n51716;
  assign n8701 = n51714 | ~n51717;
  assign n51719 = n50852 & n51374;
  assign n51720 = P1_P1_STATE2_REG_3_ & ~n51719;
  assign n51721 = n44042 & ~n51720;
  assign n51722 = n50677 & n51467;
  assign n51723 = n50679 & n51469;
  assign n51724 = ~n51722 & ~n51723;
  assign n51725 = n44059 & ~n51724;
  assign n51726 = n44053 & n51464;
  assign n51727 = ~n51725 & ~n51726;
  assign n51728 = n51721 & ~n51727;
  assign n51729 = P1_P1_INSTQUEUE_REG_0__7_ & ~n51728;
  assign n51730 = n44095 & n51719;
  assign n51731 = ~n51387 & n51726;
  assign n51732 = n44369 & n51731;
  assign n51733 = n47261 & n51723;
  assign n51734 = ~n51729 & ~n51730;
  assign n51735 = ~n51732 & n51734;
  assign n51736 = ~n51733 & n51735;
  assign n51737 = ~n50187 & n51736;
  assign n51738 = ~n51722 & n51736;
  assign n8706 = ~n51737 & ~n51738;
  assign n51740 = P1_P1_INSTQUEUE_REG_0__6_ & ~n51728;
  assign n51741 = n50204 & n51731;
  assign n51742 = n50206 & n51719;
  assign n51743 = n50220 & n51723;
  assign n51744 = n50234 & n51722;
  assign n51745 = ~n51740 & ~n51741;
  assign n51746 = ~n51742 & n51745;
  assign n51747 = ~n51743 & n51746;
  assign n8711 = n51744 | ~n51747;
  assign n51749 = P1_P1_INSTQUEUE_REG_0__5_ & ~n51728;
  assign n51750 = n50251 & n51731;
  assign n51751 = n50253 & n51719;
  assign n51752 = n50264 & n51723;
  assign n51753 = n50276 & n51722;
  assign n51754 = ~n51749 & ~n51750;
  assign n51755 = ~n51751 & n51754;
  assign n51756 = ~n51752 & n51755;
  assign n8716 = n51753 | ~n51756;
  assign n51758 = P1_P1_INSTQUEUE_REG_0__4_ & ~n51728;
  assign n51759 = n50295 & n51731;
  assign n51760 = n50297 & n51719;
  assign n51761 = n50310 & n51723;
  assign n51762 = n50322 & n51722;
  assign n51763 = ~n51758 & ~n51759;
  assign n51764 = ~n51760 & n51763;
  assign n51765 = ~n51761 & n51764;
  assign n8721 = n51762 | ~n51765;
  assign n51767 = P1_P1_INSTQUEUE_REG_0__3_ & ~n51728;
  assign n51768 = n50339 & n51731;
  assign n51769 = n50341 & n51719;
  assign n51770 = n50353 & n51723;
  assign n51771 = n50363 & n51722;
  assign n51772 = ~n51767 & ~n51768;
  assign n51773 = ~n51769 & n51772;
  assign n51774 = ~n51770 & n51773;
  assign n8726 = n51771 | ~n51774;
  assign n51776 = P1_P1_INSTQUEUE_REG_0__2_ & ~n51728;
  assign n51777 = n50381 & n51731;
  assign n51778 = n50383 & n51719;
  assign n51779 = n50397 & n51723;
  assign n51780 = n50411 & n51722;
  assign n51781 = ~n51776 & ~n51777;
  assign n51782 = ~n51778 & n51781;
  assign n51783 = ~n51779 & n51782;
  assign n8731 = n51780 | ~n51783;
  assign n51785 = P1_P1_INSTQUEUE_REG_0__1_ & ~n51728;
  assign n51786 = n50426 & n51731;
  assign n51787 = n50428 & n51719;
  assign n51788 = n50437 & n51723;
  assign n51789 = n50449 & n51722;
  assign n51790 = ~n51785 & ~n51786;
  assign n51791 = ~n51787 & n51790;
  assign n51792 = ~n51788 & n51791;
  assign n8736 = n51789 | ~n51792;
  assign n51794 = P1_P1_INSTQUEUE_REG_0__0_ & ~n51728;
  assign n51795 = n50459 & n51731;
  assign n51796 = n50461 & n51719;
  assign n51797 = n50474 & n51723;
  assign n51798 = n50488 & n51722;
  assign n51799 = ~n51794 & ~n51795;
  assign n51800 = ~n51796 & n51799;
  assign n51801 = ~n51797 & n51800;
  assign n8741 = n51798 | ~n51801;
  assign n51803 = P1_P1_STATE2_REG_3_ & ~P1_P1_STATE2_REG_0_;
  assign n51804 = P1_P1_STATE2_REG_0_ & P1_P1_FLUSH_REG;
  assign n51805 = n43336 & n51804;
  assign n51806 = ~n51803 & ~n51805;
  assign n51807 = ~n43868 & n43979;
  assign n51808 = n51806 & ~n51807;
  assign n51809 = P1_P1_INSTQUEUERD_ADDR_REG_4_ & n51808;
  assign n51810 = ~n43911 & n43985;
  assign n51811 = n43703 & n51810;
  assign n51812 = ~n51808 & n51811;
  assign n8746 = n51809 | n51812;
  assign n51814 = ~n43902 & n43985;
  assign n51815 = ~n43375 & ~n43875;
  assign n51816 = n43994 & ~n51815;
  assign n51817 = ~n51814 & ~n51816;
  assign n51818 = ~n51808 & ~n51817;
  assign n51819 = P1_P1_INSTQUEUERD_ADDR_REG_3_ & n51808;
  assign n8751 = n51818 | n51819;
  assign n51821 = ~n43826 & n43994;
  assign n51822 = P1_P1_STATE2_REG_1_ & ~n44001;
  assign n51823 = ~n44010 & n51822;
  assign n51824 = ~n51821 & ~n51823;
  assign n51825 = ~n43842 & n43985;
  assign n51826 = n51824 & ~n51825;
  assign n51827 = ~n51808 & ~n51826;
  assign n51828 = P1_P1_INSTQUEUERD_ADDR_REG_2_ & n51808;
  assign n8756 = n51827 | n51828;
  assign n51830 = n43940 & n43994;
  assign n51831 = n44010 & n51822;
  assign n51832 = ~n51830 & ~n51831;
  assign n51833 = ~n43945 & n43985;
  assign n51834 = n51832 & ~n51833;
  assign n51835 = ~n51808 & ~n51834;
  assign n51836 = P1_P1_INSTQUEUERD_ADDR_REG_1_ & n51808;
  assign n8761 = n51835 | n51836;
  assign n51838 = P1_P1_STATE2_REG_1_ & n44001;
  assign n51839 = ~P1_P1_INSTQUEUERD_ADDR_REG_0_ & n43994;
  assign n51840 = ~n51838 & ~n51839;
  assign n51841 = ~n43932 & n43985;
  assign n51842 = n51840 & ~n51841;
  assign n51843 = ~n51808 & ~n51842;
  assign n51844 = P1_P1_INSTQUEUERD_ADDR_REG_0_ & n51808;
  assign n8766 = n51843 | n51844;
  assign n51846 = P1_P1_STATE2_REG_0_ & n43336;
  assign n51847 = ~n44024 & n51846;
  assign n51848 = ~n44042 & ~n51805;
  assign n51849 = ~n51847 & n51848;
  assign n8771 = P1_P1_INSTQUEUEWR_ADDR_REG_4_ & n51849;
  assign n51851 = P1_P1_STATE2_REG_3_ & ~n44036;
  assign n51852 = ~n51849 & ~n51851;
  assign n51853 = P1_P1_INSTQUEUEWR_ADDR_REG_3_ & ~n51852;
  assign n51854 = ~n43985 & ~n44058;
  assign n51855 = ~n44078 & ~n51854;
  assign n51856 = P1_P1_STATE2_REG_3_ & n44047;
  assign n51857 = ~n51855 & ~n51856;
  assign n51858 = n44066 & ~n44073;
  assign n51859 = ~n44084 & ~n51858;
  assign n51860 = ~n51117 & ~n51859;
  assign n51861 = n44097 & ~n51860;
  assign n51862 = n51857 & ~n51861;
  assign n51863 = ~n51849 & ~n51862;
  assign n8776 = n51853 | n51863;
  assign n51865 = ~n44069 & ~n51854;
  assign n51866 = P1_P1_STATE2_REG_3_ & ~P1_P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n51867 = n44035 & n51866;
  assign n51868 = ~n51865 & ~n51867;
  assign n51869 = ~n44066 & ~n44073;
  assign n51870 = n44066 & n44073;
  assign n51871 = ~n51869 & ~n51870;
  assign n51872 = n44097 & ~n51871;
  assign n51873 = n51868 & ~n51872;
  assign n51874 = ~n51849 & ~n51873;
  assign n51875 = P1_P1_STATE2_REG_3_ & ~n44035;
  assign n51876 = ~n51849 & ~n51875;
  assign n51877 = P1_P1_INSTQUEUEWR_ADDR_REG_2_ & ~n51876;
  assign n8781 = n51874 | n51877;
  assign n51879 = ~n44062 & ~n51854;
  assign n51880 = P1_P1_STATE2_REG_3_ & ~P1_P1_INSTQUEUEWR_ADDR_REG_1_;
  assign n51881 = ~n44065 & n44097;
  assign n51882 = ~n51880 & ~n51881;
  assign n51883 = P1_P1_INSTQUEUEWR_ADDR_REG_0_ & ~n51882;
  assign n51884 = n44097 & n50590;
  assign n51885 = ~n51879 & ~n51883;
  assign n51886 = ~n51884 & n51885;
  assign n51887 = ~n51849 & ~n51886;
  assign n51888 = P1_P1_STATE2_REG_3_ & ~P1_P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n51889 = ~n51849 & ~n51888;
  assign n51890 = P1_P1_INSTQUEUEWR_ADDR_REG_1_ & ~n51889;
  assign n8786 = n51887 | n51890;
  assign n51892 = ~n43985 & ~n44057;
  assign n51893 = ~n51849 & n51892;
  assign n51894 = P1_P1_INSTQUEUEWR_ADDR_REG_0_ & ~n51893;
  assign n51895 = ~n44025 & ~n51888;
  assign n51896 = ~n51849 & ~n51895;
  assign n8791 = n51894 | n51896;
  assign n51898 = ~P1_P1_STATE2_REG_1_ & n44057;
  assign n51899 = ~P1_P1_STATE2_REG_0_ & n51898;
  assign n51900 = n43632 & n43676;
  assign n51901 = n43630 & n43676;
  assign n51902 = ~n43464 & ~n43623;
  assign n51903 = n43721 & n51902;
  assign n51904 = ~n43860 & ~n51901;
  assign n51905 = ~n51903 & n51904;
  assign n51906 = n43681 & n43729;
  assign n51907 = n43433 & n43628;
  assign n51908 = n43676 & n51907;
  assign n51909 = ~n51906 & ~n51908;
  assign n51910 = n43592 & ~n51909;
  assign n51911 = ~n43432 & n43735;
  assign n51912 = ~n43251 & n43401;
  assign n51913 = n43676 & n51912;
  assign n51914 = ~n51911 & ~n51913;
  assign n51915 = ~n43592 & ~n51914;
  assign n51916 = n43623 & n43721;
  assign n51917 = ~n51910 & ~n51915;
  assign n51918 = ~n51916 & n51917;
  assign n51919 = n43557 & ~n51918;
  assign n51920 = n43852 & ~n51900;
  assign n51921 = n51905 & n51920;
  assign n51922 = ~n51919 & n51921;
  assign n51923 = n43979 & ~n51922;
  assign n51924 = ~n51899 & ~n51923;
  assign n51925 = P1_P1_STATE2_REG_2_ & ~n51924;
  assign n51926 = ~P1_P1_INSTADDRPOINTER_REG_0_ & n43925;
  assign n51927 = ~P1_P1_INSTADDRPOINTER_REG_0_ & n43765;
  assign n51928 = ~n51926 & ~n51927;
  assign n51929 = ~P1_P1_INSTADDRPOINTER_REG_0_ & ~n43812;
  assign n51930 = P1_P1_INSTADDRPOINTER_REG_0_ & n43883;
  assign n51931 = P1_P1_INSTADDRPOINTER_REG_0_ & n43884;
  assign n51932 = n43624 & n43755;
  assign n51933 = n43761 & n51932;
  assign n51934 = ~P1_P1_INSTADDRPOINTER_REG_0_ & n51933;
  assign n51935 = n43701 & n43755;
  assign n51936 = n43761 & n51935;
  assign n51937 = ~P1_P1_INSTADDRPOINTER_REG_0_ & n51936;
  assign n51938 = ~n51934 & ~n51937;
  assign n51939 = P1_P1_INSTADDRPOINTER_REG_0_ & n43699;
  assign n51940 = n51938 & ~n51939;
  assign n51941 = n43826 & n51815;
  assign n51942 = P1_P1_INSTQUEUERD_ADDR_REG_0_ & ~n43940;
  assign n51943 = n51941 & n51942;
  assign n51944 = P1_P1_INSTQUEUE_REG_0__0_ & n51943;
  assign n51945 = ~P1_P1_INSTQUEUERD_ADDR_REG_0_ & ~n43940;
  assign n51946 = n51941 & n51945;
  assign n51947 = P1_P1_INSTQUEUE_REG_1__0_ & n51946;
  assign n51948 = P1_P1_INSTQUEUERD_ADDR_REG_0_ & n43940;
  assign n51949 = n51941 & n51948;
  assign n51950 = P1_P1_INSTQUEUE_REG_2__0_ & n51949;
  assign n51951 = ~P1_P1_INSTQUEUERD_ADDR_REG_0_ & n43940;
  assign n51952 = n51941 & n51951;
  assign n51953 = P1_P1_INSTQUEUE_REG_3__0_ & n51952;
  assign n51954 = ~n51944 & ~n51947;
  assign n51955 = ~n51950 & n51954;
  assign n51956 = ~n51953 & n51955;
  assign n51957 = ~n43826 & n51815;
  assign n51958 = n51942 & n51957;
  assign n51959 = P1_P1_INSTQUEUE_REG_4__0_ & n51958;
  assign n51960 = n51945 & n51957;
  assign n51961 = P1_P1_INSTQUEUE_REG_5__0_ & n51960;
  assign n51962 = n51948 & n51957;
  assign n51963 = P1_P1_INSTQUEUE_REG_6__0_ & n51962;
  assign n51964 = n51951 & n51957;
  assign n51965 = P1_P1_INSTQUEUE_REG_7__0_ & n51964;
  assign n51966 = ~n51959 & ~n51961;
  assign n51967 = ~n51963 & n51966;
  assign n51968 = ~n51965 & n51967;
  assign n51969 = n43826 & ~n51815;
  assign n51970 = n51942 & n51969;
  assign n51971 = P1_P1_INSTQUEUE_REG_8__0_ & n51970;
  assign n51972 = n51945 & n51969;
  assign n51973 = P1_P1_INSTQUEUE_REG_9__0_ & n51972;
  assign n51974 = n51948 & n51969;
  assign n51975 = P1_P1_INSTQUEUE_REG_10__0_ & n51974;
  assign n51976 = n51951 & n51969;
  assign n51977 = P1_P1_INSTQUEUE_REG_11__0_ & n51976;
  assign n51978 = ~n51971 & ~n51973;
  assign n51979 = ~n51975 & n51978;
  assign n51980 = ~n51977 & n51979;
  assign n51981 = ~n43826 & ~n51815;
  assign n51982 = n51942 & n51981;
  assign n51983 = P1_P1_INSTQUEUE_REG_12__0_ & n51982;
  assign n51984 = n51945 & n51981;
  assign n51985 = P1_P1_INSTQUEUE_REG_13__0_ & n51984;
  assign n51986 = n51948 & n51981;
  assign n51987 = P1_P1_INSTQUEUE_REG_14__0_ & n51986;
  assign n51988 = n51951 & n51981;
  assign n51989 = P1_P1_INSTQUEUE_REG_15__0_ & n51988;
  assign n51990 = ~n51983 & ~n51985;
  assign n51991 = ~n51987 & n51990;
  assign n51992 = ~n51989 & n51991;
  assign n51993 = n51956 & n51968;
  assign n51994 = n51980 & n51993;
  assign n51995 = n51992 & n51994;
  assign n51996 = P1_P1_INSTADDRPOINTER_REG_0_ & n51995;
  assign n51997 = ~P1_P1_INSTADDRPOINTER_REG_0_ & ~n51995;
  assign n51998 = ~n51996 & ~n51997;
  assign n51999 = P1_P1_INSTQUEUE_REG_0__7_ & n51943;
  assign n52000 = P1_P1_INSTQUEUE_REG_1__7_ & n51946;
  assign n52001 = P1_P1_INSTQUEUE_REG_2__7_ & n51949;
  assign n52002 = P1_P1_INSTQUEUE_REG_3__7_ & n51952;
  assign n52003 = ~n51999 & ~n52000;
  assign n52004 = ~n52001 & n52003;
  assign n52005 = ~n52002 & n52004;
  assign n52006 = P1_P1_INSTQUEUE_REG_4__7_ & n51958;
  assign n52007 = P1_P1_INSTQUEUE_REG_5__7_ & n51960;
  assign n52008 = P1_P1_INSTQUEUE_REG_6__7_ & n51962;
  assign n52009 = P1_P1_INSTQUEUE_REG_7__7_ & n51964;
  assign n52010 = ~n52006 & ~n52007;
  assign n52011 = ~n52008 & n52010;
  assign n52012 = ~n52009 & n52011;
  assign n52013 = P1_P1_INSTQUEUE_REG_8__7_ & n51970;
  assign n52014 = P1_P1_INSTQUEUE_REG_9__7_ & n51972;
  assign n52015 = P1_P1_INSTQUEUE_REG_10__7_ & n51974;
  assign n52016 = P1_P1_INSTQUEUE_REG_11__7_ & n51976;
  assign n52017 = ~n52013 & ~n52014;
  assign n52018 = ~n52015 & n52017;
  assign n52019 = ~n52016 & n52018;
  assign n52020 = P1_P1_INSTQUEUE_REG_12__7_ & n51982;
  assign n52021 = P1_P1_INSTQUEUE_REG_13__7_ & n51984;
  assign n52022 = P1_P1_INSTQUEUE_REG_14__7_ & n51986;
  assign n52023 = P1_P1_INSTQUEUE_REG_15__7_ & n51988;
  assign n52024 = ~n52020 & ~n52021;
  assign n52025 = ~n52022 & n52024;
  assign n52026 = ~n52023 & n52025;
  assign n52027 = n52005 & n52012;
  assign n52028 = n52019 & n52027;
  assign n52029 = n52026 & n52028;
  assign n52030 = n43731 & ~n52029;
  assign n52031 = ~n51998 & n52030;
  assign n52032 = n43731 & n52029;
  assign n52033 = ~n51998 & n52032;
  assign n52034 = ~n51930 & ~n51931;
  assign n52035 = n51940 & n52034;
  assign n52036 = ~n52031 & n52035;
  assign n52037 = ~n52033 & n52036;
  assign n52038 = n43697 & n43725;
  assign n52039 = ~P1_P1_INSTADDRPOINTER_REG_0_ & n52038;
  assign n52040 = ~P1_P1_INSTADDRPOINTER_REG_0_ & n43769;
  assign n52041 = n43526 & n43712;
  assign n52042 = n43758 & n52041;
  assign n52043 = ~P1_P1_INSTADDRPOINTER_REG_0_ & n52042;
  assign n52044 = ~P1_P1_INSTADDRPOINTER_REG_0_ & n51995;
  assign n52045 = P1_P1_INSTADDRPOINTER_REG_0_ & ~n51995;
  assign n52046 = ~n52044 & ~n52045;
  assign n52047 = n43726 & ~n52046;
  assign n52048 = n43401 & n43755;
  assign n52049 = n43758 & n52048;
  assign n52050 = ~P1_P1_INSTADDRPOINTER_REG_0_ & n52049;
  assign n52051 = ~n52039 & ~n52040;
  assign n52052 = ~n52043 & n52051;
  assign n52053 = ~n52047 & n52052;
  assign n52054 = ~n52050 & n52053;
  assign n52055 = P1_P1_INSTADDRPOINTER_REG_0_ & n43625;
  assign n52056 = P1_P1_INSTADDRPOINTER_REG_0_ & n43703;
  assign n52057 = P1_P1_INSTADDRPOINTER_REG_0_ & n43707;
  assign n52058 = ~P1_P1_INSTADDRPOINTER_REG_0_ & n43723;
  assign n52059 = ~P1_P1_INSTADDRPOINTER_REG_0_ & n43715;
  assign n52060 = ~n52055 & ~n52056;
  assign n52061 = ~n52057 & n52060;
  assign n52062 = ~n52058 & n52061;
  assign n52063 = ~n52059 & n52062;
  assign n52064 = n52054 & n52063;
  assign n52065 = n51928 & ~n51929;
  assign n52066 = n52037 & n52065;
  assign n52067 = n52064 & n52066;
  assign n52068 = n51925 & ~n52067;
  assign n52069 = ~P1_P1_STATE2_REG_2_ & ~n51924;
  assign n52070 = P1_P1_REIP_REG_0_ & n52069;
  assign n52071 = P1_P1_INSTADDRPOINTER_REG_0_ & n51924;
  assign n52072 = ~n52068 & ~n52070;
  assign n8796 = n52071 | ~n52072;
  assign n52074 = n43925 & ~n44007;
  assign n52075 = n43765 & ~n44007;
  assign n52076 = ~n52074 & ~n52075;
  assign n52077 = ~n43812 & ~n44007;
  assign n52078 = ~P1_P1_INSTADDRPOINTER_REG_1_ & n43883;
  assign n52079 = ~P1_P1_INSTADDRPOINTER_REG_1_ & n43884;
  assign n52080 = ~n44007 & n51933;
  assign n52081 = ~n44007 & n51936;
  assign n52082 = ~n52080 & ~n52081;
  assign n52083 = ~P1_P1_INSTADDRPOINTER_REG_1_ & n43699;
  assign n52084 = n52082 & ~n52083;
  assign n52085 = ~n52078 & ~n52079;
  assign n52086 = n52084 & n52085;
  assign n52087 = P1_P1_INSTADDRPOINTER_REG_1_ & n52045;
  assign n52088 = P1_P1_INSTQUEUE_REG_0__1_ & n51943;
  assign n52089 = P1_P1_INSTQUEUE_REG_1__1_ & n51946;
  assign n52090 = P1_P1_INSTQUEUE_REG_2__1_ & n51949;
  assign n52091 = P1_P1_INSTQUEUE_REG_3__1_ & n51952;
  assign n52092 = ~n52088 & ~n52089;
  assign n52093 = ~n52090 & n52092;
  assign n52094 = ~n52091 & n52093;
  assign n52095 = P1_P1_INSTQUEUE_REG_4__1_ & n51958;
  assign n52096 = P1_P1_INSTQUEUE_REG_5__1_ & n51960;
  assign n52097 = P1_P1_INSTQUEUE_REG_6__1_ & n51962;
  assign n52098 = P1_P1_INSTQUEUE_REG_7__1_ & n51964;
  assign n52099 = ~n52095 & ~n52096;
  assign n52100 = ~n52097 & n52099;
  assign n52101 = ~n52098 & n52100;
  assign n52102 = P1_P1_INSTQUEUE_REG_8__1_ & n51970;
  assign n52103 = P1_P1_INSTQUEUE_REG_9__1_ & n51972;
  assign n52104 = P1_P1_INSTQUEUE_REG_10__1_ & n51974;
  assign n52105 = P1_P1_INSTQUEUE_REG_11__1_ & n51976;
  assign n52106 = ~n52102 & ~n52103;
  assign n52107 = ~n52104 & n52106;
  assign n52108 = ~n52105 & n52107;
  assign n52109 = P1_P1_INSTQUEUE_REG_12__1_ & n51982;
  assign n52110 = P1_P1_INSTQUEUE_REG_13__1_ & n51984;
  assign n52111 = P1_P1_INSTQUEUE_REG_14__1_ & n51986;
  assign n52112 = P1_P1_INSTQUEUE_REG_15__1_ & n51988;
  assign n52113 = ~n52109 & ~n52110;
  assign n52114 = ~n52111 & n52113;
  assign n52115 = ~n52112 & n52114;
  assign n52116 = n52094 & n52101;
  assign n52117 = n52108 & n52116;
  assign n52118 = n52115 & n52117;
  assign n52119 = n52087 & n52118;
  assign n52120 = P1_P1_INSTADDRPOINTER_REG_1_ & ~n52045;
  assign n52121 = ~n52118 & n52120;
  assign n52122 = ~n52119 & ~n52121;
  assign n52123 = n52045 & ~n52118;
  assign n52124 = ~n52045 & n52118;
  assign n52125 = ~n52123 & ~n52124;
  assign n52126 = ~P1_P1_INSTADDRPOINTER_REG_1_ & ~n52125;
  assign n52127 = n52122 & ~n52126;
  assign n52128 = n52030 & ~n52127;
  assign n52129 = ~P1_P1_INSTADDRPOINTER_REG_1_ & n52045;
  assign n52130 = ~n52120 & ~n52129;
  assign n52131 = ~n52118 & ~n52130;
  assign n52132 = ~P1_P1_INSTADDRPOINTER_REG_1_ & ~n52045;
  assign n52133 = n52118 & n52132;
  assign n52134 = n52045 & n52118;
  assign n52135 = P1_P1_INSTADDRPOINTER_REG_1_ & n52134;
  assign n52136 = ~n52131 & ~n52133;
  assign n52137 = ~n52135 & n52136;
  assign n52138 = n52032 & ~n52137;
  assign n52139 = ~n52128 & ~n52138;
  assign n52140 = ~n44007 & n52049;
  assign n52141 = ~n44007 & n52042;
  assign n52142 = ~n44007 & n52038;
  assign n52143 = n43769 & ~n44007;
  assign n52144 = ~n52140 & ~n52141;
  assign n52145 = ~n52142 & n52144;
  assign n52146 = ~n52143 & n52145;
  assign n52147 = ~P1_P1_INSTADDRPOINTER_REG_1_ & n43625;
  assign n52148 = ~P1_P1_INSTADDRPOINTER_REG_1_ & n43703;
  assign n52149 = ~P1_P1_INSTADDRPOINTER_REG_1_ & n43707;
  assign n52150 = n43723 & ~n44007;
  assign n52151 = n43715 & ~n44007;
  assign n52152 = ~n52147 & ~n52148;
  assign n52153 = ~n52149 & n52152;
  assign n52154 = ~n52150 & n52153;
  assign n52155 = ~n52151 & n52154;
  assign n52156 = ~P1_P1_INSTADDRPOINTER_REG_1_ & n51996;
  assign n52157 = P1_P1_INSTADDRPOINTER_REG_1_ & ~n51996;
  assign n52158 = ~n52156 & ~n52157;
  assign n52159 = ~n51995 & n52118;
  assign n52160 = n51995 & ~n52118;
  assign n52161 = ~n52159 & ~n52160;
  assign n52162 = ~n52158 & n52161;
  assign n52163 = ~P1_P1_INSTADDRPOINTER_REG_1_ & ~n51996;
  assign n52164 = ~n52161 & n52163;
  assign n52165 = n51996 & ~n52161;
  assign n52166 = P1_P1_INSTADDRPOINTER_REG_1_ & n52165;
  assign n52167 = ~n52162 & ~n52164;
  assign n52168 = ~n52166 & n52167;
  assign n52169 = n43726 & ~n52168;
  assign n52170 = n52146 & n52155;
  assign n52171 = ~n52169 & n52170;
  assign n52172 = n52076 & ~n52077;
  assign n52173 = n52086 & n52172;
  assign n52174 = n52139 & n52173;
  assign n52175 = n52171 & n52174;
  assign n52176 = n51925 & ~n52175;
  assign n52177 = P1_P1_REIP_REG_1_ & n52069;
  assign n52178 = P1_P1_INSTADDRPOINTER_REG_1_ & n51924;
  assign n52179 = ~n52176 & ~n52177;
  assign n8801 = n52178 | ~n52179;
  assign n52181 = P1_P1_INSTADDRPOINTER_REG_2_ & n51924;
  assign n52182 = P1_P1_REIP_REG_2_ & n52069;
  assign n52183 = P1_P1_INSTADDRPOINTER_REG_0_ & P1_P1_INSTADDRPOINTER_REG_1_;
  assign n52184 = ~P1_P1_INSTADDRPOINTER_REG_2_ & n52183;
  assign n52185 = P1_P1_INSTADDRPOINTER_REG_2_ & ~n52183;
  assign n52186 = ~n52184 & ~n52185;
  assign n52187 = ~n43812 & ~n52186;
  assign n52188 = P1_P1_INSTADDRPOINTER_REG_1_ & ~P1_P1_INSTADDRPOINTER_REG_2_;
  assign n52189 = ~P1_P1_INSTADDRPOINTER_REG_1_ & P1_P1_INSTADDRPOINTER_REG_2_;
  assign n52190 = ~n52188 & ~n52189;
  assign n52191 = n43883 & ~n52190;
  assign n52192 = n43884 & ~n52190;
  assign n52193 = n51933 & ~n52186;
  assign n52194 = n51936 & ~n52186;
  assign n52195 = ~n52193 & ~n52194;
  assign n52196 = n43699 & ~n52190;
  assign n52197 = n52195 & ~n52196;
  assign n52198 = ~n52191 & ~n52192;
  assign n52199 = n52197 & n52198;
  assign n52200 = ~n52045 & ~n52118;
  assign n52201 = P1_P1_INSTADDRPOINTER_REG_1_ & ~n52200;
  assign n52202 = ~n52134 & ~n52201;
  assign n52203 = P1_P1_INSTQUEUE_REG_0__2_ & n51943;
  assign n52204 = P1_P1_INSTQUEUE_REG_1__2_ & n51946;
  assign n52205 = P1_P1_INSTQUEUE_REG_2__2_ & n51949;
  assign n52206 = P1_P1_INSTQUEUE_REG_3__2_ & n51952;
  assign n52207 = ~n52203 & ~n52204;
  assign n52208 = ~n52205 & n52207;
  assign n52209 = ~n52206 & n52208;
  assign n52210 = P1_P1_INSTQUEUE_REG_4__2_ & n51958;
  assign n52211 = P1_P1_INSTQUEUE_REG_5__2_ & n51960;
  assign n52212 = P1_P1_INSTQUEUE_REG_6__2_ & n51962;
  assign n52213 = P1_P1_INSTQUEUE_REG_7__2_ & n51964;
  assign n52214 = ~n52210 & ~n52211;
  assign n52215 = ~n52212 & n52214;
  assign n52216 = ~n52213 & n52215;
  assign n52217 = P1_P1_INSTQUEUE_REG_8__2_ & n51970;
  assign n52218 = P1_P1_INSTQUEUE_REG_9__2_ & n51972;
  assign n52219 = P1_P1_INSTQUEUE_REG_10__2_ & n51974;
  assign n52220 = P1_P1_INSTQUEUE_REG_11__2_ & n51976;
  assign n52221 = ~n52217 & ~n52218;
  assign n52222 = ~n52219 & n52221;
  assign n52223 = ~n52220 & n52222;
  assign n52224 = P1_P1_INSTQUEUE_REG_12__2_ & n51982;
  assign n52225 = P1_P1_INSTQUEUE_REG_13__2_ & n51984;
  assign n52226 = P1_P1_INSTQUEUE_REG_14__2_ & n51986;
  assign n52227 = P1_P1_INSTQUEUE_REG_15__2_ & n51988;
  assign n52228 = ~n52224 & ~n52225;
  assign n52229 = ~n52226 & n52228;
  assign n52230 = ~n52227 & n52229;
  assign n52231 = n52209 & n52216;
  assign n52232 = n52223 & n52231;
  assign n52233 = n52230 & n52232;
  assign n52234 = ~n52118 & n52233;
  assign n52235 = n52118 & ~n52233;
  assign n52236 = ~n52234 & ~n52235;
  assign n52237 = ~P1_P1_INSTADDRPOINTER_REG_2_ & ~n52236;
  assign n52238 = P1_P1_INSTADDRPOINTER_REG_2_ & n52236;
  assign n52239 = ~n52237 & ~n52238;
  assign n52240 = n52202 & ~n52239;
  assign n52241 = ~n52202 & n52239;
  assign n52242 = ~n52240 & ~n52241;
  assign n52243 = n52032 & ~n52242;
  assign n52244 = n52049 & ~n52186;
  assign n52245 = n52042 & ~n52186;
  assign n52246 = n52038 & ~n52186;
  assign n52247 = n43769 & ~n52186;
  assign n52248 = ~n52244 & ~n52245;
  assign n52249 = ~n52246 & n52248;
  assign n52250 = ~n52247 & n52249;
  assign n52251 = n43625 & ~n52190;
  assign n52252 = n43703 & ~n52190;
  assign n52253 = n43707 & ~n52190;
  assign n52254 = ~P1_P1_INSTADDRPOINTER_REG_2_ & ~n52183;
  assign n52255 = P1_P1_INSTADDRPOINTER_REG_2_ & n52183;
  assign n52256 = ~n52254 & ~n52255;
  assign n52257 = n43723 & ~n52256;
  assign n52258 = n43715 & ~n52256;
  assign n52259 = ~n52251 & ~n52252;
  assign n52260 = ~n52253 & n52259;
  assign n52261 = ~n52257 & n52260;
  assign n52262 = ~n52258 & n52261;
  assign n52263 = ~n51995 & ~n52118;
  assign n52264 = n52233 & ~n52263;
  assign n52265 = ~n52233 & n52263;
  assign n52266 = ~n52264 & ~n52265;
  assign n52267 = ~P1_P1_INSTADDRPOINTER_REG_2_ & ~n52266;
  assign n52268 = P1_P1_INSTADDRPOINTER_REG_2_ & n52266;
  assign n52269 = ~n52267 & ~n52268;
  assign n52270 = ~n51996 & n52161;
  assign n52271 = P1_P1_INSTADDRPOINTER_REG_1_ & ~n52270;
  assign n52272 = ~n52165 & ~n52271;
  assign n52273 = ~n52269 & n52272;
  assign n52274 = ~P1_P1_INSTADDRPOINTER_REG_2_ & n52266;
  assign n52275 = P1_P1_INSTADDRPOINTER_REG_2_ & ~n52266;
  assign n52276 = ~n52274 & ~n52275;
  assign n52277 = ~n52272 & ~n52276;
  assign n52278 = ~n52273 & ~n52277;
  assign n52279 = n43726 & ~n52278;
  assign n52280 = n52250 & n52262;
  assign n52281 = ~n52279 & n52280;
  assign n52282 = n43925 & ~n52186;
  assign n52283 = n43765 & ~n52186;
  assign n52284 = ~n52282 & ~n52283;
  assign n52285 = P1_P1_INSTADDRPOINTER_REG_1_ & n52118;
  assign n52286 = ~n52087 & ~n52134;
  assign n52287 = ~n52285 & n52286;
  assign n52288 = ~n52239 & n52287;
  assign n52289 = ~P1_P1_INSTADDRPOINTER_REG_2_ & n52236;
  assign n52290 = P1_P1_INSTADDRPOINTER_REG_2_ & ~n52236;
  assign n52291 = ~n52289 & ~n52290;
  assign n52292 = ~n52287 & ~n52291;
  assign n52293 = ~n52288 & ~n52292;
  assign n52294 = n52030 & ~n52293;
  assign n52295 = n52284 & ~n52294;
  assign n52296 = ~n52187 & n52199;
  assign n52297 = ~n52243 & n52296;
  assign n52298 = n52281 & n52297;
  assign n52299 = n52295 & n52298;
  assign n52300 = n51925 & ~n52299;
  assign n52301 = ~n52181 & ~n52182;
  assign n8806 = n52300 | ~n52301;
  assign n52303 = P1_P1_INSTADDRPOINTER_REG_3_ & n51924;
  assign n52304 = P1_P1_REIP_REG_3_ & n52069;
  assign n52305 = ~P1_P1_INSTADDRPOINTER_REG_3_ & n52255;
  assign n52306 = P1_P1_INSTADDRPOINTER_REG_3_ & ~n52255;
  assign n52307 = ~n52305 & ~n52306;
  assign n52308 = ~n43812 & ~n52307;
  assign n52309 = P1_P1_INSTADDRPOINTER_REG_1_ & P1_P1_INSTADDRPOINTER_REG_2_;
  assign n52310 = ~P1_P1_INSTADDRPOINTER_REG_3_ & n52309;
  assign n52311 = P1_P1_INSTADDRPOINTER_REG_3_ & ~n52309;
  assign n52312 = ~n52310 & ~n52311;
  assign n52313 = n43883 & ~n52312;
  assign n52314 = n43884 & ~n52312;
  assign n52315 = n51933 & ~n52307;
  assign n52316 = n51936 & ~n52307;
  assign n52317 = ~n52315 & ~n52316;
  assign n52318 = n43699 & ~n52312;
  assign n52319 = n52317 & ~n52318;
  assign n52320 = ~n52313 & ~n52314;
  assign n52321 = n52319 & n52320;
  assign n52322 = ~n52202 & ~n52289;
  assign n52323 = ~n52290 & ~n52322;
  assign n52324 = ~n52118 & ~n52233;
  assign n52325 = P1_P1_INSTQUEUE_REG_0__3_ & n51943;
  assign n52326 = P1_P1_INSTQUEUE_REG_1__3_ & n51946;
  assign n52327 = P1_P1_INSTQUEUE_REG_2__3_ & n51949;
  assign n52328 = P1_P1_INSTQUEUE_REG_3__3_ & n51952;
  assign n52329 = ~n52325 & ~n52326;
  assign n52330 = ~n52327 & n52329;
  assign n52331 = ~n52328 & n52330;
  assign n52332 = P1_P1_INSTQUEUE_REG_4__3_ & n51958;
  assign n52333 = P1_P1_INSTQUEUE_REG_5__3_ & n51960;
  assign n52334 = P1_P1_INSTQUEUE_REG_6__3_ & n51962;
  assign n52335 = P1_P1_INSTQUEUE_REG_7__3_ & n51964;
  assign n52336 = ~n52332 & ~n52333;
  assign n52337 = ~n52334 & n52336;
  assign n52338 = ~n52335 & n52337;
  assign n52339 = P1_P1_INSTQUEUE_REG_8__3_ & n51970;
  assign n52340 = P1_P1_INSTQUEUE_REG_9__3_ & n51972;
  assign n52341 = P1_P1_INSTQUEUE_REG_10__3_ & n51974;
  assign n52342 = P1_P1_INSTQUEUE_REG_11__3_ & n51976;
  assign n52343 = ~n52339 & ~n52340;
  assign n52344 = ~n52341 & n52343;
  assign n52345 = ~n52342 & n52344;
  assign n52346 = P1_P1_INSTQUEUE_REG_12__3_ & n51982;
  assign n52347 = P1_P1_INSTQUEUE_REG_13__3_ & n51984;
  assign n52348 = P1_P1_INSTQUEUE_REG_14__3_ & n51986;
  assign n52349 = P1_P1_INSTQUEUE_REG_15__3_ & n51988;
  assign n52350 = ~n52346 & ~n52347;
  assign n52351 = ~n52348 & n52350;
  assign n52352 = ~n52349 & n52351;
  assign n52353 = n52331 & n52338;
  assign n52354 = n52345 & n52353;
  assign n52355 = n52352 & n52354;
  assign n52356 = n52324 & n52355;
  assign n52357 = ~n52324 & ~n52355;
  assign n52358 = ~n52356 & ~n52357;
  assign n52359 = ~P1_P1_INSTADDRPOINTER_REG_3_ & n52358;
  assign n52360 = ~n52323 & ~n52359;
  assign n52361 = P1_P1_INSTADDRPOINTER_REG_3_ & ~n52358;
  assign n52362 = n52360 & ~n52361;
  assign n52363 = ~P1_P1_INSTADDRPOINTER_REG_3_ & ~n52358;
  assign n52364 = P1_P1_INSTADDRPOINTER_REG_3_ & n52358;
  assign n52365 = ~n52363 & ~n52364;
  assign n52366 = n52323 & n52365;
  assign n52367 = ~n52362 & ~n52366;
  assign n52368 = n52032 & n52367;
  assign n52369 = n43925 & ~n52307;
  assign n52370 = n43765 & ~n52307;
  assign n52371 = ~n52369 & ~n52370;
  assign n52372 = ~n52287 & ~n52289;
  assign n52373 = ~n52290 & ~n52372;
  assign n52374 = ~n52324 & n52355;
  assign n52375 = n52324 & ~n52355;
  assign n52376 = ~n52374 & ~n52375;
  assign n52377 = P1_P1_INSTADDRPOINTER_REG_3_ & ~n52376;
  assign n52378 = ~P1_P1_INSTADDRPOINTER_REG_3_ & n52376;
  assign n52379 = ~n52377 & ~n52378;
  assign n52380 = n52373 & ~n52379;
  assign n52381 = P1_P1_INSTADDRPOINTER_REG_3_ & n52376;
  assign n52382 = ~P1_P1_INSTADDRPOINTER_REG_3_ & ~n52376;
  assign n52383 = ~n52381 & ~n52382;
  assign n52384 = ~n52373 & ~n52383;
  assign n52385 = ~n52380 & ~n52384;
  assign n52386 = n52030 & ~n52385;
  assign n52387 = n52371 & ~n52386;
  assign n52388 = n52049 & ~n52307;
  assign n52389 = n52042 & ~n52307;
  assign n52390 = n52038 & ~n52307;
  assign n52391 = n43769 & ~n52307;
  assign n52392 = ~n52388 & ~n52389;
  assign n52393 = ~n52390 & n52392;
  assign n52394 = ~n52391 & n52393;
  assign n52395 = n43625 & ~n52312;
  assign n52396 = n43703 & ~n52312;
  assign n52397 = n43707 & ~n52312;
  assign n52398 = ~P1_P1_INSTADDRPOINTER_REG_3_ & n52254;
  assign n52399 = P1_P1_INSTADDRPOINTER_REG_3_ & ~n52254;
  assign n52400 = ~n52398 & ~n52399;
  assign n52401 = n43723 & n52400;
  assign n52402 = n43715 & n52400;
  assign n52403 = ~n52395 & ~n52396;
  assign n52404 = ~n52397 & n52403;
  assign n52405 = ~n52401 & n52404;
  assign n52406 = ~n52402 & n52405;
  assign n52407 = n52272 & ~n52275;
  assign n52408 = n52264 & n52355;
  assign n52409 = ~n52264 & ~n52355;
  assign n52410 = ~n52408 & ~n52409;
  assign n52411 = P1_P1_INSTADDRPOINTER_REG_3_ & n52410;
  assign n52412 = ~n52274 & n52410;
  assign n52413 = P1_P1_INSTADDRPOINTER_REG_3_ & ~n52274;
  assign n52414 = ~n52412 & ~n52413;
  assign n52415 = ~n52407 & ~n52411;
  assign n52416 = ~n52414 & n52415;
  assign n52417 = ~P1_P1_INSTADDRPOINTER_REG_3_ & n52410;
  assign n52418 = P1_P1_INSTADDRPOINTER_REG_3_ & ~n52410;
  assign n52419 = ~n52417 & ~n52418;
  assign n52420 = ~n52275 & n52419;
  assign n52421 = ~n52272 & ~n52274;
  assign n52422 = n52420 & ~n52421;
  assign n52423 = ~n52416 & ~n52422;
  assign n52424 = n43726 & n52423;
  assign n52425 = n52394 & n52406;
  assign n52426 = ~n52424 & n52425;
  assign n52427 = ~n52308 & n52321;
  assign n52428 = ~n52368 & n52427;
  assign n52429 = n52387 & n52428;
  assign n52430 = n52426 & n52429;
  assign n52431 = n51925 & ~n52430;
  assign n52432 = ~n52303 & ~n52304;
  assign n8811 = n52431 | ~n52432;
  assign n52434 = P1_P1_INSTADDRPOINTER_REG_4_ & n51924;
  assign n52435 = P1_P1_REIP_REG_4_ & n52069;
  assign n52436 = P1_P1_INSTADDRPOINTER_REG_3_ & n52255;
  assign n52437 = ~P1_P1_INSTADDRPOINTER_REG_4_ & n52436;
  assign n52438 = P1_P1_INSTADDRPOINTER_REG_4_ & ~n52436;
  assign n52439 = ~n52437 & ~n52438;
  assign n52440 = ~n43812 & ~n52439;
  assign n52441 = P1_P1_INSTADDRPOINTER_REG_3_ & n52309;
  assign n52442 = ~P1_P1_INSTADDRPOINTER_REG_4_ & n52441;
  assign n52443 = P1_P1_INSTADDRPOINTER_REG_4_ & ~n52441;
  assign n52444 = ~n52442 & ~n52443;
  assign n52445 = n43883 & ~n52444;
  assign n52446 = n43884 & ~n52444;
  assign n52447 = n51933 & ~n52439;
  assign n52448 = n51936 & ~n52439;
  assign n52449 = ~n52447 & ~n52448;
  assign n52450 = n43699 & ~n52444;
  assign n52451 = n52449 & ~n52450;
  assign n52452 = ~n52445 & ~n52446;
  assign n52453 = n52451 & n52452;
  assign n52454 = P1_P1_INSTQUEUE_REG_0__4_ & n51943;
  assign n52455 = P1_P1_INSTQUEUE_REG_1__4_ & n51946;
  assign n52456 = P1_P1_INSTQUEUE_REG_2__4_ & n51949;
  assign n52457 = P1_P1_INSTQUEUE_REG_3__4_ & n51952;
  assign n52458 = ~n52454 & ~n52455;
  assign n52459 = ~n52456 & n52458;
  assign n52460 = ~n52457 & n52459;
  assign n52461 = P1_P1_INSTQUEUE_REG_4__4_ & n51958;
  assign n52462 = P1_P1_INSTQUEUE_REG_5__4_ & n51960;
  assign n52463 = P1_P1_INSTQUEUE_REG_6__4_ & n51962;
  assign n52464 = P1_P1_INSTQUEUE_REG_7__4_ & n51964;
  assign n52465 = ~n52461 & ~n52462;
  assign n52466 = ~n52463 & n52465;
  assign n52467 = ~n52464 & n52466;
  assign n52468 = P1_P1_INSTQUEUE_REG_8__4_ & n51970;
  assign n52469 = P1_P1_INSTQUEUE_REG_9__4_ & n51972;
  assign n52470 = P1_P1_INSTQUEUE_REG_10__4_ & n51974;
  assign n52471 = P1_P1_INSTQUEUE_REG_11__4_ & n51976;
  assign n52472 = ~n52468 & ~n52469;
  assign n52473 = ~n52470 & n52472;
  assign n52474 = ~n52471 & n52473;
  assign n52475 = P1_P1_INSTQUEUE_REG_12__4_ & n51982;
  assign n52476 = P1_P1_INSTQUEUE_REG_13__4_ & n51984;
  assign n52477 = P1_P1_INSTQUEUE_REG_14__4_ & n51986;
  assign n52478 = P1_P1_INSTQUEUE_REG_15__4_ & n51988;
  assign n52479 = ~n52475 & ~n52476;
  assign n52480 = ~n52477 & n52479;
  assign n52481 = ~n52478 & n52480;
  assign n52482 = n52460 & n52467;
  assign n52483 = n52474 & n52482;
  assign n52484 = n52481 & n52483;
  assign n52485 = n52375 & n52484;
  assign n52486 = ~n52375 & ~n52484;
  assign n52487 = ~n52485 & ~n52486;
  assign n52488 = P1_P1_INSTADDRPOINTER_REG_4_ & ~n52487;
  assign n52489 = ~P1_P1_INSTADDRPOINTER_REG_4_ & n52487;
  assign n52490 = ~n52488 & ~n52489;
  assign n52491 = ~n52360 & ~n52361;
  assign n52492 = n52490 & ~n52491;
  assign n52493 = ~P1_P1_INSTADDRPOINTER_REG_4_ & ~n52487;
  assign n52494 = P1_P1_INSTADDRPOINTER_REG_4_ & n52487;
  assign n52495 = ~n52493 & ~n52494;
  assign n52496 = ~n52361 & n52495;
  assign n52497 = ~n52360 & n52496;
  assign n52498 = ~n52492 & ~n52497;
  assign n52499 = n52032 & n52498;
  assign n52500 = n43925 & ~n52439;
  assign n52501 = n43765 & ~n52439;
  assign n52502 = ~n52500 & ~n52501;
  assign n52503 = ~n52289 & ~n52382;
  assign n52504 = ~n52134 & ~n52285;
  assign n52505 = ~n52290 & n52504;
  assign n52506 = ~n52087 & n52505;
  assign n52507 = n52503 & ~n52506;
  assign n52508 = ~n52381 & ~n52507;
  assign n52509 = n52375 & ~n52484;
  assign n52510 = ~n52375 & n52484;
  assign n52511 = ~n52509 & ~n52510;
  assign n52512 = P1_P1_INSTADDRPOINTER_REG_4_ & ~n52511;
  assign n52513 = ~P1_P1_INSTADDRPOINTER_REG_4_ & n52511;
  assign n52514 = ~n52512 & ~n52513;
  assign n52515 = n52508 & ~n52514;
  assign n52516 = P1_P1_INSTADDRPOINTER_REG_4_ & n52511;
  assign n52517 = ~P1_P1_INSTADDRPOINTER_REG_4_ & ~n52511;
  assign n52518 = ~n52516 & ~n52517;
  assign n52519 = ~n52508 & ~n52518;
  assign n52520 = ~n52515 & ~n52519;
  assign n52521 = n52030 & ~n52520;
  assign n52522 = n52502 & ~n52521;
  assign n52523 = n52049 & ~n52439;
  assign n52524 = n52042 & ~n52439;
  assign n52525 = n52038 & ~n52439;
  assign n52526 = n43769 & ~n52439;
  assign n52527 = ~n52523 & ~n52524;
  assign n52528 = ~n52525 & n52527;
  assign n52529 = ~n52526 & n52528;
  assign n52530 = n43625 & ~n52444;
  assign n52531 = n43703 & ~n52444;
  assign n52532 = n43707 & ~n52444;
  assign n52533 = ~P1_P1_INSTADDRPOINTER_REG_4_ & n52399;
  assign n52534 = P1_P1_INSTADDRPOINTER_REG_4_ & ~n52399;
  assign n52535 = ~n52533 & ~n52534;
  assign n52536 = n43723 & ~n52535;
  assign n52537 = n43715 & ~n52535;
  assign n52538 = ~n52530 & ~n52531;
  assign n52539 = ~n52532 & n52538;
  assign n52540 = ~n52536 & n52539;
  assign n52541 = ~n52537 & n52540;
  assign n52542 = n52409 & n52484;
  assign n52543 = ~n52409 & ~n52484;
  assign n52544 = ~n52542 & ~n52543;
  assign n52545 = ~P1_P1_INSTADDRPOINTER_REG_4_ & ~n52544;
  assign n52546 = P1_P1_INSTADDRPOINTER_REG_4_ & n52544;
  assign n52547 = ~n52545 & ~n52546;
  assign n52548 = n52275 & n52410;
  assign n52549 = ~n52275 & ~n52410;
  assign n52550 = P1_P1_INSTADDRPOINTER_REG_3_ & ~n52549;
  assign n52551 = ~n52548 & ~n52550;
  assign n52552 = ~n52272 & ~n52414;
  assign n52553 = n52551 & ~n52552;
  assign n52554 = ~n52547 & n52553;
  assign n52555 = ~P1_P1_INSTADDRPOINTER_REG_4_ & n52544;
  assign n52556 = P1_P1_INSTADDRPOINTER_REG_4_ & ~n52544;
  assign n52557 = ~n52555 & ~n52556;
  assign n52558 = ~n52553 & ~n52557;
  assign n52559 = ~n52554 & ~n52558;
  assign n52560 = n43726 & ~n52559;
  assign n52561 = n52529 & n52541;
  assign n52562 = ~n52560 & n52561;
  assign n52563 = ~n52440 & n52453;
  assign n52564 = ~n52499 & n52563;
  assign n52565 = n52522 & n52564;
  assign n52566 = n52562 & n52565;
  assign n52567 = n51925 & ~n52566;
  assign n52568 = ~n52434 & ~n52435;
  assign n8816 = n52567 | ~n52568;
  assign n52570 = P1_P1_INSTADDRPOINTER_REG_5_ & n51924;
  assign n52571 = P1_P1_REIP_REG_5_ & n52069;
  assign n52572 = P1_P1_INSTADDRPOINTER_REG_4_ & n52436;
  assign n52573 = ~P1_P1_INSTADDRPOINTER_REG_5_ & n52572;
  assign n52574 = P1_P1_INSTADDRPOINTER_REG_5_ & ~n52572;
  assign n52575 = ~n52573 & ~n52574;
  assign n52576 = ~n43812 & ~n52575;
  assign n52577 = P1_P1_INSTADDRPOINTER_REG_4_ & n52441;
  assign n52578 = ~P1_P1_INSTADDRPOINTER_REG_5_ & n52577;
  assign n52579 = P1_P1_INSTADDRPOINTER_REG_5_ & ~n52577;
  assign n52580 = ~n52578 & ~n52579;
  assign n52581 = n43883 & ~n52580;
  assign n52582 = n43884 & ~n52580;
  assign n52583 = n51933 & ~n52575;
  assign n52584 = n51936 & ~n52575;
  assign n52585 = ~n52583 & ~n52584;
  assign n52586 = n43699 & ~n52580;
  assign n52587 = n52585 & ~n52586;
  assign n52588 = ~n52581 & ~n52582;
  assign n52589 = n52587 & n52588;
  assign n52590 = n52361 & ~n52489;
  assign n52591 = ~n52488 & ~n52590;
  assign n52592 = ~n52359 & ~n52489;
  assign n52593 = ~n52323 & n52592;
  assign n52594 = n52591 & ~n52593;
  assign n52595 = P1_P1_INSTQUEUE_REG_0__5_ & n51943;
  assign n52596 = P1_P1_INSTQUEUE_REG_1__5_ & n51946;
  assign n52597 = P1_P1_INSTQUEUE_REG_2__5_ & n51949;
  assign n52598 = P1_P1_INSTQUEUE_REG_3__5_ & n51952;
  assign n52599 = ~n52595 & ~n52596;
  assign n52600 = ~n52597 & n52599;
  assign n52601 = ~n52598 & n52600;
  assign n52602 = P1_P1_INSTQUEUE_REG_4__5_ & n51958;
  assign n52603 = P1_P1_INSTQUEUE_REG_5__5_ & n51960;
  assign n52604 = P1_P1_INSTQUEUE_REG_6__5_ & n51962;
  assign n52605 = P1_P1_INSTQUEUE_REG_7__5_ & n51964;
  assign n52606 = ~n52602 & ~n52603;
  assign n52607 = ~n52604 & n52606;
  assign n52608 = ~n52605 & n52607;
  assign n52609 = P1_P1_INSTQUEUE_REG_8__5_ & n51970;
  assign n52610 = P1_P1_INSTQUEUE_REG_9__5_ & n51972;
  assign n52611 = P1_P1_INSTQUEUE_REG_10__5_ & n51974;
  assign n52612 = P1_P1_INSTQUEUE_REG_11__5_ & n51976;
  assign n52613 = ~n52609 & ~n52610;
  assign n52614 = ~n52611 & n52613;
  assign n52615 = ~n52612 & n52614;
  assign n52616 = P1_P1_INSTQUEUE_REG_12__5_ & n51982;
  assign n52617 = P1_P1_INSTQUEUE_REG_13__5_ & n51984;
  assign n52618 = P1_P1_INSTQUEUE_REG_14__5_ & n51986;
  assign n52619 = P1_P1_INSTQUEUE_REG_15__5_ & n51988;
  assign n52620 = ~n52616 & ~n52617;
  assign n52621 = ~n52618 & n52620;
  assign n52622 = ~n52619 & n52621;
  assign n52623 = n52601 & n52608;
  assign n52624 = n52615 & n52623;
  assign n52625 = n52622 & n52624;
  assign n52626 = n52509 & n52625;
  assign n52627 = ~n52509 & ~n52625;
  assign n52628 = ~n52626 & ~n52627;
  assign n52629 = ~P1_P1_INSTADDRPOINTER_REG_5_ & ~n52628;
  assign n52630 = P1_P1_INSTADDRPOINTER_REG_5_ & n52628;
  assign n52631 = ~n52629 & ~n52630;
  assign n52632 = n52594 & ~n52631;
  assign n52633 = ~n52594 & n52631;
  assign n52634 = ~n52632 & ~n52633;
  assign n52635 = n52032 & ~n52634;
  assign n52636 = n43925 & ~n52575;
  assign n52637 = n43765 & ~n52575;
  assign n52638 = ~n52636 & ~n52637;
  assign n52639 = n52381 & ~n52517;
  assign n52640 = ~n52516 & ~n52639;
  assign n52641 = n52503 & ~n52517;
  assign n52642 = ~n52506 & n52641;
  assign n52643 = n52640 & ~n52642;
  assign n52644 = ~n52509 & n52625;
  assign n52645 = ~n52484 & ~n52625;
  assign n52646 = n52375 & n52645;
  assign n52647 = ~n52644 & ~n52646;
  assign n52648 = P1_P1_INSTADDRPOINTER_REG_5_ & ~n52647;
  assign n52649 = ~P1_P1_INSTADDRPOINTER_REG_5_ & n52647;
  assign n52650 = ~n52648 & ~n52649;
  assign n52651 = n52643 & ~n52650;
  assign n52652 = ~n52643 & n52650;
  assign n52653 = ~n52651 & ~n52652;
  assign n52654 = n52030 & ~n52653;
  assign n52655 = n52638 & ~n52654;
  assign n52656 = n52049 & ~n52575;
  assign n52657 = n52042 & ~n52575;
  assign n52658 = n52038 & ~n52575;
  assign n52659 = n43769 & ~n52575;
  assign n52660 = ~n52656 & ~n52657;
  assign n52661 = ~n52658 & n52660;
  assign n52662 = ~n52659 & n52661;
  assign n52663 = n43625 & ~n52580;
  assign n52664 = n43703 & ~n52580;
  assign n52665 = n43707 & ~n52580;
  assign n52666 = P1_P1_INSTADDRPOINTER_REG_4_ & n52399;
  assign n52667 = ~P1_P1_INSTADDRPOINTER_REG_5_ & n52666;
  assign n52668 = P1_P1_INSTADDRPOINTER_REG_5_ & ~n52666;
  assign n52669 = ~n52667 & ~n52668;
  assign n52670 = n43723 & ~n52669;
  assign n52671 = n43715 & ~n52669;
  assign n52672 = ~n52663 & ~n52664;
  assign n52673 = ~n52665 & n52672;
  assign n52674 = ~n52670 & n52673;
  assign n52675 = ~n52671 & n52674;
  assign n52676 = n52409 & ~n52484;
  assign n52677 = n52625 & n52676;
  assign n52678 = ~n52625 & ~n52676;
  assign n52679 = ~n52677 & ~n52678;
  assign n52680 = P1_P1_INSTADDRPOINTER_REG_5_ & ~n52679;
  assign n52681 = ~P1_P1_INSTADDRPOINTER_REG_5_ & n52679;
  assign n52682 = ~n52555 & ~n52681;
  assign n52683 = ~n52680 & n52682;
  assign n52684 = n52553 & ~n52556;
  assign n52685 = n52683 & ~n52684;
  assign n52686 = ~P1_P1_INSTADDRPOINTER_REG_5_ & ~n52679;
  assign n52687 = P1_P1_INSTADDRPOINTER_REG_5_ & n52679;
  assign n52688 = ~n52686 & ~n52687;
  assign n52689 = ~n52556 & n52688;
  assign n52690 = ~n52553 & ~n52555;
  assign n52691 = n52689 & ~n52690;
  assign n52692 = ~n52685 & ~n52691;
  assign n52693 = n43726 & n52692;
  assign n52694 = n52662 & n52675;
  assign n52695 = ~n52693 & n52694;
  assign n52696 = ~n52576 & n52589;
  assign n52697 = ~n52635 & n52696;
  assign n52698 = n52655 & n52697;
  assign n52699 = n52695 & n52698;
  assign n52700 = n51925 & ~n52699;
  assign n52701 = ~n52570 & ~n52571;
  assign n8821 = n52700 | ~n52701;
  assign n52703 = P1_P1_INSTADDRPOINTER_REG_6_ & n51924;
  assign n52704 = P1_P1_REIP_REG_6_ & n52069;
  assign n52705 = P1_P1_INSTADDRPOINTER_REG_5_ & n52572;
  assign n52706 = ~P1_P1_INSTADDRPOINTER_REG_6_ & n52705;
  assign n52707 = P1_P1_INSTADDRPOINTER_REG_6_ & ~n52705;
  assign n52708 = ~n52706 & ~n52707;
  assign n52709 = ~n43812 & ~n52708;
  assign n52710 = P1_P1_INSTADDRPOINTER_REG_5_ & n52577;
  assign n52711 = ~P1_P1_INSTADDRPOINTER_REG_6_ & n52710;
  assign n52712 = P1_P1_INSTADDRPOINTER_REG_6_ & ~n52710;
  assign n52713 = ~n52711 & ~n52712;
  assign n52714 = n43883 & ~n52713;
  assign n52715 = n43884 & ~n52713;
  assign n52716 = n51933 & ~n52708;
  assign n52717 = n51936 & ~n52708;
  assign n52718 = ~n52716 & ~n52717;
  assign n52719 = n43699 & ~n52713;
  assign n52720 = n52718 & ~n52719;
  assign n52721 = ~n52714 & ~n52715;
  assign n52722 = n52720 & n52721;
  assign n52723 = ~n52594 & ~n52628;
  assign n52724 = P1_P1_INSTADDRPOINTER_REG_5_ & ~n52594;
  assign n52725 = P1_P1_INSTADDRPOINTER_REG_5_ & ~n52628;
  assign n52726 = ~n52723 & ~n52724;
  assign n52727 = ~n52725 & n52726;
  assign n52728 = n52509 & ~n52625;
  assign n52729 = P1_P1_INSTQUEUE_REG_0__6_ & n51943;
  assign n52730 = P1_P1_INSTQUEUE_REG_1__6_ & n51946;
  assign n52731 = P1_P1_INSTQUEUE_REG_2__6_ & n51949;
  assign n52732 = P1_P1_INSTQUEUE_REG_3__6_ & n51952;
  assign n52733 = ~n52729 & ~n52730;
  assign n52734 = ~n52731 & n52733;
  assign n52735 = ~n52732 & n52734;
  assign n52736 = P1_P1_INSTQUEUE_REG_4__6_ & n51958;
  assign n52737 = P1_P1_INSTQUEUE_REG_5__6_ & n51960;
  assign n52738 = P1_P1_INSTQUEUE_REG_6__6_ & n51962;
  assign n52739 = P1_P1_INSTQUEUE_REG_7__6_ & n51964;
  assign n52740 = ~n52736 & ~n52737;
  assign n52741 = ~n52738 & n52740;
  assign n52742 = ~n52739 & n52741;
  assign n52743 = P1_P1_INSTQUEUE_REG_8__6_ & n51970;
  assign n52744 = P1_P1_INSTQUEUE_REG_9__6_ & n51972;
  assign n52745 = P1_P1_INSTQUEUE_REG_10__6_ & n51974;
  assign n52746 = P1_P1_INSTQUEUE_REG_11__6_ & n51976;
  assign n52747 = ~n52743 & ~n52744;
  assign n52748 = ~n52745 & n52747;
  assign n52749 = ~n52746 & n52748;
  assign n52750 = P1_P1_INSTQUEUE_REG_12__6_ & n51982;
  assign n52751 = P1_P1_INSTQUEUE_REG_13__6_ & n51984;
  assign n52752 = P1_P1_INSTQUEUE_REG_14__6_ & n51986;
  assign n52753 = P1_P1_INSTQUEUE_REG_15__6_ & n51988;
  assign n52754 = ~n52750 & ~n52751;
  assign n52755 = ~n52752 & n52754;
  assign n52756 = ~n52753 & n52755;
  assign n52757 = n52735 & n52742;
  assign n52758 = n52749 & n52757;
  assign n52759 = n52756 & n52758;
  assign n52760 = n52728 & n52759;
  assign n52761 = ~n52728 & ~n52759;
  assign n52762 = ~n52760 & ~n52761;
  assign n52763 = ~P1_P1_INSTADDRPOINTER_REG_6_ & ~n52762;
  assign n52764 = P1_P1_INSTADDRPOINTER_REG_6_ & n52762;
  assign n52765 = ~n52763 & ~n52764;
  assign n52766 = n52727 & ~n52765;
  assign n52767 = ~n52727 & n52765;
  assign n52768 = ~n52766 & ~n52767;
  assign n52769 = n52032 & ~n52768;
  assign n52770 = n52049 & ~n52708;
  assign n52771 = n52042 & ~n52708;
  assign n52772 = n52038 & ~n52708;
  assign n52773 = n43769 & ~n52708;
  assign n52774 = ~n52770 & ~n52771;
  assign n52775 = ~n52772 & n52774;
  assign n52776 = ~n52773 & n52775;
  assign n52777 = n43625 & ~n52713;
  assign n52778 = n43703 & ~n52713;
  assign n52779 = n43707 & ~n52713;
  assign n52780 = P1_P1_INSTADDRPOINTER_REG_5_ & n52666;
  assign n52781 = ~P1_P1_INSTADDRPOINTER_REG_6_ & n52780;
  assign n52782 = P1_P1_INSTADDRPOINTER_REG_6_ & ~n52780;
  assign n52783 = ~n52781 & ~n52782;
  assign n52784 = n43723 & ~n52783;
  assign n52785 = n43715 & ~n52783;
  assign n52786 = ~n52777 & ~n52778;
  assign n52787 = ~n52779 & n52786;
  assign n52788 = ~n52784 & n52787;
  assign n52789 = ~n52785 & n52788;
  assign n52790 = n52556 & ~n52679;
  assign n52791 = ~n52556 & n52679;
  assign n52792 = P1_P1_INSTADDRPOINTER_REG_5_ & ~n52791;
  assign n52793 = ~n52790 & ~n52792;
  assign n52794 = ~n52553 & n52682;
  assign n52795 = n52793 & ~n52794;
  assign n52796 = ~n52625 & n52676;
  assign n52797 = n52759 & n52796;
  assign n52798 = ~n52759 & ~n52796;
  assign n52799 = ~n52797 & ~n52798;
  assign n52800 = ~P1_P1_INSTADDRPOINTER_REG_6_ & ~n52799;
  assign n52801 = P1_P1_INSTADDRPOINTER_REG_6_ & n52799;
  assign n52802 = ~n52800 & ~n52801;
  assign n52803 = n52795 & ~n52802;
  assign n52804 = ~n52795 & n52802;
  assign n52805 = ~n52803 & ~n52804;
  assign n52806 = n43726 & ~n52805;
  assign n52807 = n43925 & ~n52708;
  assign n52808 = n43765 & ~n52708;
  assign n52809 = ~n52807 & ~n52808;
  assign n52810 = P1_P1_INSTADDRPOINTER_REG_5_ & ~n52643;
  assign n52811 = ~n52643 & n52647;
  assign n52812 = P1_P1_INSTADDRPOINTER_REG_5_ & n52647;
  assign n52813 = ~n52810 & ~n52811;
  assign n52814 = ~n52812 & n52813;
  assign n52815 = n52646 & ~n52759;
  assign n52816 = ~n52646 & n52759;
  assign n52817 = ~n52815 & ~n52816;
  assign n52818 = P1_P1_INSTADDRPOINTER_REG_6_ & ~n52817;
  assign n52819 = ~P1_P1_INSTADDRPOINTER_REG_6_ & n52817;
  assign n52820 = ~n52818 & ~n52819;
  assign n52821 = n52814 & ~n52820;
  assign n52822 = ~n52814 & n52820;
  assign n52823 = ~n52821 & ~n52822;
  assign n52824 = n52030 & ~n52823;
  assign n52825 = n52776 & n52789;
  assign n52826 = ~n52806 & n52825;
  assign n52827 = n52809 & n52826;
  assign n52828 = ~n52824 & n52827;
  assign n52829 = ~n52709 & n52722;
  assign n52830 = ~n52769 & n52829;
  assign n52831 = n52828 & n52830;
  assign n52832 = n51925 & ~n52831;
  assign n52833 = ~n52703 & ~n52704;
  assign n8826 = n52832 | ~n52833;
  assign n52835 = P1_P1_INSTADDRPOINTER_REG_7_ & n51924;
  assign n52836 = P1_P1_REIP_REG_7_ & n52069;
  assign n52837 = P1_P1_INSTADDRPOINTER_REG_6_ & n52705;
  assign n52838 = ~P1_P1_INSTADDRPOINTER_REG_7_ & n52837;
  assign n52839 = P1_P1_INSTADDRPOINTER_REG_7_ & ~n52837;
  assign n52840 = ~n52838 & ~n52839;
  assign n52841 = ~n43812 & ~n52840;
  assign n52842 = P1_P1_INSTADDRPOINTER_REG_6_ & n52710;
  assign n52843 = ~P1_P1_INSTADDRPOINTER_REG_7_ & n52842;
  assign n52844 = P1_P1_INSTADDRPOINTER_REG_7_ & ~n52842;
  assign n52845 = ~n52843 & ~n52844;
  assign n52846 = n43883 & ~n52845;
  assign n52847 = n43884 & ~n52845;
  assign n52848 = n51933 & ~n52840;
  assign n52849 = n51936 & ~n52840;
  assign n52850 = ~n52848 & ~n52849;
  assign n52851 = n43699 & ~n52845;
  assign n52852 = n52850 & ~n52851;
  assign n52853 = ~n52846 & ~n52847;
  assign n52854 = n52852 & n52853;
  assign n52855 = P1_P1_INSTADDRPOINTER_REG_6_ & ~n52762;
  assign n52856 = ~P1_P1_INSTADDRPOINTER_REG_6_ & n52762;
  assign n52857 = ~n52727 & ~n52856;
  assign n52858 = ~n52855 & ~n52857;
  assign n52859 = n52728 & ~n52759;
  assign n52860 = n52029 & n52859;
  assign n52861 = ~n52029 & ~n52859;
  assign n52862 = ~n52860 & ~n52861;
  assign n52863 = ~P1_P1_INSTADDRPOINTER_REG_7_ & ~n52862;
  assign n52864 = P1_P1_INSTADDRPOINTER_REG_7_ & n52862;
  assign n52865 = ~n52863 & ~n52864;
  assign n52866 = n52858 & ~n52865;
  assign n52867 = ~n52858 & n52865;
  assign n52868 = ~n52866 & ~n52867;
  assign n52869 = n52032 & ~n52868;
  assign n52870 = n52049 & ~n52840;
  assign n52871 = n52042 & ~n52840;
  assign n52872 = n52038 & ~n52840;
  assign n52873 = n43769 & ~n52840;
  assign n52874 = ~n52870 & ~n52871;
  assign n52875 = ~n52872 & n52874;
  assign n52876 = ~n52873 & n52875;
  assign n52877 = n43625 & ~n52845;
  assign n52878 = n43703 & ~n52845;
  assign n52879 = n43707 & ~n52845;
  assign n52880 = P1_P1_INSTADDRPOINTER_REG_6_ & n52780;
  assign n52881 = ~P1_P1_INSTADDRPOINTER_REG_7_ & n52880;
  assign n52882 = P1_P1_INSTADDRPOINTER_REG_7_ & ~n52880;
  assign n52883 = ~n52881 & ~n52882;
  assign n52884 = n43723 & ~n52883;
  assign n52885 = n43715 & ~n52883;
  assign n52886 = ~n52877 & ~n52878;
  assign n52887 = ~n52879 & n52886;
  assign n52888 = ~n52884 & n52887;
  assign n52889 = ~n52885 & n52888;
  assign n52890 = P1_P1_INSTADDRPOINTER_REG_6_ & ~n52799;
  assign n52891 = ~P1_P1_INSTADDRPOINTER_REG_6_ & n52799;
  assign n52892 = ~n52795 & ~n52891;
  assign n52893 = ~n52890 & ~n52892;
  assign n52894 = ~n52759 & n52796;
  assign n52895 = n52029 & n52894;
  assign n52896 = ~n52029 & ~n52894;
  assign n52897 = ~n52895 & ~n52896;
  assign n52898 = ~P1_P1_INSTADDRPOINTER_REG_7_ & ~n52897;
  assign n52899 = P1_P1_INSTADDRPOINTER_REG_7_ & n52897;
  assign n52900 = ~n52898 & ~n52899;
  assign n52901 = n52893 & ~n52900;
  assign n52902 = ~n52893 & n52900;
  assign n52903 = ~n52901 & ~n52902;
  assign n52904 = n43726 & ~n52903;
  assign n52905 = n43925 & ~n52840;
  assign n52906 = n43765 & ~n52840;
  assign n52907 = ~n52905 & ~n52906;
  assign n52908 = ~P1_P1_INSTADDRPOINTER_REG_6_ & ~n52817;
  assign n52909 = n52812 & ~n52908;
  assign n52910 = P1_P1_INSTADDRPOINTER_REG_5_ & ~n52908;
  assign n52911 = ~n52643 & n52910;
  assign n52912 = n52647 & ~n52908;
  assign n52913 = ~n52643 & n52912;
  assign n52914 = P1_P1_INSTADDRPOINTER_REG_6_ & n52817;
  assign n52915 = ~n52909 & ~n52911;
  assign n52916 = ~n52913 & n52915;
  assign n52917 = ~n52914 & n52916;
  assign n52918 = n52029 & ~n52815;
  assign n52919 = ~n52029 & ~n52759;
  assign n52920 = n52646 & n52919;
  assign n52921 = ~n52918 & ~n52920;
  assign n52922 = P1_P1_INSTADDRPOINTER_REG_7_ & ~n52921;
  assign n52923 = ~P1_P1_INSTADDRPOINTER_REG_7_ & n52921;
  assign n52924 = ~n52922 & ~n52923;
  assign n52925 = n52917 & ~n52924;
  assign n52926 = ~n52917 & n52924;
  assign n52927 = ~n52925 & ~n52926;
  assign n52928 = n52030 & ~n52927;
  assign n52929 = n52876 & n52889;
  assign n52930 = ~n52904 & n52929;
  assign n52931 = n52907 & n52930;
  assign n52932 = ~n52928 & n52931;
  assign n52933 = ~n52841 & n52854;
  assign n52934 = ~n52869 & n52933;
  assign n52935 = n52932 & n52934;
  assign n52936 = n51925 & ~n52935;
  assign n52937 = ~n52835 & ~n52836;
  assign n8831 = n52936 | ~n52937;
  assign n52939 = P1_P1_INSTADDRPOINTER_REG_8_ & n51924;
  assign n52940 = P1_P1_REIP_REG_8_ & n52069;
  assign n52941 = P1_P1_INSTADDRPOINTER_REG_7_ & n52837;
  assign n52942 = ~P1_P1_INSTADDRPOINTER_REG_8_ & n52941;
  assign n52943 = P1_P1_INSTADDRPOINTER_REG_8_ & ~n52941;
  assign n52944 = ~n52942 & ~n52943;
  assign n52945 = ~n43812 & ~n52944;
  assign n52946 = P1_P1_INSTADDRPOINTER_REG_7_ & n52842;
  assign n52947 = ~P1_P1_INSTADDRPOINTER_REG_8_ & n52946;
  assign n52948 = P1_P1_INSTADDRPOINTER_REG_8_ & ~n52946;
  assign n52949 = ~n52947 & ~n52948;
  assign n52950 = n43883 & ~n52949;
  assign n52951 = n43884 & ~n52949;
  assign n52952 = n51933 & ~n52944;
  assign n52953 = n51936 & ~n52944;
  assign n52954 = ~n52952 & ~n52953;
  assign n52955 = n43699 & ~n52949;
  assign n52956 = n52954 & ~n52955;
  assign n52957 = ~n52950 & ~n52951;
  assign n52958 = n52956 & n52957;
  assign n52959 = ~n52858 & ~n52862;
  assign n52960 = P1_P1_INSTADDRPOINTER_REG_7_ & ~n52858;
  assign n52961 = P1_P1_INSTADDRPOINTER_REG_7_ & ~n52862;
  assign n52962 = ~n52959 & ~n52960;
  assign n52963 = ~n52961 & n52962;
  assign n52964 = n52728 & n52919;
  assign n52965 = ~P1_P1_INSTADDRPOINTER_REG_8_ & n52964;
  assign n52966 = P1_P1_INSTADDRPOINTER_REG_8_ & ~n52964;
  assign n52967 = ~n52965 & ~n52966;
  assign n52968 = n52963 & ~n52967;
  assign n52969 = ~n52963 & n52967;
  assign n52970 = ~n52968 & ~n52969;
  assign n52971 = n52032 & ~n52970;
  assign n52972 = n52049 & ~n52944;
  assign n52973 = n52042 & ~n52944;
  assign n52974 = n52038 & ~n52944;
  assign n52975 = n43769 & ~n52944;
  assign n52976 = ~n52972 & ~n52973;
  assign n52977 = ~n52974 & n52976;
  assign n52978 = ~n52975 & n52977;
  assign n52979 = n43625 & ~n52949;
  assign n52980 = n43703 & ~n52949;
  assign n52981 = n43707 & ~n52949;
  assign n52982 = P1_P1_INSTADDRPOINTER_REG_7_ & n52880;
  assign n52983 = ~P1_P1_INSTADDRPOINTER_REG_8_ & n52982;
  assign n52984 = P1_P1_INSTADDRPOINTER_REG_8_ & ~n52982;
  assign n52985 = ~n52983 & ~n52984;
  assign n52986 = n43723 & ~n52985;
  assign n52987 = n43715 & ~n52985;
  assign n52988 = ~n52979 & ~n52980;
  assign n52989 = ~n52981 & n52988;
  assign n52990 = ~n52986 & n52989;
  assign n52991 = ~n52987 & n52990;
  assign n52992 = ~n52893 & ~n52897;
  assign n52993 = P1_P1_INSTADDRPOINTER_REG_7_ & ~n52893;
  assign n52994 = P1_P1_INSTADDRPOINTER_REG_7_ & ~n52897;
  assign n52995 = ~n52992 & ~n52993;
  assign n52996 = ~n52994 & n52995;
  assign n52997 = n52796 & n52919;
  assign n52998 = ~P1_P1_INSTADDRPOINTER_REG_8_ & n52997;
  assign n52999 = P1_P1_INSTADDRPOINTER_REG_8_ & ~n52997;
  assign n53000 = ~n52998 & ~n52999;
  assign n53001 = n52996 & ~n53000;
  assign n53002 = ~n52996 & n53000;
  assign n53003 = ~n53001 & ~n53002;
  assign n53004 = n43726 & ~n53003;
  assign n53005 = n43925 & ~n52944;
  assign n53006 = n43765 & ~n52944;
  assign n53007 = ~n53005 & ~n53006;
  assign n53008 = ~P1_P1_INSTADDRPOINTER_REG_7_ & ~n52921;
  assign n53009 = ~n52917 & ~n53008;
  assign n53010 = P1_P1_INSTADDRPOINTER_REG_7_ & n52921;
  assign n53011 = ~n53009 & ~n53010;
  assign n53012 = ~P1_P1_INSTADDRPOINTER_REG_8_ & ~n52920;
  assign n53013 = P1_P1_INSTADDRPOINTER_REG_8_ & n52920;
  assign n53014 = ~n53012 & ~n53013;
  assign n53015 = n53011 & ~n53014;
  assign n53016 = ~n53011 & n53014;
  assign n53017 = ~n53015 & ~n53016;
  assign n53018 = n52030 & ~n53017;
  assign n53019 = n52978 & n52991;
  assign n53020 = ~n53004 & n53019;
  assign n53021 = n53007 & n53020;
  assign n53022 = ~n53018 & n53021;
  assign n53023 = ~n52945 & n52958;
  assign n53024 = ~n52971 & n53023;
  assign n53025 = n53022 & n53024;
  assign n53026 = n51925 & ~n53025;
  assign n53027 = ~n52939 & ~n52940;
  assign n8836 = n53026 | ~n53027;
  assign n53029 = P1_P1_INSTADDRPOINTER_REG_9_ & n51924;
  assign n53030 = P1_P1_REIP_REG_9_ & n52069;
  assign n53031 = P1_P1_INSTADDRPOINTER_REG_8_ & n52941;
  assign n53032 = ~P1_P1_INSTADDRPOINTER_REG_9_ & n53031;
  assign n53033 = P1_P1_INSTADDRPOINTER_REG_9_ & ~n53031;
  assign n53034 = ~n53032 & ~n53033;
  assign n53035 = ~n43812 & ~n53034;
  assign n53036 = P1_P1_INSTADDRPOINTER_REG_8_ & n52946;
  assign n53037 = ~P1_P1_INSTADDRPOINTER_REG_9_ & n53036;
  assign n53038 = P1_P1_INSTADDRPOINTER_REG_9_ & ~n53036;
  assign n53039 = ~n53037 & ~n53038;
  assign n53040 = n43883 & ~n53039;
  assign n53041 = n43884 & ~n53039;
  assign n53042 = n51933 & ~n53034;
  assign n53043 = n51936 & ~n53034;
  assign n53044 = ~n53042 & ~n53043;
  assign n53045 = n43699 & ~n53039;
  assign n53046 = n53044 & ~n53045;
  assign n53047 = ~n53040 & ~n53041;
  assign n53048 = n53046 & n53047;
  assign n53049 = P1_P1_INSTADDRPOINTER_REG_8_ & n52964;
  assign n53050 = ~P1_P1_INSTADDRPOINTER_REG_8_ & ~n52964;
  assign n53051 = ~n52963 & ~n53050;
  assign n53052 = ~n53049 & ~n53051;
  assign n53053 = ~P1_P1_INSTADDRPOINTER_REG_9_ & n53052;
  assign n53054 = P1_P1_INSTADDRPOINTER_REG_9_ & ~n53052;
  assign n53055 = ~n53053 & ~n53054;
  assign n53056 = n52032 & n53055;
  assign n53057 = n52049 & ~n53034;
  assign n53058 = n52042 & ~n53034;
  assign n53059 = n52038 & ~n53034;
  assign n53060 = n43769 & ~n53034;
  assign n53061 = ~n53057 & ~n53058;
  assign n53062 = ~n53059 & n53061;
  assign n53063 = ~n53060 & n53062;
  assign n53064 = n43625 & ~n53039;
  assign n53065 = n43703 & ~n53039;
  assign n53066 = n43707 & ~n53039;
  assign n53067 = P1_P1_INSTADDRPOINTER_REG_8_ & n52982;
  assign n53068 = ~P1_P1_INSTADDRPOINTER_REG_9_ & n53067;
  assign n53069 = P1_P1_INSTADDRPOINTER_REG_9_ & ~n53067;
  assign n53070 = ~n53068 & ~n53069;
  assign n53071 = n43723 & ~n53070;
  assign n53072 = n43715 & ~n53070;
  assign n53073 = ~n53064 & ~n53065;
  assign n53074 = ~n53066 & n53073;
  assign n53075 = ~n53071 & n53074;
  assign n53076 = ~n53072 & n53075;
  assign n53077 = P1_P1_INSTADDRPOINTER_REG_8_ & n52997;
  assign n53078 = ~P1_P1_INSTADDRPOINTER_REG_8_ & ~n52997;
  assign n53079 = ~n52996 & ~n53078;
  assign n53080 = ~n53077 & ~n53079;
  assign n53081 = ~P1_P1_INSTADDRPOINTER_REG_9_ & n53080;
  assign n53082 = P1_P1_INSTADDRPOINTER_REG_9_ & ~n53080;
  assign n53083 = ~n53081 & ~n53082;
  assign n53084 = n43726 & n53083;
  assign n53085 = n53063 & n53076;
  assign n53086 = ~n53084 & n53085;
  assign n53087 = n43925 & ~n53034;
  assign n53088 = n43765 & ~n53034;
  assign n53089 = ~n53087 & ~n53088;
  assign n53090 = P1_P1_INSTADDRPOINTER_REG_8_ & ~n52920;
  assign n53091 = ~P1_P1_INSTADDRPOINTER_REG_8_ & n52920;
  assign n53092 = ~n53011 & ~n53091;
  assign n53093 = ~n53090 & ~n53092;
  assign n53094 = P1_P1_INSTADDRPOINTER_REG_9_ & n52920;
  assign n53095 = ~P1_P1_INSTADDRPOINTER_REG_9_ & ~n52920;
  assign n53096 = ~n53094 & ~n53095;
  assign n53097 = n53093 & ~n53096;
  assign n53098 = P1_P1_INSTADDRPOINTER_REG_9_ & ~n52920;
  assign n53099 = ~P1_P1_INSTADDRPOINTER_REG_9_ & n52920;
  assign n53100 = ~n53098 & ~n53099;
  assign n53101 = ~n53093 & ~n53100;
  assign n53102 = ~n53097 & ~n53101;
  assign n53103 = n52030 & ~n53102;
  assign n53104 = n53089 & ~n53103;
  assign n53105 = ~n53035 & n53048;
  assign n53106 = ~n53056 & n53105;
  assign n53107 = n53086 & n53106;
  assign n53108 = n53104 & n53107;
  assign n53109 = n51925 & ~n53108;
  assign n53110 = ~n53029 & ~n53030;
  assign n8841 = n53109 | ~n53110;
  assign n53112 = P1_P1_INSTADDRPOINTER_REG_10_ & n51924;
  assign n53113 = P1_P1_REIP_REG_10_ & n52069;
  assign n53114 = P1_P1_INSTADDRPOINTER_REG_9_ & n53031;
  assign n53115 = ~P1_P1_INSTADDRPOINTER_REG_10_ & n53114;
  assign n53116 = P1_P1_INSTADDRPOINTER_REG_10_ & ~n53114;
  assign n53117 = ~n53115 & ~n53116;
  assign n53118 = ~n43812 & ~n53117;
  assign n53119 = P1_P1_INSTADDRPOINTER_REG_9_ & n53036;
  assign n53120 = ~P1_P1_INSTADDRPOINTER_REG_10_ & n53119;
  assign n53121 = P1_P1_INSTADDRPOINTER_REG_10_ & ~n53119;
  assign n53122 = ~n53120 & ~n53121;
  assign n53123 = n43883 & ~n53122;
  assign n53124 = n43884 & ~n53122;
  assign n53125 = n51933 & ~n53117;
  assign n53126 = n51936 & ~n53117;
  assign n53127 = ~n53125 & ~n53126;
  assign n53128 = n43699 & ~n53122;
  assign n53129 = n53127 & ~n53128;
  assign n53130 = ~n53123 & ~n53124;
  assign n53131 = n53129 & n53130;
  assign n53132 = ~P1_P1_INSTADDRPOINTER_REG_10_ & ~n53054;
  assign n53133 = P1_P1_INSTADDRPOINTER_REG_9_ & P1_P1_INSTADDRPOINTER_REG_10_;
  assign n53134 = ~n53052 & n53133;
  assign n53135 = ~n53132 & ~n53134;
  assign n53136 = n52032 & n53135;
  assign n53137 = n52049 & ~n53117;
  assign n53138 = n52042 & ~n53117;
  assign n53139 = n52038 & ~n53117;
  assign n53140 = n43769 & ~n53117;
  assign n53141 = ~n53137 & ~n53138;
  assign n53142 = ~n53139 & n53141;
  assign n53143 = ~n53140 & n53142;
  assign n53144 = n43625 & ~n53122;
  assign n53145 = n43703 & ~n53122;
  assign n53146 = n43707 & ~n53122;
  assign n53147 = P1_P1_INSTADDRPOINTER_REG_9_ & n53067;
  assign n53148 = ~P1_P1_INSTADDRPOINTER_REG_10_ & n53147;
  assign n53149 = P1_P1_INSTADDRPOINTER_REG_10_ & ~n53147;
  assign n53150 = ~n53148 & ~n53149;
  assign n53151 = n43723 & ~n53150;
  assign n53152 = n43715 & ~n53150;
  assign n53153 = ~n53144 & ~n53145;
  assign n53154 = ~n53146 & n53153;
  assign n53155 = ~n53151 & n53154;
  assign n53156 = ~n53152 & n53155;
  assign n53157 = ~P1_P1_INSTADDRPOINTER_REG_10_ & ~n53082;
  assign n53158 = ~n53080 & n53133;
  assign n53159 = ~n53157 & ~n53158;
  assign n53160 = n43726 & n53159;
  assign n53161 = n53143 & n53156;
  assign n53162 = ~n53160 & n53161;
  assign n53163 = n43925 & ~n53117;
  assign n53164 = n43765 & ~n53117;
  assign n53165 = ~n53163 & ~n53164;
  assign n53166 = ~n53090 & ~n53098;
  assign n53167 = ~n53091 & ~n53099;
  assign n53168 = ~n53011 & n53167;
  assign n53169 = n53166 & ~n53168;
  assign n53170 = ~P1_P1_INSTADDRPOINTER_REG_10_ & ~n52920;
  assign n53171 = P1_P1_INSTADDRPOINTER_REG_10_ & n52920;
  assign n53172 = ~n53170 & ~n53171;
  assign n53173 = n53169 & ~n53172;
  assign n53174 = P1_P1_INSTADDRPOINTER_REG_10_ & ~n52920;
  assign n53175 = ~P1_P1_INSTADDRPOINTER_REG_10_ & n52920;
  assign n53176 = ~n53174 & ~n53175;
  assign n53177 = ~n53169 & ~n53176;
  assign n53178 = ~n53173 & ~n53177;
  assign n53179 = n52030 & ~n53178;
  assign n53180 = n53165 & ~n53179;
  assign n53181 = ~n53118 & n53131;
  assign n53182 = ~n53136 & n53181;
  assign n53183 = n53162 & n53182;
  assign n53184 = n53180 & n53183;
  assign n53185 = n51925 & ~n53184;
  assign n53186 = ~n53112 & ~n53113;
  assign n8846 = n53185 | ~n53186;
  assign n53188 = P1_P1_INSTADDRPOINTER_REG_11_ & n51924;
  assign n53189 = P1_P1_REIP_REG_11_ & n52069;
  assign n53190 = P1_P1_INSTADDRPOINTER_REG_10_ & n53114;
  assign n53191 = ~P1_P1_INSTADDRPOINTER_REG_11_ & n53190;
  assign n53192 = P1_P1_INSTADDRPOINTER_REG_11_ & ~n53190;
  assign n53193 = ~n53191 & ~n53192;
  assign n53194 = ~n43812 & ~n53193;
  assign n53195 = P1_P1_INSTADDRPOINTER_REG_10_ & n53119;
  assign n53196 = ~P1_P1_INSTADDRPOINTER_REG_11_ & n53195;
  assign n53197 = P1_P1_INSTADDRPOINTER_REG_11_ & ~n53195;
  assign n53198 = ~n53196 & ~n53197;
  assign n53199 = n43883 & ~n53198;
  assign n53200 = n43884 & ~n53198;
  assign n53201 = n51933 & ~n53193;
  assign n53202 = n51936 & ~n53193;
  assign n53203 = ~n53201 & ~n53202;
  assign n53204 = n43699 & ~n53198;
  assign n53205 = n53203 & ~n53204;
  assign n53206 = ~n53199 & ~n53200;
  assign n53207 = n53205 & n53206;
  assign n53208 = P1_P1_INSTADDRPOINTER_REG_11_ & ~n53134;
  assign n53209 = ~P1_P1_INSTADDRPOINTER_REG_11_ & n53134;
  assign n53210 = ~n53208 & ~n53209;
  assign n53211 = n52032 & ~n53210;
  assign n53212 = n52049 & ~n53193;
  assign n53213 = n52042 & ~n53193;
  assign n53214 = n52038 & ~n53193;
  assign n53215 = n43769 & ~n53193;
  assign n53216 = ~n53212 & ~n53213;
  assign n53217 = ~n53214 & n53216;
  assign n53218 = ~n53215 & n53217;
  assign n53219 = n43625 & ~n53198;
  assign n53220 = n43703 & ~n53198;
  assign n53221 = n43707 & ~n53198;
  assign n53222 = P1_P1_INSTADDRPOINTER_REG_10_ & n53147;
  assign n53223 = ~P1_P1_INSTADDRPOINTER_REG_11_ & n53222;
  assign n53224 = P1_P1_INSTADDRPOINTER_REG_11_ & ~n53222;
  assign n53225 = ~n53223 & ~n53224;
  assign n53226 = n43723 & ~n53225;
  assign n53227 = n43715 & ~n53225;
  assign n53228 = ~n53219 & ~n53220;
  assign n53229 = ~n53221 & n53228;
  assign n53230 = ~n53226 & n53229;
  assign n53231 = ~n53227 & n53230;
  assign n53232 = P1_P1_INSTADDRPOINTER_REG_11_ & ~n53158;
  assign n53233 = ~P1_P1_INSTADDRPOINTER_REG_11_ & n53158;
  assign n53234 = ~n53232 & ~n53233;
  assign n53235 = n43726 & ~n53234;
  assign n53236 = n53218 & n53231;
  assign n53237 = ~n53235 & n53236;
  assign n53238 = n43925 & ~n53193;
  assign n53239 = n43765 & ~n53193;
  assign n53240 = ~n53238 & ~n53239;
  assign n53241 = n53166 & ~n53174;
  assign n53242 = n53167 & ~n53175;
  assign n53243 = ~n53011 & n53242;
  assign n53244 = n53241 & ~n53243;
  assign n53245 = ~P1_P1_INSTADDRPOINTER_REG_11_ & ~n52920;
  assign n53246 = P1_P1_INSTADDRPOINTER_REG_11_ & n52920;
  assign n53247 = ~n53245 & ~n53246;
  assign n53248 = n53244 & ~n53247;
  assign n53249 = ~n53244 & n53247;
  assign n53250 = ~n53248 & ~n53249;
  assign n53251 = n52030 & ~n53250;
  assign n53252 = n53240 & ~n53251;
  assign n53253 = ~n53194 & n53207;
  assign n53254 = ~n53211 & n53253;
  assign n53255 = n53237 & n53254;
  assign n53256 = n53252 & n53255;
  assign n53257 = n51925 & ~n53256;
  assign n53258 = ~n53188 & ~n53189;
  assign n8851 = n53257 | ~n53258;
  assign n53260 = P1_P1_INSTADDRPOINTER_REG_12_ & n51924;
  assign n53261 = P1_P1_REIP_REG_12_ & n52069;
  assign n53262 = P1_P1_INSTADDRPOINTER_REG_11_ & n53190;
  assign n53263 = ~P1_P1_INSTADDRPOINTER_REG_12_ & n53262;
  assign n53264 = P1_P1_INSTADDRPOINTER_REG_12_ & ~n53262;
  assign n53265 = ~n53263 & ~n53264;
  assign n53266 = ~n43812 & ~n53265;
  assign n53267 = P1_P1_INSTADDRPOINTER_REG_11_ & n53195;
  assign n53268 = ~P1_P1_INSTADDRPOINTER_REG_12_ & n53267;
  assign n53269 = P1_P1_INSTADDRPOINTER_REG_12_ & ~n53267;
  assign n53270 = ~n53268 & ~n53269;
  assign n53271 = n43883 & ~n53270;
  assign n53272 = n43884 & ~n53270;
  assign n53273 = n51933 & ~n53265;
  assign n53274 = n51936 & ~n53265;
  assign n53275 = ~n53273 & ~n53274;
  assign n53276 = n43699 & ~n53270;
  assign n53277 = n53275 & ~n53276;
  assign n53278 = ~n53271 & ~n53272;
  assign n53279 = n53277 & n53278;
  assign n53280 = P1_P1_INSTADDRPOINTER_REG_11_ & n53134;
  assign n53281 = ~P1_P1_INSTADDRPOINTER_REG_12_ & ~n53280;
  assign n53282 = P1_P1_INSTADDRPOINTER_REG_12_ & n53133;
  assign n53283 = P1_P1_INSTADDRPOINTER_REG_11_ & n53282;
  assign n53284 = ~n53052 & n53283;
  assign n53285 = ~n53281 & ~n53284;
  assign n53286 = n52032 & n53285;
  assign n53287 = n52049 & ~n53265;
  assign n53288 = n52042 & ~n53265;
  assign n53289 = n52038 & ~n53265;
  assign n53290 = n43769 & ~n53265;
  assign n53291 = ~n53287 & ~n53288;
  assign n53292 = ~n53289 & n53291;
  assign n53293 = ~n53290 & n53292;
  assign n53294 = n43625 & ~n53270;
  assign n53295 = n43703 & ~n53270;
  assign n53296 = n43707 & ~n53270;
  assign n53297 = P1_P1_INSTADDRPOINTER_REG_11_ & n53222;
  assign n53298 = ~P1_P1_INSTADDRPOINTER_REG_12_ & n53297;
  assign n53299 = P1_P1_INSTADDRPOINTER_REG_12_ & ~n53297;
  assign n53300 = ~n53298 & ~n53299;
  assign n53301 = n43723 & ~n53300;
  assign n53302 = n43715 & ~n53300;
  assign n53303 = ~n53294 & ~n53295;
  assign n53304 = ~n53296 & n53303;
  assign n53305 = ~n53301 & n53304;
  assign n53306 = ~n53302 & n53305;
  assign n53307 = P1_P1_INSTADDRPOINTER_REG_11_ & n53158;
  assign n53308 = ~P1_P1_INSTADDRPOINTER_REG_12_ & ~n53307;
  assign n53309 = ~n53080 & n53283;
  assign n53310 = ~n53308 & ~n53309;
  assign n53311 = n43726 & n53310;
  assign n53312 = n53293 & n53306;
  assign n53313 = ~n53311 & n53312;
  assign n53314 = n43925 & ~n53265;
  assign n53315 = n43765 & ~n53265;
  assign n53316 = ~n53314 & ~n53315;
  assign n53317 = ~P1_P1_INSTADDRPOINTER_REG_12_ & ~n52920;
  assign n53318 = P1_P1_INSTADDRPOINTER_REG_12_ & n52920;
  assign n53319 = ~n53317 & ~n53318;
  assign n53320 = ~P1_P1_INSTADDRPOINTER_REG_11_ & n52920;
  assign n53321 = ~n53244 & ~n53320;
  assign n53322 = P1_P1_INSTADDRPOINTER_REG_11_ & ~n52920;
  assign n53323 = ~n53321 & ~n53322;
  assign n53324 = ~n53319 & n53323;
  assign n53325 = ~P1_P1_INSTADDRPOINTER_REG_12_ & n52920;
  assign n53326 = P1_P1_INSTADDRPOINTER_REG_12_ & ~n52920;
  assign n53327 = ~n53325 & ~n53326;
  assign n53328 = ~n53323 & ~n53327;
  assign n53329 = ~n53324 & ~n53328;
  assign n53330 = n52030 & ~n53329;
  assign n53331 = n53316 & ~n53330;
  assign n53332 = ~n53266 & n53279;
  assign n53333 = ~n53286 & n53332;
  assign n53334 = n53313 & n53333;
  assign n53335 = n53331 & n53334;
  assign n53336 = n51925 & ~n53335;
  assign n53337 = ~n53260 & ~n53261;
  assign n8856 = n53336 | ~n53337;
  assign n53339 = P1_P1_INSTADDRPOINTER_REG_13_ & n51924;
  assign n53340 = P1_P1_REIP_REG_13_ & n52069;
  assign n53341 = P1_P1_INSTADDRPOINTER_REG_12_ & n53262;
  assign n53342 = ~P1_P1_INSTADDRPOINTER_REG_13_ & n53341;
  assign n53343 = P1_P1_INSTADDRPOINTER_REG_13_ & ~n53341;
  assign n53344 = ~n53342 & ~n53343;
  assign n53345 = ~n43812 & ~n53344;
  assign n53346 = n43925 & ~n53344;
  assign n53347 = n43765 & ~n53344;
  assign n53348 = ~n53346 & ~n53347;
  assign n53349 = ~P1_P1_INSTADDRPOINTER_REG_13_ & ~n53284;
  assign n53350 = P1_P1_INSTADDRPOINTER_REG_13_ & n53284;
  assign n53351 = ~n53349 & ~n53350;
  assign n53352 = n52032 & n53351;
  assign n53353 = n52049 & ~n53344;
  assign n53354 = n43769 & ~n53344;
  assign n53355 = n52038 & ~n53344;
  assign n53356 = n52042 & ~n53344;
  assign n53357 = ~n53353 & ~n53354;
  assign n53358 = ~n53355 & n53357;
  assign n53359 = ~n53356 & n53358;
  assign n53360 = P1_P1_INSTADDRPOINTER_REG_12_ & n53267;
  assign n53361 = ~P1_P1_INSTADDRPOINTER_REG_13_ & n53360;
  assign n53362 = P1_P1_INSTADDRPOINTER_REG_13_ & ~n53360;
  assign n53363 = ~n53361 & ~n53362;
  assign n53364 = n43625 & ~n53363;
  assign n53365 = n43703 & ~n53363;
  assign n53366 = n43707 & ~n53363;
  assign n53367 = P1_P1_INSTADDRPOINTER_REG_12_ & n53297;
  assign n53368 = ~P1_P1_INSTADDRPOINTER_REG_13_ & n53367;
  assign n53369 = P1_P1_INSTADDRPOINTER_REG_13_ & ~n53367;
  assign n53370 = ~n53368 & ~n53369;
  assign n53371 = n43723 & ~n53370;
  assign n53372 = n43715 & ~n53370;
  assign n53373 = ~n53364 & ~n53365;
  assign n53374 = ~n53366 & n53373;
  assign n53375 = ~n53371 & n53374;
  assign n53376 = ~n53372 & n53375;
  assign n53377 = ~P1_P1_INSTADDRPOINTER_REG_13_ & ~n53309;
  assign n53378 = P1_P1_INSTADDRPOINTER_REG_13_ & n53309;
  assign n53379 = ~n53377 & ~n53378;
  assign n53380 = n43726 & n53379;
  assign n53381 = n53359 & n53376;
  assign n53382 = ~n53380 & n53381;
  assign n53383 = n43883 & ~n53363;
  assign n53384 = n43884 & ~n53363;
  assign n53385 = n43699 & ~n53363;
  assign n53386 = n51936 & ~n53344;
  assign n53387 = n51933 & ~n53344;
  assign n53388 = ~n53385 & ~n53386;
  assign n53389 = ~n53387 & n53388;
  assign n53390 = P1_P1_INSTADDRPOINTER_REG_13_ & ~n52920;
  assign n53391 = P1_P1_INSTADDRPOINTER_REG_12_ & P1_P1_INSTADDRPOINTER_REG_13_;
  assign n53392 = n52920 & ~n53391;
  assign n53393 = ~n53390 & ~n53392;
  assign n53394 = n53323 & ~n53326;
  assign n53395 = n53393 & ~n53394;
  assign n53396 = ~P1_P1_INSTADDRPOINTER_REG_13_ & ~n52920;
  assign n53397 = P1_P1_INSTADDRPOINTER_REG_13_ & n52920;
  assign n53398 = ~n53396 & ~n53397;
  assign n53399 = ~n53326 & n53398;
  assign n53400 = ~n53323 & ~n53325;
  assign n53401 = n53399 & ~n53400;
  assign n53402 = ~n53395 & ~n53401;
  assign n53403 = n52030 & n53402;
  assign n53404 = ~n53383 & ~n53384;
  assign n53405 = n53389 & n53404;
  assign n53406 = ~n53403 & n53405;
  assign n53407 = ~n53345 & n53348;
  assign n53408 = ~n53352 & n53407;
  assign n53409 = n53382 & n53408;
  assign n53410 = n53406 & n53409;
  assign n53411 = n51925 & ~n53410;
  assign n53412 = ~n53339 & ~n53340;
  assign n8861 = n53411 | ~n53412;
  assign n53414 = P1_P1_INSTADDRPOINTER_REG_14_ & n51924;
  assign n53415 = P1_P1_REIP_REG_14_ & n52069;
  assign n53416 = P1_P1_INSTADDRPOINTER_REG_13_ & n53341;
  assign n53417 = ~P1_P1_INSTADDRPOINTER_REG_14_ & n53416;
  assign n53418 = P1_P1_INSTADDRPOINTER_REG_14_ & ~n53416;
  assign n53419 = ~n53417 & ~n53418;
  assign n53420 = ~n43812 & ~n53419;
  assign n53421 = P1_P1_INSTADDRPOINTER_REG_13_ & n53360;
  assign n53422 = ~P1_P1_INSTADDRPOINTER_REG_14_ & n53421;
  assign n53423 = P1_P1_INSTADDRPOINTER_REG_14_ & ~n53421;
  assign n53424 = ~n53422 & ~n53423;
  assign n53425 = n43883 & ~n53424;
  assign n53426 = n43884 & ~n53424;
  assign n53427 = n43699 & ~n53424;
  assign n53428 = n51936 & ~n53419;
  assign n53429 = n51933 & ~n53419;
  assign n53430 = ~n53427 & ~n53428;
  assign n53431 = ~n53429 & n53430;
  assign n53432 = ~n53425 & ~n53426;
  assign n53433 = n53431 & n53432;
  assign n53434 = ~P1_P1_INSTADDRPOINTER_REG_14_ & n53350;
  assign n53435 = P1_P1_INSTADDRPOINTER_REG_14_ & ~n53350;
  assign n53436 = ~n53434 & ~n53435;
  assign n53437 = n52032 & ~n53436;
  assign n53438 = n52049 & ~n53419;
  assign n53439 = n43769 & ~n53419;
  assign n53440 = n52038 & ~n53419;
  assign n53441 = n52042 & ~n53419;
  assign n53442 = ~n53438 & ~n53439;
  assign n53443 = ~n53440 & n53442;
  assign n53444 = ~n53441 & n53443;
  assign n53445 = n43625 & ~n53424;
  assign n53446 = n43703 & ~n53424;
  assign n53447 = n43707 & ~n53424;
  assign n53448 = P1_P1_INSTADDRPOINTER_REG_13_ & n53367;
  assign n53449 = ~P1_P1_INSTADDRPOINTER_REG_14_ & n53448;
  assign n53450 = P1_P1_INSTADDRPOINTER_REG_14_ & ~n53448;
  assign n53451 = ~n53449 & ~n53450;
  assign n53452 = n43723 & ~n53451;
  assign n53453 = n43715 & ~n53451;
  assign n53454 = ~n53445 & ~n53446;
  assign n53455 = ~n53447 & n53454;
  assign n53456 = ~n53452 & n53455;
  assign n53457 = ~n53453 & n53456;
  assign n53458 = ~P1_P1_INSTADDRPOINTER_REG_14_ & n53378;
  assign n53459 = P1_P1_INSTADDRPOINTER_REG_14_ & ~n53378;
  assign n53460 = ~n53458 & ~n53459;
  assign n53461 = n43726 & ~n53460;
  assign n53462 = n53444 & n53457;
  assign n53463 = ~n53461 & n53462;
  assign n53464 = n43925 & ~n53419;
  assign n53465 = n43765 & ~n53419;
  assign n53466 = ~n53464 & ~n53465;
  assign n53467 = ~n53320 & ~n53392;
  assign n53468 = ~n53244 & n53467;
  assign n53469 = ~n53326 & ~n53390;
  assign n53470 = ~n53322 & n53469;
  assign n53471 = ~n53468 & n53470;
  assign n53472 = ~P1_P1_INSTADDRPOINTER_REG_14_ & ~n52920;
  assign n53473 = P1_P1_INSTADDRPOINTER_REG_14_ & n52920;
  assign n53474 = ~n53472 & ~n53473;
  assign n53475 = n53471 & ~n53474;
  assign n53476 = ~n53471 & n53474;
  assign n53477 = ~n53475 & ~n53476;
  assign n53478 = n52030 & ~n53477;
  assign n53479 = n53466 & ~n53478;
  assign n53480 = ~n53420 & n53433;
  assign n53481 = ~n53437 & n53480;
  assign n53482 = n53463 & n53481;
  assign n53483 = n53479 & n53482;
  assign n53484 = n51925 & ~n53483;
  assign n53485 = ~n53414 & ~n53415;
  assign n8866 = n53484 | ~n53485;
  assign n53487 = P1_P1_INSTADDRPOINTER_REG_15_ & n51924;
  assign n53488 = P1_P1_REIP_REG_15_ & n52069;
  assign n53489 = P1_P1_INSTADDRPOINTER_REG_14_ & n53416;
  assign n53490 = ~P1_P1_INSTADDRPOINTER_REG_15_ & n53489;
  assign n53491 = P1_P1_INSTADDRPOINTER_REG_15_ & ~n53489;
  assign n53492 = ~n53490 & ~n53491;
  assign n53493 = ~n43812 & ~n53492;
  assign n53494 = n43925 & ~n53492;
  assign n53495 = n43765 & ~n53492;
  assign n53496 = ~n53494 & ~n53495;
  assign n53497 = P1_P1_INSTADDRPOINTER_REG_14_ & n53350;
  assign n53498 = ~P1_P1_INSTADDRPOINTER_REG_15_ & ~n53497;
  assign n53499 = P1_P1_INSTADDRPOINTER_REG_14_ & P1_P1_INSTADDRPOINTER_REG_15_;
  assign n53500 = P1_P1_INSTADDRPOINTER_REG_13_ & n53499;
  assign n53501 = n53284 & n53500;
  assign n53502 = ~n53498 & ~n53501;
  assign n53503 = n52032 & n53502;
  assign n53504 = n52049 & ~n53492;
  assign n53505 = n43769 & ~n53492;
  assign n53506 = n52038 & ~n53492;
  assign n53507 = n52042 & ~n53492;
  assign n53508 = ~n53504 & ~n53505;
  assign n53509 = ~n53506 & n53508;
  assign n53510 = ~n53507 & n53509;
  assign n53511 = P1_P1_INSTADDRPOINTER_REG_14_ & n53421;
  assign n53512 = ~P1_P1_INSTADDRPOINTER_REG_15_ & n53511;
  assign n53513 = P1_P1_INSTADDRPOINTER_REG_15_ & ~n53511;
  assign n53514 = ~n53512 & ~n53513;
  assign n53515 = n43625 & ~n53514;
  assign n53516 = n43703 & ~n53514;
  assign n53517 = n43707 & ~n53514;
  assign n53518 = P1_P1_INSTADDRPOINTER_REG_14_ & n53448;
  assign n53519 = ~P1_P1_INSTADDRPOINTER_REG_15_ & n53518;
  assign n53520 = P1_P1_INSTADDRPOINTER_REG_15_ & ~n53518;
  assign n53521 = ~n53519 & ~n53520;
  assign n53522 = n43723 & ~n53521;
  assign n53523 = n43715 & ~n53521;
  assign n53524 = ~n53515 & ~n53516;
  assign n53525 = ~n53517 & n53524;
  assign n53526 = ~n53522 & n53525;
  assign n53527 = ~n53523 & n53526;
  assign n53528 = P1_P1_INSTADDRPOINTER_REG_14_ & n53378;
  assign n53529 = ~P1_P1_INSTADDRPOINTER_REG_15_ & ~n53528;
  assign n53530 = n53309 & n53500;
  assign n53531 = ~n53529 & ~n53530;
  assign n53532 = n43726 & n53531;
  assign n53533 = n53510 & n53527;
  assign n53534 = ~n53532 & n53533;
  assign n53535 = n43883 & ~n53514;
  assign n53536 = n43884 & ~n53514;
  assign n53537 = n51933 & ~n53492;
  assign n53538 = n43699 & ~n53514;
  assign n53539 = n51936 & ~n53492;
  assign n53540 = ~n53538 & ~n53539;
  assign n53541 = P1_P1_INSTADDRPOINTER_REG_14_ & ~n52920;
  assign n53542 = n53470 & ~n53541;
  assign n53543 = ~P1_P1_INSTADDRPOINTER_REG_14_ & n52920;
  assign n53544 = n53467 & ~n53543;
  assign n53545 = ~n53244 & n53544;
  assign n53546 = n53542 & ~n53545;
  assign n53547 = ~P1_P1_INSTADDRPOINTER_REG_15_ & ~n52920;
  assign n53548 = P1_P1_INSTADDRPOINTER_REG_15_ & n52920;
  assign n53549 = ~n53547 & ~n53548;
  assign n53550 = n53546 & ~n53549;
  assign n53551 = ~n53546 & n53549;
  assign n53552 = ~n53550 & ~n53551;
  assign n53553 = n52030 & ~n53552;
  assign n53554 = ~n53535 & ~n53536;
  assign n53555 = ~n53537 & n53554;
  assign n53556 = n53540 & n53555;
  assign n53557 = ~n53553 & n53556;
  assign n53558 = ~n53493 & n53496;
  assign n53559 = ~n53503 & n53558;
  assign n53560 = n53534 & n53559;
  assign n53561 = n53557 & n53560;
  assign n53562 = n51925 & ~n53561;
  assign n53563 = ~n53487 & ~n53488;
  assign n8871 = n53562 | ~n53563;
  assign n53565 = P1_P1_INSTADDRPOINTER_REG_16_ & n51924;
  assign n53566 = P1_P1_REIP_REG_16_ & n52069;
  assign n53567 = P1_P1_INSTADDRPOINTER_REG_15_ & n53489;
  assign n53568 = ~P1_P1_INSTADDRPOINTER_REG_16_ & n53567;
  assign n53569 = P1_P1_INSTADDRPOINTER_REG_16_ & ~n53567;
  assign n53570 = ~n53568 & ~n53569;
  assign n53571 = ~n43812 & ~n53570;
  assign n53572 = n43925 & ~n53570;
  assign n53573 = n43765 & ~n53570;
  assign n53574 = ~n53572 & ~n53573;
  assign n53575 = ~P1_P1_INSTADDRPOINTER_REG_16_ & n53501;
  assign n53576 = P1_P1_INSTADDRPOINTER_REG_16_ & ~n53501;
  assign n53577 = ~n53575 & ~n53576;
  assign n53578 = n52032 & ~n53577;
  assign n53579 = n52049 & ~n53570;
  assign n53580 = n43769 & ~n53570;
  assign n53581 = n52038 & ~n53570;
  assign n53582 = n52042 & ~n53570;
  assign n53583 = ~n53579 & ~n53580;
  assign n53584 = ~n53581 & n53583;
  assign n53585 = ~n53582 & n53584;
  assign n53586 = P1_P1_INSTADDRPOINTER_REG_15_ & n53511;
  assign n53587 = ~P1_P1_INSTADDRPOINTER_REG_16_ & n53586;
  assign n53588 = P1_P1_INSTADDRPOINTER_REG_16_ & ~n53586;
  assign n53589 = ~n53587 & ~n53588;
  assign n53590 = n43625 & ~n53589;
  assign n53591 = n43703 & ~n53589;
  assign n53592 = n43707 & ~n53589;
  assign n53593 = P1_P1_INSTADDRPOINTER_REG_15_ & n53518;
  assign n53594 = ~P1_P1_INSTADDRPOINTER_REG_16_ & n53593;
  assign n53595 = P1_P1_INSTADDRPOINTER_REG_16_ & ~n53593;
  assign n53596 = ~n53594 & ~n53595;
  assign n53597 = n43723 & ~n53596;
  assign n53598 = n43715 & ~n53596;
  assign n53599 = ~n53590 & ~n53591;
  assign n53600 = ~n53592 & n53599;
  assign n53601 = ~n53597 & n53600;
  assign n53602 = ~n53598 & n53601;
  assign n53603 = ~P1_P1_INSTADDRPOINTER_REG_16_ & n53530;
  assign n53604 = P1_P1_INSTADDRPOINTER_REG_16_ & ~n53530;
  assign n53605 = ~n53603 & ~n53604;
  assign n53606 = n43726 & ~n53605;
  assign n53607 = n53585 & n53602;
  assign n53608 = ~n53606 & n53607;
  assign n53609 = n43883 & ~n53589;
  assign n53610 = n43884 & ~n53589;
  assign n53611 = n51933 & ~n53570;
  assign n53612 = n43699 & ~n53589;
  assign n53613 = n51936 & ~n53570;
  assign n53614 = ~n53612 & ~n53613;
  assign n53615 = P1_P1_INSTADDRPOINTER_REG_15_ & ~n52920;
  assign n53616 = ~P1_P1_INSTADDRPOINTER_REG_15_ & n52920;
  assign n53617 = ~n53546 & ~n53616;
  assign n53618 = ~n53615 & ~n53617;
  assign n53619 = ~P1_P1_INSTADDRPOINTER_REG_16_ & ~n52920;
  assign n53620 = P1_P1_INSTADDRPOINTER_REG_16_ & n52920;
  assign n53621 = ~n53619 & ~n53620;
  assign n53622 = n53618 & ~n53621;
  assign n53623 = ~n53618 & n53621;
  assign n53624 = ~n53622 & ~n53623;
  assign n53625 = n52030 & ~n53624;
  assign n53626 = ~n53609 & ~n53610;
  assign n53627 = ~n53611 & n53626;
  assign n53628 = n53614 & n53627;
  assign n53629 = ~n53625 & n53628;
  assign n53630 = ~n53571 & n53574;
  assign n53631 = ~n53578 & n53630;
  assign n53632 = n53608 & n53631;
  assign n53633 = n53629 & n53632;
  assign n53634 = n51925 & ~n53633;
  assign n53635 = ~n53565 & ~n53566;
  assign n8876 = n53634 | ~n53635;
  assign n53637 = P1_P1_INSTADDRPOINTER_REG_17_ & n51924;
  assign n53638 = P1_P1_REIP_REG_17_ & n52069;
  assign n53639 = P1_P1_INSTADDRPOINTER_REG_16_ & n53567;
  assign n53640 = ~P1_P1_INSTADDRPOINTER_REG_17_ & n53639;
  assign n53641 = P1_P1_INSTADDRPOINTER_REG_17_ & ~n53639;
  assign n53642 = ~n53640 & ~n53641;
  assign n53643 = ~n43812 & ~n53642;
  assign n53644 = n43925 & ~n53642;
  assign n53645 = n43765 & ~n53642;
  assign n53646 = ~n53644 & ~n53645;
  assign n53647 = P1_P1_INSTADDRPOINTER_REG_16_ & n53501;
  assign n53648 = ~P1_P1_INSTADDRPOINTER_REG_17_ & ~n53647;
  assign n53649 = P1_P1_INSTADDRPOINTER_REG_16_ & P1_P1_INSTADDRPOINTER_REG_17_;
  assign n53650 = n53501 & n53649;
  assign n53651 = ~n53648 & ~n53650;
  assign n53652 = n52032 & n53651;
  assign n53653 = n52049 & ~n53642;
  assign n53654 = n43769 & ~n53642;
  assign n53655 = n52038 & ~n53642;
  assign n53656 = n52042 & ~n53642;
  assign n53657 = ~n53653 & ~n53654;
  assign n53658 = ~n53655 & n53657;
  assign n53659 = ~n53656 & n53658;
  assign n53660 = P1_P1_INSTADDRPOINTER_REG_16_ & n53586;
  assign n53661 = ~P1_P1_INSTADDRPOINTER_REG_17_ & n53660;
  assign n53662 = P1_P1_INSTADDRPOINTER_REG_17_ & ~n53660;
  assign n53663 = ~n53661 & ~n53662;
  assign n53664 = n43625 & ~n53663;
  assign n53665 = n43703 & ~n53663;
  assign n53666 = n43707 & ~n53663;
  assign n53667 = P1_P1_INSTADDRPOINTER_REG_16_ & n53593;
  assign n53668 = ~P1_P1_INSTADDRPOINTER_REG_17_ & n53667;
  assign n53669 = P1_P1_INSTADDRPOINTER_REG_17_ & ~n53667;
  assign n53670 = ~n53668 & ~n53669;
  assign n53671 = n43723 & ~n53670;
  assign n53672 = n43715 & ~n53670;
  assign n53673 = ~n53664 & ~n53665;
  assign n53674 = ~n53666 & n53673;
  assign n53675 = ~n53671 & n53674;
  assign n53676 = ~n53672 & n53675;
  assign n53677 = P1_P1_INSTADDRPOINTER_REG_16_ & n53530;
  assign n53678 = ~P1_P1_INSTADDRPOINTER_REG_17_ & ~n53677;
  assign n53679 = n53530 & n53649;
  assign n53680 = ~n53678 & ~n53679;
  assign n53681 = n43726 & n53680;
  assign n53682 = n53659 & n53676;
  assign n53683 = ~n53681 & n53682;
  assign n53684 = n43883 & ~n53663;
  assign n53685 = n43884 & ~n53663;
  assign n53686 = n51933 & ~n53642;
  assign n53687 = n43699 & ~n53663;
  assign n53688 = n51936 & ~n53642;
  assign n53689 = ~n53687 & ~n53688;
  assign n53690 = ~n53618 & n53649;
  assign n53691 = n52920 & ~n53690;
  assign n53692 = P1_P1_INSTADDRPOINTER_REG_17_ & ~n52920;
  assign n53693 = ~P1_P1_INSTADDRPOINTER_REG_16_ & ~n53615;
  assign n53694 = ~n53617 & n53693;
  assign n53695 = ~n53691 & ~n53692;
  assign n53696 = ~n53694 & n53695;
  assign n53697 = P1_P1_INSTADDRPOINTER_REG_17_ & n53694;
  assign n53698 = ~n52920 & ~n53697;
  assign n53699 = P1_P1_INSTADDRPOINTER_REG_17_ & n52920;
  assign n53700 = P1_P1_INSTADDRPOINTER_REG_16_ & ~n53618;
  assign n53701 = ~n53698 & ~n53699;
  assign n53702 = ~n53700 & n53701;
  assign n53703 = ~n53696 & ~n53702;
  assign n53704 = n52030 & n53703;
  assign n53705 = ~n53684 & ~n53685;
  assign n53706 = ~n53686 & n53705;
  assign n53707 = n53689 & n53706;
  assign n53708 = ~n53704 & n53707;
  assign n53709 = ~n53643 & n53646;
  assign n53710 = ~n53652 & n53709;
  assign n53711 = n53683 & n53710;
  assign n53712 = n53708 & n53711;
  assign n53713 = n51925 & ~n53712;
  assign n53714 = ~n53637 & ~n53638;
  assign n8881 = n53713 | ~n53714;
  assign n53716 = P1_P1_INSTADDRPOINTER_REG_18_ & n51924;
  assign n53717 = P1_P1_REIP_REG_18_ & n52069;
  assign n53718 = P1_P1_INSTADDRPOINTER_REG_17_ & n53639;
  assign n53719 = ~P1_P1_INSTADDRPOINTER_REG_18_ & n53718;
  assign n53720 = P1_P1_INSTADDRPOINTER_REG_18_ & ~n53718;
  assign n53721 = ~n53719 & ~n53720;
  assign n53722 = ~n43812 & ~n53721;
  assign n53723 = n43925 & ~n53721;
  assign n53724 = n43765 & ~n53721;
  assign n53725 = ~n53723 & ~n53724;
  assign n53726 = ~P1_P1_INSTADDRPOINTER_REG_18_ & n53650;
  assign n53727 = P1_P1_INSTADDRPOINTER_REG_18_ & ~n53650;
  assign n53728 = ~n53726 & ~n53727;
  assign n53729 = n52032 & ~n53728;
  assign n53730 = n52049 & ~n53721;
  assign n53731 = n43769 & ~n53721;
  assign n53732 = n52038 & ~n53721;
  assign n53733 = n52042 & ~n53721;
  assign n53734 = ~n53730 & ~n53731;
  assign n53735 = ~n53732 & n53734;
  assign n53736 = ~n53733 & n53735;
  assign n53737 = P1_P1_INSTADDRPOINTER_REG_17_ & n53660;
  assign n53738 = ~P1_P1_INSTADDRPOINTER_REG_18_ & n53737;
  assign n53739 = P1_P1_INSTADDRPOINTER_REG_18_ & ~n53737;
  assign n53740 = ~n53738 & ~n53739;
  assign n53741 = n43625 & ~n53740;
  assign n53742 = n43703 & ~n53740;
  assign n53743 = n43707 & ~n53740;
  assign n53744 = P1_P1_INSTADDRPOINTER_REG_17_ & n53667;
  assign n53745 = ~P1_P1_INSTADDRPOINTER_REG_18_ & n53744;
  assign n53746 = P1_P1_INSTADDRPOINTER_REG_18_ & ~n53744;
  assign n53747 = ~n53745 & ~n53746;
  assign n53748 = n43723 & ~n53747;
  assign n53749 = n43715 & ~n53747;
  assign n53750 = ~n53741 & ~n53742;
  assign n53751 = ~n53743 & n53750;
  assign n53752 = ~n53748 & n53751;
  assign n53753 = ~n53749 & n53752;
  assign n53754 = ~P1_P1_INSTADDRPOINTER_REG_18_ & n53679;
  assign n53755 = P1_P1_INSTADDRPOINTER_REG_18_ & ~n53679;
  assign n53756 = ~n53754 & ~n53755;
  assign n53757 = n43726 & ~n53756;
  assign n53758 = n53736 & n53753;
  assign n53759 = ~n53757 & n53758;
  assign n53760 = n43883 & ~n53740;
  assign n53761 = n43884 & ~n53740;
  assign n53762 = n51933 & ~n53721;
  assign n53763 = n43699 & ~n53740;
  assign n53764 = n51936 & ~n53721;
  assign n53765 = ~n53763 & ~n53764;
  assign n53766 = ~n52920 & ~n53694;
  assign n53767 = ~n53690 & ~n53766;
  assign n53768 = ~n53692 & n53767;
  assign n53769 = ~P1_P1_INSTADDRPOINTER_REG_18_ & ~n52920;
  assign n53770 = P1_P1_INSTADDRPOINTER_REG_18_ & n52920;
  assign n53771 = ~n53769 & ~n53770;
  assign n53772 = n53768 & ~n53771;
  assign n53773 = ~n53768 & n53771;
  assign n53774 = ~n53772 & ~n53773;
  assign n53775 = n52030 & ~n53774;
  assign n53776 = ~n53760 & ~n53761;
  assign n53777 = ~n53762 & n53776;
  assign n53778 = n53765 & n53777;
  assign n53779 = ~n53775 & n53778;
  assign n53780 = ~n53722 & n53725;
  assign n53781 = ~n53729 & n53780;
  assign n53782 = n53759 & n53781;
  assign n53783 = n53779 & n53782;
  assign n53784 = n51925 & ~n53783;
  assign n53785 = ~n53716 & ~n53717;
  assign n8886 = n53784 | ~n53785;
  assign n53787 = P1_P1_INSTADDRPOINTER_REG_19_ & n51924;
  assign n53788 = P1_P1_REIP_REG_19_ & n52069;
  assign n53789 = P1_P1_INSTADDRPOINTER_REG_18_ & n53718;
  assign n53790 = ~P1_P1_INSTADDRPOINTER_REG_19_ & n53789;
  assign n53791 = P1_P1_INSTADDRPOINTER_REG_19_ & ~n53789;
  assign n53792 = ~n53790 & ~n53791;
  assign n53793 = ~n43812 & ~n53792;
  assign n53794 = n43925 & ~n53792;
  assign n53795 = n43765 & ~n53792;
  assign n53796 = ~n53794 & ~n53795;
  assign n53797 = P1_P1_INSTADDRPOINTER_REG_18_ & n53650;
  assign n53798 = ~P1_P1_INSTADDRPOINTER_REG_19_ & ~n53797;
  assign n53799 = P1_P1_INSTADDRPOINTER_REG_18_ & P1_P1_INSTADDRPOINTER_REG_19_;
  assign n53800 = P1_P1_INSTADDRPOINTER_REG_16_ & n53799;
  assign n53801 = P1_P1_INSTADDRPOINTER_REG_17_ & n53800;
  assign n53802 = n53501 & n53801;
  assign n53803 = ~n53798 & ~n53802;
  assign n53804 = n52032 & n53803;
  assign n53805 = n52049 & ~n53792;
  assign n53806 = n43769 & ~n53792;
  assign n53807 = n52038 & ~n53792;
  assign n53808 = n52042 & ~n53792;
  assign n53809 = ~n53805 & ~n53806;
  assign n53810 = ~n53807 & n53809;
  assign n53811 = ~n53808 & n53810;
  assign n53812 = P1_P1_INSTADDRPOINTER_REG_18_ & n53737;
  assign n53813 = ~P1_P1_INSTADDRPOINTER_REG_19_ & n53812;
  assign n53814 = P1_P1_INSTADDRPOINTER_REG_19_ & ~n53812;
  assign n53815 = ~n53813 & ~n53814;
  assign n53816 = n43625 & ~n53815;
  assign n53817 = n43703 & ~n53815;
  assign n53818 = n43707 & ~n53815;
  assign n53819 = P1_P1_INSTADDRPOINTER_REG_18_ & n53744;
  assign n53820 = ~P1_P1_INSTADDRPOINTER_REG_19_ & n53819;
  assign n53821 = P1_P1_INSTADDRPOINTER_REG_19_ & ~n53819;
  assign n53822 = ~n53820 & ~n53821;
  assign n53823 = n43723 & ~n53822;
  assign n53824 = n43715 & ~n53822;
  assign n53825 = ~n53816 & ~n53817;
  assign n53826 = ~n53818 & n53825;
  assign n53827 = ~n53823 & n53826;
  assign n53828 = ~n53824 & n53827;
  assign n53829 = P1_P1_INSTADDRPOINTER_REG_18_ & n53679;
  assign n53830 = ~P1_P1_INSTADDRPOINTER_REG_19_ & ~n53829;
  assign n53831 = n53530 & n53801;
  assign n53832 = ~n53830 & ~n53831;
  assign n53833 = n43726 & n53832;
  assign n53834 = n53811 & n53828;
  assign n53835 = ~n53833 & n53834;
  assign n53836 = n43883 & ~n53815;
  assign n53837 = n43884 & ~n53815;
  assign n53838 = n51933 & ~n53792;
  assign n53839 = n43699 & ~n53815;
  assign n53840 = n51936 & ~n53792;
  assign n53841 = ~n53839 & ~n53840;
  assign n53842 = ~P1_P1_INSTADDRPOINTER_REG_19_ & ~n52920;
  assign n53843 = P1_P1_INSTADDRPOINTER_REG_19_ & n52920;
  assign n53844 = ~n53842 & ~n53843;
  assign n53845 = ~P1_P1_INSTADDRPOINTER_REG_18_ & n52920;
  assign n53846 = ~n53768 & ~n53845;
  assign n53847 = P1_P1_INSTADDRPOINTER_REG_18_ & ~n52920;
  assign n53848 = ~n53846 & ~n53847;
  assign n53849 = ~n53844 & n53848;
  assign n53850 = ~P1_P1_INSTADDRPOINTER_REG_19_ & n52920;
  assign n53851 = P1_P1_INSTADDRPOINTER_REG_19_ & ~n52920;
  assign n53852 = ~n53850 & ~n53851;
  assign n53853 = ~n53848 & ~n53852;
  assign n53854 = ~n53849 & ~n53853;
  assign n53855 = n52030 & ~n53854;
  assign n53856 = ~n53836 & ~n53837;
  assign n53857 = ~n53838 & n53856;
  assign n53858 = n53841 & n53857;
  assign n53859 = ~n53855 & n53858;
  assign n53860 = ~n53793 & n53796;
  assign n53861 = ~n53804 & n53860;
  assign n53862 = n53835 & n53861;
  assign n53863 = n53859 & n53862;
  assign n53864 = n51925 & ~n53863;
  assign n53865 = ~n53787 & ~n53788;
  assign n8891 = n53864 | ~n53865;
  assign n53867 = P1_P1_INSTADDRPOINTER_REG_20_ & n51924;
  assign n53868 = P1_P1_REIP_REG_20_ & n52069;
  assign n53869 = P1_P1_INSTADDRPOINTER_REG_19_ & n53789;
  assign n53870 = ~P1_P1_INSTADDRPOINTER_REG_20_ & n53869;
  assign n53871 = P1_P1_INSTADDRPOINTER_REG_20_ & ~n53869;
  assign n53872 = ~n53870 & ~n53871;
  assign n53873 = ~n43812 & ~n53872;
  assign n53874 = n43925 & ~n53872;
  assign n53875 = n43765 & ~n53872;
  assign n53876 = ~n53874 & ~n53875;
  assign n53877 = ~P1_P1_INSTADDRPOINTER_REG_20_ & ~n53802;
  assign n53878 = P1_P1_INSTADDRPOINTER_REG_20_ & n53802;
  assign n53879 = ~n53877 & ~n53878;
  assign n53880 = n52032 & n53879;
  assign n53881 = n52049 & ~n53872;
  assign n53882 = n43769 & ~n53872;
  assign n53883 = n52038 & ~n53872;
  assign n53884 = n52042 & ~n53872;
  assign n53885 = ~n53881 & ~n53882;
  assign n53886 = ~n53883 & n53885;
  assign n53887 = ~n53884 & n53886;
  assign n53888 = P1_P1_INSTADDRPOINTER_REG_19_ & n53812;
  assign n53889 = ~P1_P1_INSTADDRPOINTER_REG_20_ & n53888;
  assign n53890 = P1_P1_INSTADDRPOINTER_REG_20_ & ~n53888;
  assign n53891 = ~n53889 & ~n53890;
  assign n53892 = n43625 & ~n53891;
  assign n53893 = n43703 & ~n53891;
  assign n53894 = n43707 & ~n53891;
  assign n53895 = P1_P1_INSTADDRPOINTER_REG_19_ & n53819;
  assign n53896 = ~P1_P1_INSTADDRPOINTER_REG_20_ & n53895;
  assign n53897 = P1_P1_INSTADDRPOINTER_REG_20_ & ~n53895;
  assign n53898 = ~n53896 & ~n53897;
  assign n53899 = n43723 & ~n53898;
  assign n53900 = n43715 & ~n53898;
  assign n53901 = ~n53892 & ~n53893;
  assign n53902 = ~n53894 & n53901;
  assign n53903 = ~n53899 & n53902;
  assign n53904 = ~n53900 & n53903;
  assign n53905 = ~P1_P1_INSTADDRPOINTER_REG_20_ & ~n53831;
  assign n53906 = P1_P1_INSTADDRPOINTER_REG_20_ & n53831;
  assign n53907 = ~n53905 & ~n53906;
  assign n53908 = n43726 & n53907;
  assign n53909 = n53887 & n53904;
  assign n53910 = ~n53908 & n53909;
  assign n53911 = n43883 & ~n53891;
  assign n53912 = n43884 & ~n53891;
  assign n53913 = n51933 & ~n53872;
  assign n53914 = n43699 & ~n53891;
  assign n53915 = n51936 & ~n53872;
  assign n53916 = ~n53914 & ~n53915;
  assign n53917 = P1_P1_INSTADDRPOINTER_REG_19_ & P1_P1_INSTADDRPOINTER_REG_20_;
  assign n53918 = n52920 & ~n53917;
  assign n53919 = P1_P1_INSTADDRPOINTER_REG_20_ & ~n52920;
  assign n53920 = ~n53918 & ~n53919;
  assign n53921 = n53848 & ~n53851;
  assign n53922 = n53920 & ~n53921;
  assign n53923 = ~P1_P1_INSTADDRPOINTER_REG_19_ & n53848;
  assign n53924 = P1_P1_INSTADDRPOINTER_REG_20_ & n53923;
  assign n53925 = ~n52920 & ~n53924;
  assign n53926 = P1_P1_INSTADDRPOINTER_REG_20_ & n52920;
  assign n53927 = P1_P1_INSTADDRPOINTER_REG_19_ & ~n53848;
  assign n53928 = ~n53925 & ~n53926;
  assign n53929 = ~n53927 & n53928;
  assign n53930 = ~n53922 & ~n53929;
  assign n53931 = n52030 & n53930;
  assign n53932 = ~n53911 & ~n53912;
  assign n53933 = ~n53913 & n53932;
  assign n53934 = n53916 & n53933;
  assign n53935 = ~n53931 & n53934;
  assign n53936 = ~n53873 & n53876;
  assign n53937 = ~n53880 & n53936;
  assign n53938 = n53910 & n53937;
  assign n53939 = n53935 & n53938;
  assign n53940 = n51925 & ~n53939;
  assign n53941 = ~n53867 & ~n53868;
  assign n8896 = n53940 | ~n53941;
  assign n53943 = P1_P1_INSTADDRPOINTER_REG_21_ & n51924;
  assign n53944 = P1_P1_REIP_REG_21_ & n52069;
  assign n53945 = P1_P1_INSTADDRPOINTER_REG_20_ & n53869;
  assign n53946 = ~P1_P1_INSTADDRPOINTER_REG_21_ & n53945;
  assign n53947 = P1_P1_INSTADDRPOINTER_REG_21_ & ~n53945;
  assign n53948 = ~n53946 & ~n53947;
  assign n53949 = ~n43812 & ~n53948;
  assign n53950 = n43925 & ~n53948;
  assign n53951 = n43765 & ~n53948;
  assign n53952 = ~n53950 & ~n53951;
  assign n53953 = ~P1_P1_INSTADDRPOINTER_REG_21_ & ~n53878;
  assign n53954 = P1_P1_INSTADDRPOINTER_REG_20_ & P1_P1_INSTADDRPOINTER_REG_21_;
  assign n53955 = n53802 & n53954;
  assign n53956 = ~n53953 & ~n53955;
  assign n53957 = n52032 & n53956;
  assign n53958 = n52049 & ~n53948;
  assign n53959 = n43769 & ~n53948;
  assign n53960 = n52038 & ~n53948;
  assign n53961 = n52042 & ~n53948;
  assign n53962 = ~n53958 & ~n53959;
  assign n53963 = ~n53960 & n53962;
  assign n53964 = ~n53961 & n53963;
  assign n53965 = P1_P1_INSTADDRPOINTER_REG_20_ & n53888;
  assign n53966 = ~P1_P1_INSTADDRPOINTER_REG_21_ & n53965;
  assign n53967 = P1_P1_INSTADDRPOINTER_REG_21_ & ~n53965;
  assign n53968 = ~n53966 & ~n53967;
  assign n53969 = n43625 & ~n53968;
  assign n53970 = n43703 & ~n53968;
  assign n53971 = n43707 & ~n53968;
  assign n53972 = P1_P1_INSTADDRPOINTER_REG_20_ & n53895;
  assign n53973 = ~P1_P1_INSTADDRPOINTER_REG_21_ & n53972;
  assign n53974 = P1_P1_INSTADDRPOINTER_REG_21_ & ~n53972;
  assign n53975 = ~n53973 & ~n53974;
  assign n53976 = n43723 & ~n53975;
  assign n53977 = n43715 & ~n53975;
  assign n53978 = ~n53969 & ~n53970;
  assign n53979 = ~n53971 & n53978;
  assign n53980 = ~n53976 & n53979;
  assign n53981 = ~n53977 & n53980;
  assign n53982 = ~P1_P1_INSTADDRPOINTER_REG_21_ & ~n53906;
  assign n53983 = n53831 & n53954;
  assign n53984 = ~n53982 & ~n53983;
  assign n53985 = n43726 & n53984;
  assign n53986 = n53964 & n53981;
  assign n53987 = ~n53985 & n53986;
  assign n53988 = n43883 & ~n53968;
  assign n53989 = n43884 & ~n53968;
  assign n53990 = n51933 & ~n53948;
  assign n53991 = n43699 & ~n53968;
  assign n53992 = n51936 & ~n53948;
  assign n53993 = ~n53991 & ~n53992;
  assign n53994 = ~n53848 & n53917;
  assign n53995 = ~n53919 & ~n53994;
  assign n53996 = ~n52920 & ~n53923;
  assign n53997 = n53995 & ~n53996;
  assign n53998 = ~P1_P1_INSTADDRPOINTER_REG_21_ & ~n52920;
  assign n53999 = P1_P1_INSTADDRPOINTER_REG_21_ & n52920;
  assign n54000 = ~n53998 & ~n53999;
  assign n54001 = n53997 & ~n54000;
  assign n54002 = ~n53997 & n54000;
  assign n54003 = ~n54001 & ~n54002;
  assign n54004 = n52030 & ~n54003;
  assign n54005 = ~n53988 & ~n53989;
  assign n54006 = ~n53990 & n54005;
  assign n54007 = n53993 & n54006;
  assign n54008 = ~n54004 & n54007;
  assign n54009 = ~n53949 & n53952;
  assign n54010 = ~n53957 & n54009;
  assign n54011 = n53987 & n54010;
  assign n54012 = n54008 & n54011;
  assign n54013 = n51925 & ~n54012;
  assign n54014 = ~n53943 & ~n53944;
  assign n8901 = n54013 | ~n54014;
  assign n54016 = P1_P1_INSTADDRPOINTER_REG_22_ & n51924;
  assign n54017 = P1_P1_REIP_REG_22_ & n52069;
  assign n54018 = P1_P1_INSTADDRPOINTER_REG_21_ & n53945;
  assign n54019 = ~P1_P1_INSTADDRPOINTER_REG_22_ & n54018;
  assign n54020 = P1_P1_INSTADDRPOINTER_REG_22_ & ~n54018;
  assign n54021 = ~n54019 & ~n54020;
  assign n54022 = ~n43812 & ~n54021;
  assign n54023 = n43925 & ~n54021;
  assign n54024 = n43765 & ~n54021;
  assign n54025 = ~n54023 & ~n54024;
  assign n54026 = ~P1_P1_INSTADDRPOINTER_REG_22_ & n53955;
  assign n54027 = P1_P1_INSTADDRPOINTER_REG_22_ & ~n53955;
  assign n54028 = ~n54026 & ~n54027;
  assign n54029 = n52032 & ~n54028;
  assign n54030 = n52049 & ~n54021;
  assign n54031 = n43769 & ~n54021;
  assign n54032 = n52038 & ~n54021;
  assign n54033 = n52042 & ~n54021;
  assign n54034 = ~n54030 & ~n54031;
  assign n54035 = ~n54032 & n54034;
  assign n54036 = ~n54033 & n54035;
  assign n54037 = P1_P1_INSTADDRPOINTER_REG_21_ & n53965;
  assign n54038 = ~P1_P1_INSTADDRPOINTER_REG_22_ & n54037;
  assign n54039 = P1_P1_INSTADDRPOINTER_REG_22_ & ~n54037;
  assign n54040 = ~n54038 & ~n54039;
  assign n54041 = n43625 & ~n54040;
  assign n54042 = n43703 & ~n54040;
  assign n54043 = n43707 & ~n54040;
  assign n54044 = P1_P1_INSTADDRPOINTER_REG_21_ & n53972;
  assign n54045 = ~P1_P1_INSTADDRPOINTER_REG_22_ & n54044;
  assign n54046 = P1_P1_INSTADDRPOINTER_REG_22_ & ~n54044;
  assign n54047 = ~n54045 & ~n54046;
  assign n54048 = n43723 & ~n54047;
  assign n54049 = n43715 & ~n54047;
  assign n54050 = ~n54041 & ~n54042;
  assign n54051 = ~n54043 & n54050;
  assign n54052 = ~n54048 & n54051;
  assign n54053 = ~n54049 & n54052;
  assign n54054 = ~P1_P1_INSTADDRPOINTER_REG_22_ & n53983;
  assign n54055 = P1_P1_INSTADDRPOINTER_REG_22_ & ~n53983;
  assign n54056 = ~n54054 & ~n54055;
  assign n54057 = n43726 & ~n54056;
  assign n54058 = n54036 & n54053;
  assign n54059 = ~n54057 & n54058;
  assign n54060 = n43883 & ~n54040;
  assign n54061 = n43884 & ~n54040;
  assign n54062 = n51933 & ~n54021;
  assign n54063 = n43699 & ~n54040;
  assign n54064 = n51936 & ~n54021;
  assign n54065 = ~n54063 & ~n54064;
  assign n54066 = P1_P1_INSTADDRPOINTER_REG_21_ & n53917;
  assign n54067 = n52920 & ~n54066;
  assign n54068 = ~n53845 & ~n54067;
  assign n54069 = ~n53768 & n54068;
  assign n54070 = P1_P1_INSTADDRPOINTER_REG_21_ & ~n52920;
  assign n54071 = ~n53847 & ~n54070;
  assign n54072 = ~n53851 & n54071;
  assign n54073 = ~n53919 & n54072;
  assign n54074 = ~n54069 & n54073;
  assign n54075 = ~P1_P1_INSTADDRPOINTER_REG_22_ & ~n52920;
  assign n54076 = P1_P1_INSTADDRPOINTER_REG_22_ & n52920;
  assign n54077 = ~n54075 & ~n54076;
  assign n54078 = n54074 & ~n54077;
  assign n54079 = ~n54074 & n54077;
  assign n54080 = ~n54078 & ~n54079;
  assign n54081 = n52030 & ~n54080;
  assign n54082 = ~n54060 & ~n54061;
  assign n54083 = ~n54062 & n54082;
  assign n54084 = n54065 & n54083;
  assign n54085 = ~n54081 & n54084;
  assign n54086 = ~n54022 & n54025;
  assign n54087 = ~n54029 & n54086;
  assign n54088 = n54059 & n54087;
  assign n54089 = n54085 & n54088;
  assign n54090 = n51925 & ~n54089;
  assign n54091 = ~n54016 & ~n54017;
  assign n8906 = n54090 | ~n54091;
  assign n54093 = P1_P1_INSTADDRPOINTER_REG_23_ & n51924;
  assign n54094 = P1_P1_REIP_REG_23_ & n52069;
  assign n54095 = P1_P1_INSTADDRPOINTER_REG_22_ & n54018;
  assign n54096 = ~P1_P1_INSTADDRPOINTER_REG_23_ & n54095;
  assign n54097 = P1_P1_INSTADDRPOINTER_REG_23_ & ~n54095;
  assign n54098 = ~n54096 & ~n54097;
  assign n54099 = ~n43812 & ~n54098;
  assign n54100 = n43925 & ~n54098;
  assign n54101 = n43765 & ~n54098;
  assign n54102 = ~n54100 & ~n54101;
  assign n54103 = P1_P1_INSTADDRPOINTER_REG_22_ & n53955;
  assign n54104 = ~P1_P1_INSTADDRPOINTER_REG_23_ & ~n54103;
  assign n54105 = P1_P1_INSTADDRPOINTER_REG_22_ & P1_P1_INSTADDRPOINTER_REG_23_;
  assign n54106 = n53955 & n54105;
  assign n54107 = ~n54104 & ~n54106;
  assign n54108 = n52032 & n54107;
  assign n54109 = n52049 & ~n54098;
  assign n54110 = n43769 & ~n54098;
  assign n54111 = n52038 & ~n54098;
  assign n54112 = n52042 & ~n54098;
  assign n54113 = ~n54109 & ~n54110;
  assign n54114 = ~n54111 & n54113;
  assign n54115 = ~n54112 & n54114;
  assign n54116 = P1_P1_INSTADDRPOINTER_REG_22_ & n54037;
  assign n54117 = ~P1_P1_INSTADDRPOINTER_REG_23_ & n54116;
  assign n54118 = P1_P1_INSTADDRPOINTER_REG_23_ & ~n54116;
  assign n54119 = ~n54117 & ~n54118;
  assign n54120 = n43625 & ~n54119;
  assign n54121 = n43703 & ~n54119;
  assign n54122 = n43707 & ~n54119;
  assign n54123 = P1_P1_INSTADDRPOINTER_REG_22_ & n54044;
  assign n54124 = ~P1_P1_INSTADDRPOINTER_REG_23_ & n54123;
  assign n54125 = P1_P1_INSTADDRPOINTER_REG_23_ & ~n54123;
  assign n54126 = ~n54124 & ~n54125;
  assign n54127 = n43723 & ~n54126;
  assign n54128 = n43715 & ~n54126;
  assign n54129 = ~n54120 & ~n54121;
  assign n54130 = ~n54122 & n54129;
  assign n54131 = ~n54127 & n54130;
  assign n54132 = ~n54128 & n54131;
  assign n54133 = P1_P1_INSTADDRPOINTER_REG_22_ & n53983;
  assign n54134 = ~P1_P1_INSTADDRPOINTER_REG_23_ & ~n54133;
  assign n54135 = P1_P1_INSTADDRPOINTER_REG_22_ & n53954;
  assign n54136 = P1_P1_INSTADDRPOINTER_REG_23_ & n54135;
  assign n54137 = n53831 & n54136;
  assign n54138 = ~n54134 & ~n54137;
  assign n54139 = n43726 & n54138;
  assign n54140 = n54115 & n54132;
  assign n54141 = ~n54139 & n54140;
  assign n54142 = n43883 & ~n54119;
  assign n54143 = n43884 & ~n54119;
  assign n54144 = n51933 & ~n54098;
  assign n54145 = n43699 & ~n54119;
  assign n54146 = n51936 & ~n54098;
  assign n54147 = ~n54145 & ~n54146;
  assign n54148 = ~P1_P1_INSTADDRPOINTER_REG_22_ & n52920;
  assign n54149 = n54068 & ~n54148;
  assign n54150 = ~n53768 & n54149;
  assign n54151 = P1_P1_INSTADDRPOINTER_REG_22_ & ~n52920;
  assign n54152 = n54073 & ~n54151;
  assign n54153 = ~n54150 & n54152;
  assign n54154 = ~P1_P1_INSTADDRPOINTER_REG_23_ & ~n52920;
  assign n54155 = P1_P1_INSTADDRPOINTER_REG_23_ & n52920;
  assign n54156 = ~n54154 & ~n54155;
  assign n54157 = n54153 & ~n54156;
  assign n54158 = ~n54153 & n54156;
  assign n54159 = ~n54157 & ~n54158;
  assign n54160 = n52030 & ~n54159;
  assign n54161 = ~n54142 & ~n54143;
  assign n54162 = ~n54144 & n54161;
  assign n54163 = n54147 & n54162;
  assign n54164 = ~n54160 & n54163;
  assign n54165 = ~n54099 & n54102;
  assign n54166 = ~n54108 & n54165;
  assign n54167 = n54141 & n54166;
  assign n54168 = n54164 & n54167;
  assign n54169 = n51925 & ~n54168;
  assign n54170 = ~n54093 & ~n54094;
  assign n8911 = n54169 | ~n54170;
  assign n54172 = P1_P1_INSTADDRPOINTER_REG_24_ & n51924;
  assign n54173 = P1_P1_REIP_REG_24_ & n52069;
  assign n54174 = P1_P1_INSTADDRPOINTER_REG_23_ & n54095;
  assign n54175 = ~P1_P1_INSTADDRPOINTER_REG_24_ & n54174;
  assign n54176 = P1_P1_INSTADDRPOINTER_REG_24_ & ~n54174;
  assign n54177 = ~n54175 & ~n54176;
  assign n54178 = ~n43812 & ~n54177;
  assign n54179 = n43925 & ~n54177;
  assign n54180 = n43765 & ~n54177;
  assign n54181 = ~n54179 & ~n54180;
  assign n54182 = ~P1_P1_INSTADDRPOINTER_REG_24_ & n54106;
  assign n54183 = P1_P1_INSTADDRPOINTER_REG_24_ & ~n54106;
  assign n54184 = ~n54182 & ~n54183;
  assign n54185 = n52032 & ~n54184;
  assign n54186 = n52049 & ~n54177;
  assign n54187 = n43769 & ~n54177;
  assign n54188 = n52038 & ~n54177;
  assign n54189 = n52042 & ~n54177;
  assign n54190 = ~n54186 & ~n54187;
  assign n54191 = ~n54188 & n54190;
  assign n54192 = ~n54189 & n54191;
  assign n54193 = P1_P1_INSTADDRPOINTER_REG_23_ & n54116;
  assign n54194 = ~P1_P1_INSTADDRPOINTER_REG_24_ & n54193;
  assign n54195 = P1_P1_INSTADDRPOINTER_REG_24_ & ~n54193;
  assign n54196 = ~n54194 & ~n54195;
  assign n54197 = n43625 & ~n54196;
  assign n54198 = n43703 & ~n54196;
  assign n54199 = n43707 & ~n54196;
  assign n54200 = P1_P1_INSTADDRPOINTER_REG_23_ & n54123;
  assign n54201 = ~P1_P1_INSTADDRPOINTER_REG_24_ & n54200;
  assign n54202 = P1_P1_INSTADDRPOINTER_REG_24_ & ~n54200;
  assign n54203 = ~n54201 & ~n54202;
  assign n54204 = n43723 & ~n54203;
  assign n54205 = n43715 & ~n54203;
  assign n54206 = ~n54197 & ~n54198;
  assign n54207 = ~n54199 & n54206;
  assign n54208 = ~n54204 & n54207;
  assign n54209 = ~n54205 & n54208;
  assign n54210 = ~P1_P1_INSTADDRPOINTER_REG_24_ & n54137;
  assign n54211 = P1_P1_INSTADDRPOINTER_REG_24_ & ~n54137;
  assign n54212 = ~n54210 & ~n54211;
  assign n54213 = n43726 & ~n54212;
  assign n54214 = n54192 & n54209;
  assign n54215 = ~n54213 & n54214;
  assign n54216 = n43883 & ~n54196;
  assign n54217 = n43884 & ~n54196;
  assign n54218 = n51933 & ~n54177;
  assign n54219 = n43699 & ~n54196;
  assign n54220 = n51936 & ~n54177;
  assign n54221 = ~n54219 & ~n54220;
  assign n54222 = ~P1_P1_INSTADDRPOINTER_REG_23_ & n52920;
  assign n54223 = n54149 & ~n54222;
  assign n54224 = ~n53768 & n54223;
  assign n54225 = P1_P1_INSTADDRPOINTER_REG_23_ & ~n52920;
  assign n54226 = n54152 & ~n54225;
  assign n54227 = ~n54224 & n54226;
  assign n54228 = ~P1_P1_INSTADDRPOINTER_REG_24_ & ~n52920;
  assign n54229 = P1_P1_INSTADDRPOINTER_REG_24_ & n52920;
  assign n54230 = ~n54228 & ~n54229;
  assign n54231 = n54227 & ~n54230;
  assign n54232 = ~n54227 & n54230;
  assign n54233 = ~n54231 & ~n54232;
  assign n54234 = n52030 & ~n54233;
  assign n54235 = ~n54216 & ~n54217;
  assign n54236 = ~n54218 & n54235;
  assign n54237 = n54221 & n54236;
  assign n54238 = ~n54234 & n54237;
  assign n54239 = ~n54178 & n54181;
  assign n54240 = ~n54185 & n54239;
  assign n54241 = n54215 & n54240;
  assign n54242 = n54238 & n54241;
  assign n54243 = n51925 & ~n54242;
  assign n54244 = ~n54172 & ~n54173;
  assign n8916 = n54243 | ~n54244;
  assign n54246 = P1_P1_INSTADDRPOINTER_REG_25_ & n51924;
  assign n54247 = P1_P1_REIP_REG_25_ & n52069;
  assign n54248 = P1_P1_INSTADDRPOINTER_REG_24_ & n54174;
  assign n54249 = ~P1_P1_INSTADDRPOINTER_REG_25_ & n54248;
  assign n54250 = P1_P1_INSTADDRPOINTER_REG_25_ & ~n54248;
  assign n54251 = ~n54249 & ~n54250;
  assign n54252 = ~n43812 & ~n54251;
  assign n54253 = n43925 & ~n54251;
  assign n54254 = n43765 & ~n54251;
  assign n54255 = ~n54253 & ~n54254;
  assign n54256 = P1_P1_INSTADDRPOINTER_REG_24_ & n54106;
  assign n54257 = ~P1_P1_INSTADDRPOINTER_REG_25_ & ~n54256;
  assign n54258 = P1_P1_INSTADDRPOINTER_REG_24_ & P1_P1_INSTADDRPOINTER_REG_25_;
  assign n54259 = n54106 & n54258;
  assign n54260 = ~n54257 & ~n54259;
  assign n54261 = n52032 & n54260;
  assign n54262 = n52049 & ~n54251;
  assign n54263 = n43769 & ~n54251;
  assign n54264 = n52038 & ~n54251;
  assign n54265 = n52042 & ~n54251;
  assign n54266 = ~n54262 & ~n54263;
  assign n54267 = ~n54264 & n54266;
  assign n54268 = ~n54265 & n54267;
  assign n54269 = P1_P1_INSTADDRPOINTER_REG_24_ & n54193;
  assign n54270 = ~P1_P1_INSTADDRPOINTER_REG_25_ & n54269;
  assign n54271 = P1_P1_INSTADDRPOINTER_REG_25_ & ~n54269;
  assign n54272 = ~n54270 & ~n54271;
  assign n54273 = n43625 & ~n54272;
  assign n54274 = n43703 & ~n54272;
  assign n54275 = n43707 & ~n54272;
  assign n54276 = P1_P1_INSTADDRPOINTER_REG_24_ & n54200;
  assign n54277 = ~P1_P1_INSTADDRPOINTER_REG_25_ & n54276;
  assign n54278 = P1_P1_INSTADDRPOINTER_REG_25_ & ~n54276;
  assign n54279 = ~n54277 & ~n54278;
  assign n54280 = n43723 & ~n54279;
  assign n54281 = n43715 & ~n54279;
  assign n54282 = ~n54273 & ~n54274;
  assign n54283 = ~n54275 & n54282;
  assign n54284 = ~n54280 & n54283;
  assign n54285 = ~n54281 & n54284;
  assign n54286 = P1_P1_INSTADDRPOINTER_REG_24_ & n54137;
  assign n54287 = ~P1_P1_INSTADDRPOINTER_REG_25_ & ~n54286;
  assign n54288 = n54137 & n54258;
  assign n54289 = ~n54287 & ~n54288;
  assign n54290 = n43726 & n54289;
  assign n54291 = n54268 & n54285;
  assign n54292 = ~n54290 & n54291;
  assign n54293 = n43883 & ~n54272;
  assign n54294 = n43884 & ~n54272;
  assign n54295 = n51933 & ~n54251;
  assign n54296 = n43699 & ~n54272;
  assign n54297 = n51936 & ~n54251;
  assign n54298 = ~n54296 & ~n54297;
  assign n54299 = ~P1_P1_INSTADDRPOINTER_REG_25_ & ~n52920;
  assign n54300 = P1_P1_INSTADDRPOINTER_REG_25_ & n52920;
  assign n54301 = ~n54299 & ~n54300;
  assign n54302 = P1_P1_INSTADDRPOINTER_REG_24_ & ~n52920;
  assign n54303 = n54226 & ~n54302;
  assign n54304 = ~P1_P1_INSTADDRPOINTER_REG_24_ & n52920;
  assign n54305 = n54223 & ~n54304;
  assign n54306 = ~n53768 & n54305;
  assign n54307 = n54303 & ~n54306;
  assign n54308 = ~n54301 & n54307;
  assign n54309 = ~P1_P1_INSTADDRPOINTER_REG_25_ & n52920;
  assign n54310 = P1_P1_INSTADDRPOINTER_REG_25_ & ~n52920;
  assign n54311 = ~n54309 & ~n54310;
  assign n54312 = ~n54307 & ~n54311;
  assign n54313 = ~n54308 & ~n54312;
  assign n54314 = n52030 & ~n54313;
  assign n54315 = ~n54293 & ~n54294;
  assign n54316 = ~n54295 & n54315;
  assign n54317 = n54298 & n54316;
  assign n54318 = ~n54314 & n54317;
  assign n54319 = ~n54252 & n54255;
  assign n54320 = ~n54261 & n54319;
  assign n54321 = n54292 & n54320;
  assign n54322 = n54318 & n54321;
  assign n54323 = n51925 & ~n54322;
  assign n54324 = ~n54246 & ~n54247;
  assign n8921 = n54323 | ~n54324;
  assign n54326 = P1_P1_INSTADDRPOINTER_REG_26_ & n51924;
  assign n54327 = P1_P1_REIP_REG_26_ & n52069;
  assign n54328 = P1_P1_INSTADDRPOINTER_REG_25_ & n54248;
  assign n54329 = ~P1_P1_INSTADDRPOINTER_REG_26_ & n54328;
  assign n54330 = P1_P1_INSTADDRPOINTER_REG_26_ & ~n54328;
  assign n54331 = ~n54329 & ~n54330;
  assign n54332 = ~n43812 & ~n54331;
  assign n54333 = n43925 & ~n54331;
  assign n54334 = n43765 & ~n54331;
  assign n54335 = ~n54333 & ~n54334;
  assign n54336 = ~P1_P1_INSTADDRPOINTER_REG_26_ & ~n54259;
  assign n54337 = P1_P1_INSTADDRPOINTER_REG_26_ & n54259;
  assign n54338 = ~n54336 & ~n54337;
  assign n54339 = n52032 & n54338;
  assign n54340 = n52049 & ~n54331;
  assign n54341 = n43769 & ~n54331;
  assign n54342 = n52038 & ~n54331;
  assign n54343 = n52042 & ~n54331;
  assign n54344 = ~n54340 & ~n54341;
  assign n54345 = ~n54342 & n54344;
  assign n54346 = ~n54343 & n54345;
  assign n54347 = P1_P1_INSTADDRPOINTER_REG_25_ & n54269;
  assign n54348 = ~P1_P1_INSTADDRPOINTER_REG_26_ & n54347;
  assign n54349 = P1_P1_INSTADDRPOINTER_REG_26_ & ~n54347;
  assign n54350 = ~n54348 & ~n54349;
  assign n54351 = n43625 & ~n54350;
  assign n54352 = n43703 & ~n54350;
  assign n54353 = n43707 & ~n54350;
  assign n54354 = P1_P1_INSTADDRPOINTER_REG_25_ & n54276;
  assign n54355 = ~P1_P1_INSTADDRPOINTER_REG_26_ & n54354;
  assign n54356 = P1_P1_INSTADDRPOINTER_REG_26_ & ~n54354;
  assign n54357 = ~n54355 & ~n54356;
  assign n54358 = n43723 & ~n54357;
  assign n54359 = n43715 & ~n54357;
  assign n54360 = ~n54351 & ~n54352;
  assign n54361 = ~n54353 & n54360;
  assign n54362 = ~n54358 & n54361;
  assign n54363 = ~n54359 & n54362;
  assign n54364 = ~P1_P1_INSTADDRPOINTER_REG_26_ & ~n54288;
  assign n54365 = P1_P1_INSTADDRPOINTER_REG_26_ & n54288;
  assign n54366 = ~n54364 & ~n54365;
  assign n54367 = n43726 & n54366;
  assign n54368 = n54346 & n54363;
  assign n54369 = ~n54367 & n54368;
  assign n54370 = n43883 & ~n54350;
  assign n54371 = n43884 & ~n54350;
  assign n54372 = n51933 & ~n54331;
  assign n54373 = n43699 & ~n54350;
  assign n54374 = n51936 & ~n54331;
  assign n54375 = ~n54373 & ~n54374;
  assign n54376 = P1_P1_INSTADDRPOINTER_REG_26_ & ~n52920;
  assign n54377 = P1_P1_INSTADDRPOINTER_REG_25_ & P1_P1_INSTADDRPOINTER_REG_26_;
  assign n54378 = n52920 & ~n54377;
  assign n54379 = ~n54376 & ~n54378;
  assign n54380 = n54307 & ~n54310;
  assign n54381 = n54379 & ~n54380;
  assign n54382 = ~P1_P1_INSTADDRPOINTER_REG_26_ & ~n52920;
  assign n54383 = P1_P1_INSTADDRPOINTER_REG_26_ & n52920;
  assign n54384 = ~n54382 & ~n54383;
  assign n54385 = ~n54310 & n54384;
  assign n54386 = ~n54307 & ~n54309;
  assign n54387 = n54385 & ~n54386;
  assign n54388 = ~n54381 & ~n54387;
  assign n54389 = n52030 & n54388;
  assign n54390 = ~n54370 & ~n54371;
  assign n54391 = ~n54372 & n54390;
  assign n54392 = n54375 & n54391;
  assign n54393 = ~n54389 & n54392;
  assign n54394 = ~n54332 & n54335;
  assign n54395 = ~n54339 & n54394;
  assign n54396 = n54369 & n54395;
  assign n54397 = n54393 & n54396;
  assign n54398 = n51925 & ~n54397;
  assign n54399 = ~n54326 & ~n54327;
  assign n8926 = n54398 | ~n54399;
  assign n54401 = P1_P1_INSTADDRPOINTER_REG_27_ & n51924;
  assign n54402 = P1_P1_REIP_REG_27_ & n52069;
  assign n54403 = P1_P1_INSTADDRPOINTER_REG_26_ & n54328;
  assign n54404 = ~P1_P1_INSTADDRPOINTER_REG_27_ & n54403;
  assign n54405 = P1_P1_INSTADDRPOINTER_REG_27_ & ~n54403;
  assign n54406 = ~n54404 & ~n54405;
  assign n54407 = ~n43812 & ~n54406;
  assign n54408 = n43925 & ~n54406;
  assign n54409 = n43765 & ~n54406;
  assign n54410 = ~n54408 & ~n54409;
  assign n54411 = ~P1_P1_INSTADDRPOINTER_REG_27_ & n54337;
  assign n54412 = P1_P1_INSTADDRPOINTER_REG_27_ & ~n54337;
  assign n54413 = ~n54411 & ~n54412;
  assign n54414 = n52032 & ~n54413;
  assign n54415 = n52049 & ~n54406;
  assign n54416 = n43769 & ~n54406;
  assign n54417 = n52038 & ~n54406;
  assign n54418 = n52042 & ~n54406;
  assign n54419 = ~n54415 & ~n54416;
  assign n54420 = ~n54417 & n54419;
  assign n54421 = ~n54418 & n54420;
  assign n54422 = P1_P1_INSTADDRPOINTER_REG_26_ & n54347;
  assign n54423 = ~P1_P1_INSTADDRPOINTER_REG_27_ & n54422;
  assign n54424 = P1_P1_INSTADDRPOINTER_REG_27_ & ~n54422;
  assign n54425 = ~n54423 & ~n54424;
  assign n54426 = n43625 & ~n54425;
  assign n54427 = n43703 & ~n54425;
  assign n54428 = n43707 & ~n54425;
  assign n54429 = P1_P1_INSTADDRPOINTER_REG_26_ & n54354;
  assign n54430 = ~P1_P1_INSTADDRPOINTER_REG_27_ & n54429;
  assign n54431 = P1_P1_INSTADDRPOINTER_REG_27_ & ~n54429;
  assign n54432 = ~n54430 & ~n54431;
  assign n54433 = n43723 & ~n54432;
  assign n54434 = n43715 & ~n54432;
  assign n54435 = ~n54426 & ~n54427;
  assign n54436 = ~n54428 & n54435;
  assign n54437 = ~n54433 & n54436;
  assign n54438 = ~n54434 & n54437;
  assign n54439 = ~P1_P1_INSTADDRPOINTER_REG_27_ & n54365;
  assign n54440 = P1_P1_INSTADDRPOINTER_REG_27_ & ~n54365;
  assign n54441 = ~n54439 & ~n54440;
  assign n54442 = n43726 & ~n54441;
  assign n54443 = n54421 & n54438;
  assign n54444 = ~n54442 & n54443;
  assign n54445 = n43883 & ~n54425;
  assign n54446 = n43884 & ~n54425;
  assign n54447 = n51933 & ~n54406;
  assign n54448 = n43699 & ~n54425;
  assign n54449 = n51936 & ~n54406;
  assign n54450 = ~n54448 & ~n54449;
  assign n54451 = ~n54310 & ~n54376;
  assign n54452 = ~n54307 & ~n54378;
  assign n54453 = n54451 & ~n54452;
  assign n54454 = ~P1_P1_INSTADDRPOINTER_REG_27_ & ~n52920;
  assign n54455 = P1_P1_INSTADDRPOINTER_REG_27_ & n52920;
  assign n54456 = ~n54454 & ~n54455;
  assign n54457 = n54453 & ~n54456;
  assign n54458 = ~n54453 & n54456;
  assign n54459 = ~n54457 & ~n54458;
  assign n54460 = n52030 & ~n54459;
  assign n54461 = ~n54445 & ~n54446;
  assign n54462 = ~n54447 & n54461;
  assign n54463 = n54450 & n54462;
  assign n54464 = ~n54460 & n54463;
  assign n54465 = ~n54407 & n54410;
  assign n54466 = ~n54414 & n54465;
  assign n54467 = n54444 & n54466;
  assign n54468 = n54464 & n54467;
  assign n54469 = n51925 & ~n54468;
  assign n54470 = ~n54401 & ~n54402;
  assign n8931 = n54469 | ~n54470;
  assign n54472 = P1_P1_INSTADDRPOINTER_REG_28_ & n51924;
  assign n54473 = P1_P1_REIP_REG_28_ & n52069;
  assign n54474 = P1_P1_INSTADDRPOINTER_REG_27_ & n54403;
  assign n54475 = ~P1_P1_INSTADDRPOINTER_REG_28_ & n54474;
  assign n54476 = P1_P1_INSTADDRPOINTER_REG_28_ & ~n54474;
  assign n54477 = ~n54475 & ~n54476;
  assign n54478 = ~n43812 & ~n54477;
  assign n54479 = n43925 & ~n54477;
  assign n54480 = n43765 & ~n54477;
  assign n54481 = ~n54479 & ~n54480;
  assign n54482 = P1_P1_INSTADDRPOINTER_REG_27_ & n54337;
  assign n54483 = ~P1_P1_INSTADDRPOINTER_REG_28_ & ~n54482;
  assign n54484 = P1_P1_INSTADDRPOINTER_REG_27_ & P1_P1_INSTADDRPOINTER_REG_28_;
  assign n54485 = P1_P1_INSTADDRPOINTER_REG_26_ & n54484;
  assign n54486 = n54259 & n54485;
  assign n54487 = ~n54483 & ~n54486;
  assign n54488 = n52032 & n54487;
  assign n54489 = n52049 & ~n54477;
  assign n54490 = n43769 & ~n54477;
  assign n54491 = n52038 & ~n54477;
  assign n54492 = n52042 & ~n54477;
  assign n54493 = ~n54489 & ~n54490;
  assign n54494 = ~n54491 & n54493;
  assign n54495 = ~n54492 & n54494;
  assign n54496 = P1_P1_INSTADDRPOINTER_REG_27_ & n54422;
  assign n54497 = ~P1_P1_INSTADDRPOINTER_REG_28_ & n54496;
  assign n54498 = P1_P1_INSTADDRPOINTER_REG_28_ & ~n54496;
  assign n54499 = ~n54497 & ~n54498;
  assign n54500 = n43625 & ~n54499;
  assign n54501 = n43703 & ~n54499;
  assign n54502 = n43707 & ~n54499;
  assign n54503 = P1_P1_INSTADDRPOINTER_REG_27_ & n54429;
  assign n54504 = ~P1_P1_INSTADDRPOINTER_REG_28_ & n54503;
  assign n54505 = P1_P1_INSTADDRPOINTER_REG_28_ & ~n54503;
  assign n54506 = ~n54504 & ~n54505;
  assign n54507 = n43723 & ~n54506;
  assign n54508 = n43715 & ~n54506;
  assign n54509 = ~n54500 & ~n54501;
  assign n54510 = ~n54502 & n54509;
  assign n54511 = ~n54507 & n54510;
  assign n54512 = ~n54508 & n54511;
  assign n54513 = P1_P1_INSTADDRPOINTER_REG_27_ & n54365;
  assign n54514 = ~P1_P1_INSTADDRPOINTER_REG_28_ & ~n54513;
  assign n54515 = P1_P1_INSTADDRPOINTER_REG_25_ & P1_P1_INSTADDRPOINTER_REG_27_;
  assign n54516 = P1_P1_INSTADDRPOINTER_REG_24_ & n54515;
  assign n54517 = P1_P1_INSTADDRPOINTER_REG_26_ & n54516;
  assign n54518 = P1_P1_INSTADDRPOINTER_REG_28_ & n54517;
  assign n54519 = n54137 & n54518;
  assign n54520 = ~n54514 & ~n54519;
  assign n54521 = n43726 & n54520;
  assign n54522 = n54495 & n54512;
  assign n54523 = ~n54521 & n54522;
  assign n54524 = n43883 & ~n54499;
  assign n54525 = n43884 & ~n54499;
  assign n54526 = n51933 & ~n54477;
  assign n54527 = n43699 & ~n54499;
  assign n54528 = n51936 & ~n54477;
  assign n54529 = ~n54527 & ~n54528;
  assign n54530 = ~n54453 & n54484;
  assign n54531 = n52920 & ~n54530;
  assign n54532 = P1_P1_INSTADDRPOINTER_REG_28_ & ~n52920;
  assign n54533 = ~P1_P1_INSTADDRPOINTER_REG_27_ & ~n54310;
  assign n54534 = ~n54376 & n54533;
  assign n54535 = ~n54452 & n54534;
  assign n54536 = ~n54531 & ~n54532;
  assign n54537 = ~n54535 & n54536;
  assign n54538 = P1_P1_INSTADDRPOINTER_REG_28_ & n54535;
  assign n54539 = ~n52920 & ~n54538;
  assign n54540 = P1_P1_INSTADDRPOINTER_REG_28_ & n52920;
  assign n54541 = P1_P1_INSTADDRPOINTER_REG_27_ & ~n54453;
  assign n54542 = ~n54539 & ~n54540;
  assign n54543 = ~n54541 & n54542;
  assign n54544 = ~n54537 & ~n54543;
  assign n54545 = n52030 & n54544;
  assign n54546 = ~n54524 & ~n54525;
  assign n54547 = ~n54526 & n54546;
  assign n54548 = n54529 & n54547;
  assign n54549 = ~n54545 & n54548;
  assign n54550 = ~n54478 & n54481;
  assign n54551 = ~n54488 & n54550;
  assign n54552 = n54523 & n54551;
  assign n54553 = n54549 & n54552;
  assign n54554 = n51925 & ~n54553;
  assign n54555 = ~n54472 & ~n54473;
  assign n8936 = n54554 | ~n54555;
  assign n54557 = P1_P1_INSTADDRPOINTER_REG_29_ & n51924;
  assign n54558 = P1_P1_REIP_REG_29_ & n52069;
  assign n54559 = ~n54557 & ~n54558;
  assign n54560 = ~n52920 & ~n54535;
  assign n54561 = ~n54532 & ~n54560;
  assign n54562 = ~n54530 & n54561;
  assign n54563 = ~P1_P1_INSTADDRPOINTER_REG_29_ & ~n52920;
  assign n54564 = P1_P1_INSTADDRPOINTER_REG_29_ & n52920;
  assign n54565 = ~n54563 & ~n54564;
  assign n54566 = n54562 & ~n54565;
  assign n54567 = ~n54562 & n54565;
  assign n54568 = ~n54566 & ~n54567;
  assign n54569 = n52030 & ~n54568;
  assign n54570 = P1_P1_INSTADDRPOINTER_REG_28_ & n54474;
  assign n54571 = ~P1_P1_INSTADDRPOINTER_REG_29_ & n54570;
  assign n54572 = P1_P1_INSTADDRPOINTER_REG_29_ & ~n54570;
  assign n54573 = ~n54571 & ~n54572;
  assign n54574 = ~n43812 & ~n54573;
  assign n54575 = n43925 & ~n54573;
  assign n54576 = n43765 & ~n54573;
  assign n54577 = ~n54575 & ~n54576;
  assign n54578 = P1_P1_INSTADDRPOINTER_REG_28_ & n54496;
  assign n54579 = ~P1_P1_INSTADDRPOINTER_REG_29_ & n54578;
  assign n54580 = P1_P1_INSTADDRPOINTER_REG_29_ & ~n54578;
  assign n54581 = ~n54579 & ~n54580;
  assign n54582 = n43883 & ~n54581;
  assign n54583 = n43884 & ~n54581;
  assign n54584 = n51933 & ~n54573;
  assign n54585 = n43699 & ~n54581;
  assign n54586 = n51936 & ~n54573;
  assign n54587 = ~n54585 & ~n54586;
  assign n54588 = ~n54582 & ~n54583;
  assign n54589 = ~n54584 & n54588;
  assign n54590 = n54587 & n54589;
  assign n54591 = ~P1_P1_INSTADDRPOINTER_REG_29_ & ~n54486;
  assign n54592 = P1_P1_INSTADDRPOINTER_REG_29_ & n54486;
  assign n54593 = ~n54591 & ~n54592;
  assign n54594 = n52032 & n54593;
  assign n54595 = n52049 & ~n54573;
  assign n54596 = n43769 & ~n54573;
  assign n54597 = n52038 & ~n54573;
  assign n54598 = n52042 & ~n54573;
  assign n54599 = ~n54595 & ~n54596;
  assign n54600 = ~n54597 & n54599;
  assign n54601 = ~n54598 & n54600;
  assign n54602 = n43625 & ~n54581;
  assign n54603 = n43703 & ~n54581;
  assign n54604 = n43707 & ~n54581;
  assign n54605 = P1_P1_INSTADDRPOINTER_REG_28_ & n54503;
  assign n54606 = ~P1_P1_INSTADDRPOINTER_REG_29_ & n54605;
  assign n54607 = P1_P1_INSTADDRPOINTER_REG_29_ & ~n54605;
  assign n54608 = ~n54606 & ~n54607;
  assign n54609 = n43723 & ~n54608;
  assign n54610 = n43715 & ~n54608;
  assign n54611 = ~n54602 & ~n54603;
  assign n54612 = ~n54604 & n54611;
  assign n54613 = ~n54609 & n54612;
  assign n54614 = ~n54610 & n54613;
  assign n54615 = ~P1_P1_INSTADDRPOINTER_REG_29_ & ~n54519;
  assign n54616 = P1_P1_INSTADDRPOINTER_REG_29_ & n54519;
  assign n54617 = ~n54615 & ~n54616;
  assign n54618 = n43726 & n54617;
  assign n54619 = n54601 & n54614;
  assign n54620 = ~n54618 & n54619;
  assign n54621 = ~n54574 & n54577;
  assign n54622 = n54590 & n54621;
  assign n54623 = ~n54594 & n54622;
  assign n54624 = n54620 & n54623;
  assign n54625 = ~n54569 & n54624;
  assign n54626 = n51925 & ~n54625;
  assign n8941 = ~n54559 | n54626;
  assign n54628 = P1_P1_INSTADDRPOINTER_REG_30_ & n51924;
  assign n54629 = P1_P1_REIP_REG_30_ & n52069;
  assign n54630 = ~n54628 & ~n54629;
  assign n54631 = ~P1_P1_INSTADDRPOINTER_REG_30_ & ~n52920;
  assign n54632 = P1_P1_INSTADDRPOINTER_REG_30_ & n52920;
  assign n54633 = ~n54631 & ~n54632;
  assign n54634 = P1_P1_INSTADDRPOINTER_REG_29_ & ~n52920;
  assign n54635 = ~P1_P1_INSTADDRPOINTER_REG_29_ & n52920;
  assign n54636 = ~n54562 & ~n54635;
  assign n54637 = ~n54634 & ~n54636;
  assign n54638 = ~n54633 & n54637;
  assign n54639 = n54633 & ~n54637;
  assign n54640 = ~n54638 & ~n54639;
  assign n54641 = n52030 & ~n54640;
  assign n54642 = P1_P1_INSTADDRPOINTER_REG_29_ & n54570;
  assign n54643 = ~P1_P1_INSTADDRPOINTER_REG_30_ & n54642;
  assign n54644 = P1_P1_INSTADDRPOINTER_REG_30_ & ~n54642;
  assign n54645 = ~n54643 & ~n54644;
  assign n54646 = ~n43812 & ~n54645;
  assign n54647 = n43925 & ~n54645;
  assign n54648 = n43765 & ~n54645;
  assign n54649 = ~n54647 & ~n54648;
  assign n54650 = P1_P1_INSTADDRPOINTER_REG_29_ & n54578;
  assign n54651 = ~P1_P1_INSTADDRPOINTER_REG_30_ & n54650;
  assign n54652 = P1_P1_INSTADDRPOINTER_REG_30_ & ~n54650;
  assign n54653 = ~n54651 & ~n54652;
  assign n54654 = n43883 & ~n54653;
  assign n54655 = n43884 & ~n54653;
  assign n54656 = n51933 & ~n54645;
  assign n54657 = n43699 & ~n54653;
  assign n54658 = n51936 & ~n54645;
  assign n54659 = ~n54657 & ~n54658;
  assign n54660 = ~n54654 & ~n54655;
  assign n54661 = ~n54656 & n54660;
  assign n54662 = n54659 & n54661;
  assign n54663 = ~P1_P1_INSTADDRPOINTER_REG_30_ & n54592;
  assign n54664 = P1_P1_INSTADDRPOINTER_REG_30_ & ~n54592;
  assign n54665 = ~n54663 & ~n54664;
  assign n54666 = n52032 & ~n54665;
  assign n54667 = n52049 & ~n54645;
  assign n54668 = n43769 & ~n54645;
  assign n54669 = n52038 & ~n54645;
  assign n54670 = n52042 & ~n54645;
  assign n54671 = ~n54667 & ~n54668;
  assign n54672 = ~n54669 & n54671;
  assign n54673 = ~n54670 & n54672;
  assign n54674 = n43625 & ~n54653;
  assign n54675 = n43703 & ~n54653;
  assign n54676 = n43707 & ~n54653;
  assign n54677 = P1_P1_INSTADDRPOINTER_REG_29_ & n54605;
  assign n54678 = ~P1_P1_INSTADDRPOINTER_REG_30_ & n54677;
  assign n54679 = P1_P1_INSTADDRPOINTER_REG_30_ & ~n54677;
  assign n54680 = ~n54678 & ~n54679;
  assign n54681 = n43723 & ~n54680;
  assign n54682 = n43715 & ~n54680;
  assign n54683 = ~n54674 & ~n54675;
  assign n54684 = ~n54676 & n54683;
  assign n54685 = ~n54681 & n54684;
  assign n54686 = ~n54682 & n54685;
  assign n54687 = ~P1_P1_INSTADDRPOINTER_REG_30_ & n54616;
  assign n54688 = P1_P1_INSTADDRPOINTER_REG_30_ & ~n54616;
  assign n54689 = ~n54687 & ~n54688;
  assign n54690 = n43726 & ~n54689;
  assign n54691 = n54673 & n54686;
  assign n54692 = ~n54690 & n54691;
  assign n54693 = ~n54646 & n54649;
  assign n54694 = n54662 & n54693;
  assign n54695 = ~n54666 & n54694;
  assign n54696 = n54692 & n54695;
  assign n54697 = ~n54641 & n54696;
  assign n54698 = n51925 & ~n54697;
  assign n8946 = ~n54630 | n54698;
  assign n54700 = P1_P1_INSTADDRPOINTER_REG_31_ & n51924;
  assign n54701 = P1_P1_REIP_REG_31_ & n52069;
  assign n54702 = ~n54700 & ~n54701;
  assign n54703 = P1_P1_INSTADDRPOINTER_REG_31_ & ~n52920;
  assign n54704 = P1_P1_INSTADDRPOINTER_REG_30_ & P1_P1_INSTADDRPOINTER_REG_31_;
  assign n54705 = ~n54635 & n54704;
  assign n54706 = ~n54562 & n54705;
  assign n54707 = n52920 & ~n54706;
  assign n54708 = ~n54703 & ~n54707;
  assign n54709 = ~P1_P1_INSTADDRPOINTER_REG_30_ & n54637;
  assign n54710 = n54708 & ~n54709;
  assign n54711 = ~P1_P1_INSTADDRPOINTER_REG_30_ & ~n54634;
  assign n54712 = P1_P1_INSTADDRPOINTER_REG_31_ & n54711;
  assign n54713 = ~n54532 & n54712;
  assign n54714 = ~n54560 & n54713;
  assign n54715 = ~n52920 & ~n54714;
  assign n54716 = P1_P1_INSTADDRPOINTER_REG_31_ & n52920;
  assign n54717 = ~n54715 & ~n54716;
  assign n54718 = P1_P1_INSTADDRPOINTER_REG_30_ & ~n54637;
  assign n54719 = n54717 & ~n54718;
  assign n54720 = ~n54710 & ~n54719;
  assign n54721 = n52030 & n54720;
  assign n54722 = P1_P1_INSTADDRPOINTER_REG_30_ & n54642;
  assign n54723 = ~P1_P1_INSTADDRPOINTER_REG_31_ & n54722;
  assign n54724 = P1_P1_INSTADDRPOINTER_REG_31_ & ~n54722;
  assign n54725 = ~n54723 & ~n54724;
  assign n54726 = ~n43812 & ~n54725;
  assign n54727 = n43925 & ~n54725;
  assign n54728 = n43765 & ~n54725;
  assign n54729 = ~n54727 & ~n54728;
  assign n54730 = P1_P1_INSTADDRPOINTER_REG_30_ & n54650;
  assign n54731 = ~P1_P1_INSTADDRPOINTER_REG_31_ & n54730;
  assign n54732 = P1_P1_INSTADDRPOINTER_REG_31_ & ~n54730;
  assign n54733 = ~n54731 & ~n54732;
  assign n54734 = n43883 & ~n54733;
  assign n54735 = n43884 & ~n54733;
  assign n54736 = n51933 & ~n54725;
  assign n54737 = n43699 & ~n54733;
  assign n54738 = n51936 & ~n54725;
  assign n54739 = ~n54737 & ~n54738;
  assign n54740 = ~n54734 & ~n54735;
  assign n54741 = ~n54736 & n54740;
  assign n54742 = n54739 & n54741;
  assign n54743 = P1_P1_INSTADDRPOINTER_REG_29_ & P1_P1_INSTADDRPOINTER_REG_30_;
  assign n54744 = n54486 & n54743;
  assign n54745 = ~P1_P1_INSTADDRPOINTER_REG_31_ & n54744;
  assign n54746 = P1_P1_INSTADDRPOINTER_REG_31_ & ~n54744;
  assign n54747 = ~n54745 & ~n54746;
  assign n54748 = n52032 & ~n54747;
  assign n54749 = n52049 & ~n54725;
  assign n54750 = n43769 & ~n54725;
  assign n54751 = n52038 & ~n54725;
  assign n54752 = n52042 & ~n54725;
  assign n54753 = ~n54749 & ~n54750;
  assign n54754 = ~n54751 & n54753;
  assign n54755 = ~n54752 & n54754;
  assign n54756 = n43625 & ~n54733;
  assign n54757 = n43703 & ~n54733;
  assign n54758 = n43707 & ~n54733;
  assign n54759 = P1_P1_INSTADDRPOINTER_REG_30_ & n54677;
  assign n54760 = ~P1_P1_INSTADDRPOINTER_REG_31_ & n54759;
  assign n54761 = P1_P1_INSTADDRPOINTER_REG_31_ & ~n54759;
  assign n54762 = ~n54760 & ~n54761;
  assign n54763 = n43723 & ~n54762;
  assign n54764 = n43715 & ~n54762;
  assign n54765 = ~n54756 & ~n54757;
  assign n54766 = ~n54758 & n54765;
  assign n54767 = ~n54763 & n54766;
  assign n54768 = ~n54764 & n54767;
  assign n54769 = n54519 & n54743;
  assign n54770 = ~P1_P1_INSTADDRPOINTER_REG_31_ & n54769;
  assign n54771 = P1_P1_INSTADDRPOINTER_REG_31_ & ~n54769;
  assign n54772 = ~n54770 & ~n54771;
  assign n54773 = n43726 & ~n54772;
  assign n54774 = n54755 & n54768;
  assign n54775 = ~n54773 & n54774;
  assign n54776 = ~n54726 & n54729;
  assign n54777 = n54742 & n54776;
  assign n54778 = ~n54748 & n54777;
  assign n54779 = n54775 & n54778;
  assign n54780 = ~n54721 & n54779;
  assign n54781 = n51925 & ~n54780;
  assign n8951 = ~n54702 | n54781;
  assign n54783 = P1_P1_STATE2_REG_0_ & ~n43592;
  assign n54784 = ~P1_P1_STATE2_REG_0_ & ~n51892;
  assign n54785 = n43726 & n43729;
  assign n54786 = n43731 & n43735;
  assign n54787 = ~n54785 & ~n54786;
  assign n54788 = n43979 & ~n54787;
  assign n54789 = ~n54784 & ~n54788;
  assign n54790 = n54783 & ~n54789;
  assign n54791 = ~n52029 & n54790;
  assign n54792 = ~n51998 & n54791;
  assign n54793 = n52029 & n54790;
  assign n54794 = ~n51998 & n54793;
  assign n54795 = P1_P1_STATE2_REG_1_ & ~n54789;
  assign n54796 = P1_P1_STATEBS16_REG & n54795;
  assign n54797 = P1_P1_PHYADDRPOINTER_REG_0_ & n54796;
  assign n54798 = ~P1_P1_STATEBS16_REG & n54795;
  assign n54799 = P1_P1_PHYADDRPOINTER_REG_0_ & n54798;
  assign n54800 = P1_P1_PHYADDRPOINTER_REG_0_ & n54789;
  assign n54801 = P1_P1_STATE2_REG_0_ & n43592;
  assign n54802 = ~n54789 & n54801;
  assign n54803 = ~n52046 & n54802;
  assign n54804 = P1_P1_STATE2_REG_2_ & ~P1_P1_STATE2_REG_0_;
  assign n54805 = ~n54789 & n54804;
  assign n54806 = P1_P1_PHYADDRPOINTER_REG_0_ & n54805;
  assign n54807 = n43995 & ~n54789;
  assign n54808 = P1_P1_REIP_REG_0_ & n54807;
  assign n54809 = ~n54800 & ~n54803;
  assign n54810 = ~n54806 & n54809;
  assign n54811 = ~n54808 & n54810;
  assign n54812 = ~n54792 & ~n54794;
  assign n54813 = ~n54797 & n54812;
  assign n54814 = ~n54799 & n54813;
  assign n8956 = ~n54811 | ~n54814;
  assign n54816 = ~n52127 & n54791;
  assign n54817 = ~n52137 & n54793;
  assign n54818 = P1_P1_PHYADDRPOINTER_REG_1_ & n54796;
  assign n54819 = ~P1_P1_PHYADDRPOINTER_REG_1_ & n54798;
  assign n54820 = P1_P1_PHYADDRPOINTER_REG_1_ & n54789;
  assign n54821 = ~n52168 & n54802;
  assign n54822 = ~P1_P1_PHYADDRPOINTER_REG_1_ & n54805;
  assign n54823 = P1_P1_REIP_REG_1_ & n54807;
  assign n54824 = ~n54820 & ~n54821;
  assign n54825 = ~n54822 & n54824;
  assign n54826 = ~n54823 & n54825;
  assign n54827 = ~n54816 & ~n54817;
  assign n54828 = ~n54818 & n54827;
  assign n54829 = ~n54819 & n54828;
  assign n8961 = ~n54826 | ~n54829;
  assign n54831 = ~n52293 & n54791;
  assign n54832 = ~n52242 & n54793;
  assign n54833 = ~P1_P1_PHYADDRPOINTER_REG_2_ & n54796;
  assign n54834 = P1_P1_PHYADDRPOINTER_REG_1_ & ~P1_P1_PHYADDRPOINTER_REG_2_;
  assign n54835 = ~P1_P1_PHYADDRPOINTER_REG_1_ & P1_P1_PHYADDRPOINTER_REG_2_;
  assign n54836 = ~n54834 & ~n54835;
  assign n54837 = n54798 & ~n54836;
  assign n54838 = P1_P1_PHYADDRPOINTER_REG_2_ & n54789;
  assign n54839 = ~n52278 & n54802;
  assign n54840 = n54805 & ~n54836;
  assign n54841 = P1_P1_REIP_REG_2_ & n54807;
  assign n54842 = ~n54838 & ~n54839;
  assign n54843 = ~n54840 & n54842;
  assign n54844 = ~n54841 & n54843;
  assign n54845 = ~n54831 & ~n54832;
  assign n54846 = ~n54833 & n54845;
  assign n54847 = ~n54837 & n54846;
  assign n8966 = ~n54844 | ~n54847;
  assign n54849 = ~n52385 & n54791;
  assign n54850 = n52367 & n54793;
  assign n54851 = P1_P1_PHYADDRPOINTER_REG_2_ & ~P1_P1_PHYADDRPOINTER_REG_3_;
  assign n54852 = ~P1_P1_PHYADDRPOINTER_REG_2_ & P1_P1_PHYADDRPOINTER_REG_3_;
  assign n54853 = ~n54851 & ~n54852;
  assign n54854 = n54796 & ~n54853;
  assign n54855 = P1_P1_PHYADDRPOINTER_REG_1_ & P1_P1_PHYADDRPOINTER_REG_2_;
  assign n54856 = ~P1_P1_PHYADDRPOINTER_REG_3_ & n54855;
  assign n54857 = P1_P1_PHYADDRPOINTER_REG_3_ & ~n54855;
  assign n54858 = ~n54856 & ~n54857;
  assign n54859 = n54798 & ~n54858;
  assign n54860 = n54805 & ~n54858;
  assign n54861 = P1_P1_REIP_REG_3_ & n54807;
  assign n54862 = P1_P1_PHYADDRPOINTER_REG_3_ & n54789;
  assign n54863 = n52423 & n54802;
  assign n54864 = ~n54860 & ~n54861;
  assign n54865 = ~n54862 & n54864;
  assign n54866 = ~n54863 & n54865;
  assign n54867 = ~n54849 & ~n54850;
  assign n54868 = ~n54854 & n54867;
  assign n54869 = ~n54859 & n54868;
  assign n8971 = ~n54866 | ~n54869;
  assign n54871 = P1_P1_PHYADDRPOINTER_REG_2_ & P1_P1_PHYADDRPOINTER_REG_3_;
  assign n54872 = ~P1_P1_PHYADDRPOINTER_REG_4_ & n54871;
  assign n54873 = P1_P1_PHYADDRPOINTER_REG_4_ & ~n54871;
  assign n54874 = ~n54872 & ~n54873;
  assign n54875 = n54796 & ~n54874;
  assign n54876 = P1_P1_PHYADDRPOINTER_REG_3_ & n54855;
  assign n54877 = ~P1_P1_PHYADDRPOINTER_REG_4_ & n54876;
  assign n54878 = P1_P1_PHYADDRPOINTER_REG_4_ & ~n54876;
  assign n54879 = ~n54877 & ~n54878;
  assign n54880 = n54798 & ~n54879;
  assign n54881 = n52498 & n54793;
  assign n54882 = ~n52520 & n54791;
  assign n54883 = n54805 & ~n54879;
  assign n54884 = P1_P1_REIP_REG_4_ & n54807;
  assign n54885 = P1_P1_PHYADDRPOINTER_REG_4_ & n54789;
  assign n54886 = ~n52559 & n54802;
  assign n54887 = ~n54883 & ~n54884;
  assign n54888 = ~n54885 & n54887;
  assign n54889 = ~n54886 & n54888;
  assign n54890 = ~n54875 & ~n54880;
  assign n54891 = ~n54881 & n54890;
  assign n54892 = ~n54882 & n54891;
  assign n8976 = ~n54889 | ~n54892;
  assign n54894 = P1_P1_PHYADDRPOINTER_REG_4_ & n54871;
  assign n54895 = ~P1_P1_PHYADDRPOINTER_REG_5_ & n54894;
  assign n54896 = P1_P1_PHYADDRPOINTER_REG_5_ & ~n54894;
  assign n54897 = ~n54895 & ~n54896;
  assign n54898 = n54796 & ~n54897;
  assign n54899 = P1_P1_PHYADDRPOINTER_REG_4_ & n54876;
  assign n54900 = ~P1_P1_PHYADDRPOINTER_REG_5_ & n54899;
  assign n54901 = P1_P1_PHYADDRPOINTER_REG_5_ & ~n54899;
  assign n54902 = ~n54900 & ~n54901;
  assign n54903 = n54798 & ~n54902;
  assign n54904 = ~n52634 & n54793;
  assign n54905 = ~n52653 & n54791;
  assign n54906 = n54805 & ~n54902;
  assign n54907 = P1_P1_REIP_REG_5_ & n54807;
  assign n54908 = P1_P1_PHYADDRPOINTER_REG_5_ & n54789;
  assign n54909 = n52692 & n54802;
  assign n54910 = ~n54906 & ~n54907;
  assign n54911 = ~n54908 & n54910;
  assign n54912 = ~n54909 & n54911;
  assign n54913 = ~n54898 & ~n54903;
  assign n54914 = ~n54904 & n54913;
  assign n54915 = ~n54905 & n54914;
  assign n8981 = ~n54912 | ~n54915;
  assign n54917 = P1_P1_PHYADDRPOINTER_REG_5_ & n54894;
  assign n54918 = ~P1_P1_PHYADDRPOINTER_REG_6_ & n54917;
  assign n54919 = P1_P1_PHYADDRPOINTER_REG_6_ & ~n54917;
  assign n54920 = ~n54918 & ~n54919;
  assign n54921 = n54796 & ~n54920;
  assign n54922 = P1_P1_PHYADDRPOINTER_REG_5_ & n54899;
  assign n54923 = ~P1_P1_PHYADDRPOINTER_REG_6_ & n54922;
  assign n54924 = P1_P1_PHYADDRPOINTER_REG_6_ & ~n54922;
  assign n54925 = ~n54923 & ~n54924;
  assign n54926 = n54798 & ~n54925;
  assign n54927 = ~n52768 & n54793;
  assign n54928 = ~n52823 & n54791;
  assign n54929 = n54805 & ~n54925;
  assign n54930 = P1_P1_REIP_REG_6_ & n54807;
  assign n54931 = P1_P1_PHYADDRPOINTER_REG_6_ & n54789;
  assign n54932 = ~n52805 & n54802;
  assign n54933 = ~n54929 & ~n54930;
  assign n54934 = ~n54931 & n54933;
  assign n54935 = ~n54932 & n54934;
  assign n54936 = ~n54921 & ~n54926;
  assign n54937 = ~n54927 & n54936;
  assign n54938 = ~n54928 & n54937;
  assign n8986 = ~n54935 | ~n54938;
  assign n54940 = P1_P1_PHYADDRPOINTER_REG_6_ & n54917;
  assign n54941 = ~P1_P1_PHYADDRPOINTER_REG_7_ & n54940;
  assign n54942 = P1_P1_PHYADDRPOINTER_REG_7_ & ~n54940;
  assign n54943 = ~n54941 & ~n54942;
  assign n54944 = n54796 & ~n54943;
  assign n54945 = P1_P1_PHYADDRPOINTER_REG_6_ & n54922;
  assign n54946 = ~P1_P1_PHYADDRPOINTER_REG_7_ & n54945;
  assign n54947 = P1_P1_PHYADDRPOINTER_REG_7_ & ~n54945;
  assign n54948 = ~n54946 & ~n54947;
  assign n54949 = n54798 & ~n54948;
  assign n54950 = ~n52868 & n54793;
  assign n54951 = ~n52927 & n54791;
  assign n54952 = n54805 & ~n54948;
  assign n54953 = P1_P1_REIP_REG_7_ & n54807;
  assign n54954 = P1_P1_PHYADDRPOINTER_REG_7_ & n54789;
  assign n54955 = ~n52903 & n54802;
  assign n54956 = ~n54952 & ~n54953;
  assign n54957 = ~n54954 & n54956;
  assign n54958 = ~n54955 & n54957;
  assign n54959 = ~n54944 & ~n54949;
  assign n54960 = ~n54950 & n54959;
  assign n54961 = ~n54951 & n54960;
  assign n8991 = ~n54958 | ~n54961;
  assign n54963 = P1_P1_PHYADDRPOINTER_REG_7_ & n54940;
  assign n54964 = ~P1_P1_PHYADDRPOINTER_REG_8_ & n54963;
  assign n54965 = P1_P1_PHYADDRPOINTER_REG_8_ & ~n54963;
  assign n54966 = ~n54964 & ~n54965;
  assign n54967 = n54796 & ~n54966;
  assign n54968 = P1_P1_PHYADDRPOINTER_REG_7_ & n54945;
  assign n54969 = ~P1_P1_PHYADDRPOINTER_REG_8_ & n54968;
  assign n54970 = P1_P1_PHYADDRPOINTER_REG_8_ & ~n54968;
  assign n54971 = ~n54969 & ~n54970;
  assign n54972 = n54798 & ~n54971;
  assign n54973 = ~n52970 & n54793;
  assign n54974 = ~n53017 & n54791;
  assign n54975 = n54805 & ~n54971;
  assign n54976 = P1_P1_REIP_REG_8_ & n54807;
  assign n54977 = P1_P1_PHYADDRPOINTER_REG_8_ & n54789;
  assign n54978 = ~n53003 & n54802;
  assign n54979 = ~n54975 & ~n54976;
  assign n54980 = ~n54977 & n54979;
  assign n54981 = ~n54978 & n54980;
  assign n54982 = ~n54967 & ~n54972;
  assign n54983 = ~n54973 & n54982;
  assign n54984 = ~n54974 & n54983;
  assign n8996 = ~n54981 | ~n54984;
  assign n54986 = P1_P1_PHYADDRPOINTER_REG_8_ & n54963;
  assign n54987 = ~P1_P1_PHYADDRPOINTER_REG_9_ & n54986;
  assign n54988 = P1_P1_PHYADDRPOINTER_REG_9_ & ~n54986;
  assign n54989 = ~n54987 & ~n54988;
  assign n54990 = n54796 & ~n54989;
  assign n54991 = P1_P1_PHYADDRPOINTER_REG_8_ & n54968;
  assign n54992 = ~P1_P1_PHYADDRPOINTER_REG_9_ & n54991;
  assign n54993 = P1_P1_PHYADDRPOINTER_REG_9_ & ~n54991;
  assign n54994 = ~n54992 & ~n54993;
  assign n54995 = n54798 & ~n54994;
  assign n54996 = n53055 & n54793;
  assign n54997 = ~n53102 & n54791;
  assign n54998 = n54805 & ~n54994;
  assign n54999 = P1_P1_REIP_REG_9_ & n54807;
  assign n55000 = P1_P1_PHYADDRPOINTER_REG_9_ & n54789;
  assign n55001 = n53083 & n54802;
  assign n55002 = ~n54998 & ~n54999;
  assign n55003 = ~n55000 & n55002;
  assign n55004 = ~n55001 & n55003;
  assign n55005 = ~n54990 & ~n54995;
  assign n55006 = ~n54996 & n55005;
  assign n55007 = ~n54997 & n55006;
  assign n9001 = ~n55004 | ~n55007;
  assign n55009 = P1_P1_PHYADDRPOINTER_REG_9_ & n54986;
  assign n55010 = ~P1_P1_PHYADDRPOINTER_REG_10_ & n55009;
  assign n55011 = P1_P1_PHYADDRPOINTER_REG_10_ & ~n55009;
  assign n55012 = ~n55010 & ~n55011;
  assign n55013 = n54796 & ~n55012;
  assign n55014 = P1_P1_PHYADDRPOINTER_REG_9_ & n54991;
  assign n55015 = ~P1_P1_PHYADDRPOINTER_REG_10_ & n55014;
  assign n55016 = P1_P1_PHYADDRPOINTER_REG_10_ & ~n55014;
  assign n55017 = ~n55015 & ~n55016;
  assign n55018 = n54798 & ~n55017;
  assign n55019 = n53135 & n54793;
  assign n55020 = ~n53178 & n54791;
  assign n55021 = n54805 & ~n55017;
  assign n55022 = P1_P1_REIP_REG_10_ & n54807;
  assign n55023 = P1_P1_PHYADDRPOINTER_REG_10_ & n54789;
  assign n55024 = n53159 & n54802;
  assign n55025 = ~n55021 & ~n55022;
  assign n55026 = ~n55023 & n55025;
  assign n55027 = ~n55024 & n55026;
  assign n55028 = ~n55013 & ~n55018;
  assign n55029 = ~n55019 & n55028;
  assign n55030 = ~n55020 & n55029;
  assign n9006 = ~n55027 | ~n55030;
  assign n55032 = P1_P1_PHYADDRPOINTER_REG_10_ & n55009;
  assign n55033 = ~P1_P1_PHYADDRPOINTER_REG_11_ & n55032;
  assign n55034 = P1_P1_PHYADDRPOINTER_REG_11_ & ~n55032;
  assign n55035 = ~n55033 & ~n55034;
  assign n55036 = n54796 & ~n55035;
  assign n55037 = P1_P1_PHYADDRPOINTER_REG_10_ & n55014;
  assign n55038 = ~P1_P1_PHYADDRPOINTER_REG_11_ & n55037;
  assign n55039 = P1_P1_PHYADDRPOINTER_REG_11_ & ~n55037;
  assign n55040 = ~n55038 & ~n55039;
  assign n55041 = n54798 & ~n55040;
  assign n55042 = ~n53210 & n54793;
  assign n55043 = ~n53250 & n54791;
  assign n55044 = n54805 & ~n55040;
  assign n55045 = P1_P1_REIP_REG_11_ & n54807;
  assign n55046 = P1_P1_PHYADDRPOINTER_REG_11_ & n54789;
  assign n55047 = ~n53234 & n54802;
  assign n55048 = ~n55044 & ~n55045;
  assign n55049 = ~n55046 & n55048;
  assign n55050 = ~n55047 & n55049;
  assign n55051 = ~n55036 & ~n55041;
  assign n55052 = ~n55042 & n55051;
  assign n55053 = ~n55043 & n55052;
  assign n9011 = ~n55050 | ~n55053;
  assign n55055 = P1_P1_PHYADDRPOINTER_REG_11_ & n55032;
  assign n55056 = ~P1_P1_PHYADDRPOINTER_REG_12_ & n55055;
  assign n55057 = P1_P1_PHYADDRPOINTER_REG_12_ & ~n55055;
  assign n55058 = ~n55056 & ~n55057;
  assign n55059 = n54796 & ~n55058;
  assign n55060 = P1_P1_PHYADDRPOINTER_REG_11_ & n55037;
  assign n55061 = ~P1_P1_PHYADDRPOINTER_REG_12_ & n55060;
  assign n55062 = P1_P1_PHYADDRPOINTER_REG_12_ & ~n55060;
  assign n55063 = ~n55061 & ~n55062;
  assign n55064 = n54798 & ~n55063;
  assign n55065 = n53285 & n54793;
  assign n55066 = ~n53329 & n54791;
  assign n55067 = n54805 & ~n55063;
  assign n55068 = P1_P1_REIP_REG_12_ & n54807;
  assign n55069 = P1_P1_PHYADDRPOINTER_REG_12_ & n54789;
  assign n55070 = n53310 & n54802;
  assign n55071 = ~n55067 & ~n55068;
  assign n55072 = ~n55069 & n55071;
  assign n55073 = ~n55070 & n55072;
  assign n55074 = ~n55059 & ~n55064;
  assign n55075 = ~n55065 & n55074;
  assign n55076 = ~n55066 & n55075;
  assign n9016 = ~n55073 | ~n55076;
  assign n55078 = P1_P1_PHYADDRPOINTER_REG_12_ & n55055;
  assign n55079 = ~P1_P1_PHYADDRPOINTER_REG_13_ & n55078;
  assign n55080 = P1_P1_PHYADDRPOINTER_REG_13_ & ~n55078;
  assign n55081 = ~n55079 & ~n55080;
  assign n55082 = n54796 & ~n55081;
  assign n55083 = P1_P1_PHYADDRPOINTER_REG_12_ & n55060;
  assign n55084 = ~P1_P1_PHYADDRPOINTER_REG_13_ & n55083;
  assign n55085 = P1_P1_PHYADDRPOINTER_REG_13_ & ~n55083;
  assign n55086 = ~n55084 & ~n55085;
  assign n55087 = n54798 & ~n55086;
  assign n55088 = n53351 & n54793;
  assign n55089 = n53402 & n54791;
  assign n55090 = n54805 & ~n55086;
  assign n55091 = P1_P1_REIP_REG_13_ & n54807;
  assign n55092 = P1_P1_PHYADDRPOINTER_REG_13_ & n54789;
  assign n55093 = n53379 & n54802;
  assign n55094 = ~n55090 & ~n55091;
  assign n55095 = ~n55092 & n55094;
  assign n55096 = ~n55093 & n55095;
  assign n55097 = ~n55082 & ~n55087;
  assign n55098 = ~n55088 & n55097;
  assign n55099 = ~n55089 & n55098;
  assign n9021 = ~n55096 | ~n55099;
  assign n55101 = P1_P1_PHYADDRPOINTER_REG_13_ & n55078;
  assign n55102 = ~P1_P1_PHYADDRPOINTER_REG_14_ & n55101;
  assign n55103 = P1_P1_PHYADDRPOINTER_REG_14_ & ~n55101;
  assign n55104 = ~n55102 & ~n55103;
  assign n55105 = n54796 & ~n55104;
  assign n55106 = P1_P1_PHYADDRPOINTER_REG_13_ & n55083;
  assign n55107 = ~P1_P1_PHYADDRPOINTER_REG_14_ & n55106;
  assign n55108 = P1_P1_PHYADDRPOINTER_REG_14_ & ~n55106;
  assign n55109 = ~n55107 & ~n55108;
  assign n55110 = n54798 & ~n55109;
  assign n55111 = ~n53436 & n54793;
  assign n55112 = ~n53477 & n54791;
  assign n55113 = n54805 & ~n55109;
  assign n55114 = P1_P1_REIP_REG_14_ & n54807;
  assign n55115 = P1_P1_PHYADDRPOINTER_REG_14_ & n54789;
  assign n55116 = ~n53460 & n54802;
  assign n55117 = ~n55113 & ~n55114;
  assign n55118 = ~n55115 & n55117;
  assign n55119 = ~n55116 & n55118;
  assign n55120 = ~n55105 & ~n55110;
  assign n55121 = ~n55111 & n55120;
  assign n55122 = ~n55112 & n55121;
  assign n9026 = ~n55119 | ~n55122;
  assign n55124 = P1_P1_PHYADDRPOINTER_REG_14_ & n55101;
  assign n55125 = ~P1_P1_PHYADDRPOINTER_REG_15_ & n55124;
  assign n55126 = P1_P1_PHYADDRPOINTER_REG_15_ & ~n55124;
  assign n55127 = ~n55125 & ~n55126;
  assign n55128 = n54796 & ~n55127;
  assign n55129 = P1_P1_PHYADDRPOINTER_REG_14_ & n55106;
  assign n55130 = ~P1_P1_PHYADDRPOINTER_REG_15_ & n55129;
  assign n55131 = P1_P1_PHYADDRPOINTER_REG_15_ & ~n55129;
  assign n55132 = ~n55130 & ~n55131;
  assign n55133 = n54798 & ~n55132;
  assign n55134 = n53502 & n54793;
  assign n55135 = ~n53552 & n54791;
  assign n55136 = n54805 & ~n55132;
  assign n55137 = P1_P1_REIP_REG_15_ & n54807;
  assign n55138 = P1_P1_PHYADDRPOINTER_REG_15_ & n54789;
  assign n55139 = n53531 & n54802;
  assign n55140 = ~n55136 & ~n55137;
  assign n55141 = ~n55138 & n55140;
  assign n55142 = ~n55139 & n55141;
  assign n55143 = ~n55128 & ~n55133;
  assign n55144 = ~n55134 & n55143;
  assign n55145 = ~n55135 & n55144;
  assign n9031 = ~n55142 | ~n55145;
  assign n55147 = P1_P1_PHYADDRPOINTER_REG_15_ & n55124;
  assign n55148 = ~P1_P1_PHYADDRPOINTER_REG_16_ & n55147;
  assign n55149 = P1_P1_PHYADDRPOINTER_REG_16_ & ~n55147;
  assign n55150 = ~n55148 & ~n55149;
  assign n55151 = n54796 & ~n55150;
  assign n55152 = P1_P1_PHYADDRPOINTER_REG_15_ & n55129;
  assign n55153 = ~P1_P1_PHYADDRPOINTER_REG_16_ & n55152;
  assign n55154 = P1_P1_PHYADDRPOINTER_REG_16_ & ~n55152;
  assign n55155 = ~n55153 & ~n55154;
  assign n55156 = n54798 & ~n55155;
  assign n55157 = ~n53577 & n54793;
  assign n55158 = ~n53624 & n54791;
  assign n55159 = n54805 & ~n55155;
  assign n55160 = P1_P1_REIP_REG_16_ & n54807;
  assign n55161 = P1_P1_PHYADDRPOINTER_REG_16_ & n54789;
  assign n55162 = ~n53605 & n54802;
  assign n55163 = ~n55159 & ~n55160;
  assign n55164 = ~n55161 & n55163;
  assign n55165 = ~n55162 & n55164;
  assign n55166 = ~n55151 & ~n55156;
  assign n55167 = ~n55157 & n55166;
  assign n55168 = ~n55158 & n55167;
  assign n9036 = ~n55165 | ~n55168;
  assign n55170 = P1_P1_PHYADDRPOINTER_REG_16_ & n55147;
  assign n55171 = ~P1_P1_PHYADDRPOINTER_REG_17_ & n55170;
  assign n55172 = P1_P1_PHYADDRPOINTER_REG_17_ & ~n55170;
  assign n55173 = ~n55171 & ~n55172;
  assign n55174 = n54796 & ~n55173;
  assign n55175 = P1_P1_PHYADDRPOINTER_REG_16_ & n55152;
  assign n55176 = ~P1_P1_PHYADDRPOINTER_REG_17_ & n55175;
  assign n55177 = P1_P1_PHYADDRPOINTER_REG_17_ & ~n55175;
  assign n55178 = ~n55176 & ~n55177;
  assign n55179 = n54798 & ~n55178;
  assign n55180 = n53651 & n54793;
  assign n55181 = n53703 & n54791;
  assign n55182 = n54805 & ~n55178;
  assign n55183 = P1_P1_REIP_REG_17_ & n54807;
  assign n55184 = P1_P1_PHYADDRPOINTER_REG_17_ & n54789;
  assign n55185 = n53680 & n54802;
  assign n55186 = ~n55182 & ~n55183;
  assign n55187 = ~n55184 & n55186;
  assign n55188 = ~n55185 & n55187;
  assign n55189 = ~n55174 & ~n55179;
  assign n55190 = ~n55180 & n55189;
  assign n55191 = ~n55181 & n55190;
  assign n9041 = ~n55188 | ~n55191;
  assign n55193 = P1_P1_PHYADDRPOINTER_REG_17_ & n55170;
  assign n55194 = ~P1_P1_PHYADDRPOINTER_REG_18_ & n55193;
  assign n55195 = P1_P1_PHYADDRPOINTER_REG_18_ & ~n55193;
  assign n55196 = ~n55194 & ~n55195;
  assign n55197 = n54796 & ~n55196;
  assign n55198 = P1_P1_PHYADDRPOINTER_REG_17_ & n55175;
  assign n55199 = ~P1_P1_PHYADDRPOINTER_REG_18_ & n55198;
  assign n55200 = P1_P1_PHYADDRPOINTER_REG_18_ & ~n55198;
  assign n55201 = ~n55199 & ~n55200;
  assign n55202 = n54798 & ~n55201;
  assign n55203 = ~n53728 & n54793;
  assign n55204 = ~n53774 & n54791;
  assign n55205 = n54805 & ~n55201;
  assign n55206 = P1_P1_REIP_REG_18_ & n54807;
  assign n55207 = P1_P1_PHYADDRPOINTER_REG_18_ & n54789;
  assign n55208 = ~n53756 & n54802;
  assign n55209 = ~n55205 & ~n55206;
  assign n55210 = ~n55207 & n55209;
  assign n55211 = ~n55208 & n55210;
  assign n55212 = ~n55197 & ~n55202;
  assign n55213 = ~n55203 & n55212;
  assign n55214 = ~n55204 & n55213;
  assign n9046 = ~n55211 | ~n55214;
  assign n55216 = P1_P1_PHYADDRPOINTER_REG_18_ & n55193;
  assign n55217 = ~P1_P1_PHYADDRPOINTER_REG_19_ & n55216;
  assign n55218 = P1_P1_PHYADDRPOINTER_REG_19_ & ~n55216;
  assign n55219 = ~n55217 & ~n55218;
  assign n55220 = n54796 & ~n55219;
  assign n55221 = P1_P1_PHYADDRPOINTER_REG_18_ & n55198;
  assign n55222 = ~P1_P1_PHYADDRPOINTER_REG_19_ & n55221;
  assign n55223 = P1_P1_PHYADDRPOINTER_REG_19_ & ~n55221;
  assign n55224 = ~n55222 & ~n55223;
  assign n55225 = n54798 & ~n55224;
  assign n55226 = n53803 & n54793;
  assign n55227 = ~n53854 & n54791;
  assign n55228 = n54805 & ~n55224;
  assign n55229 = P1_P1_REIP_REG_19_ & n54807;
  assign n55230 = P1_P1_PHYADDRPOINTER_REG_19_ & n54789;
  assign n55231 = n53832 & n54802;
  assign n55232 = ~n55228 & ~n55229;
  assign n55233 = ~n55230 & n55232;
  assign n55234 = ~n55231 & n55233;
  assign n55235 = ~n55220 & ~n55225;
  assign n55236 = ~n55226 & n55235;
  assign n55237 = ~n55227 & n55236;
  assign n9051 = ~n55234 | ~n55237;
  assign n55239 = P1_P1_PHYADDRPOINTER_REG_19_ & n55216;
  assign n55240 = ~P1_P1_PHYADDRPOINTER_REG_20_ & n55239;
  assign n55241 = P1_P1_PHYADDRPOINTER_REG_20_ & ~n55239;
  assign n55242 = ~n55240 & ~n55241;
  assign n55243 = n54796 & ~n55242;
  assign n55244 = P1_P1_PHYADDRPOINTER_REG_19_ & n55221;
  assign n55245 = ~P1_P1_PHYADDRPOINTER_REG_20_ & n55244;
  assign n55246 = P1_P1_PHYADDRPOINTER_REG_20_ & ~n55244;
  assign n55247 = ~n55245 & ~n55246;
  assign n55248 = n54798 & ~n55247;
  assign n55249 = n53879 & n54793;
  assign n55250 = n53930 & n54791;
  assign n55251 = n54805 & ~n55247;
  assign n55252 = P1_P1_REIP_REG_20_ & n54807;
  assign n55253 = P1_P1_PHYADDRPOINTER_REG_20_ & n54789;
  assign n55254 = n53907 & n54802;
  assign n55255 = ~n55251 & ~n55252;
  assign n55256 = ~n55253 & n55255;
  assign n55257 = ~n55254 & n55256;
  assign n55258 = ~n55243 & ~n55248;
  assign n55259 = ~n55249 & n55258;
  assign n55260 = ~n55250 & n55259;
  assign n9056 = ~n55257 | ~n55260;
  assign n55262 = P1_P1_PHYADDRPOINTER_REG_20_ & n55239;
  assign n55263 = ~P1_P1_PHYADDRPOINTER_REG_21_ & n55262;
  assign n55264 = P1_P1_PHYADDRPOINTER_REG_21_ & ~n55262;
  assign n55265 = ~n55263 & ~n55264;
  assign n55266 = n54796 & ~n55265;
  assign n55267 = P1_P1_PHYADDRPOINTER_REG_20_ & n55244;
  assign n55268 = ~P1_P1_PHYADDRPOINTER_REG_21_ & n55267;
  assign n55269 = P1_P1_PHYADDRPOINTER_REG_21_ & ~n55267;
  assign n55270 = ~n55268 & ~n55269;
  assign n55271 = n54798 & ~n55270;
  assign n55272 = n53956 & n54793;
  assign n55273 = ~n54003 & n54791;
  assign n55274 = P1_P1_PHYADDRPOINTER_REG_21_ & n54789;
  assign n55275 = P1_P1_REIP_REG_21_ & n54807;
  assign n55276 = n54805 & ~n55270;
  assign n55277 = n53984 & n54802;
  assign n55278 = ~n55274 & ~n55275;
  assign n55279 = ~n55276 & n55278;
  assign n55280 = ~n55277 & n55279;
  assign n55281 = ~n55266 & ~n55271;
  assign n55282 = ~n55272 & n55281;
  assign n55283 = ~n55273 & n55282;
  assign n9061 = ~n55280 | ~n55283;
  assign n55285 = P1_P1_PHYADDRPOINTER_REG_21_ & n55262;
  assign n55286 = ~P1_P1_PHYADDRPOINTER_REG_22_ & n55285;
  assign n55287 = P1_P1_PHYADDRPOINTER_REG_22_ & ~n55285;
  assign n55288 = ~n55286 & ~n55287;
  assign n55289 = n54796 & ~n55288;
  assign n55290 = P1_P1_PHYADDRPOINTER_REG_21_ & n55267;
  assign n55291 = ~P1_P1_PHYADDRPOINTER_REG_22_ & n55290;
  assign n55292 = P1_P1_PHYADDRPOINTER_REG_22_ & ~n55290;
  assign n55293 = ~n55291 & ~n55292;
  assign n55294 = n54798 & ~n55293;
  assign n55295 = ~n54028 & n54793;
  assign n55296 = ~n54080 & n54791;
  assign n55297 = P1_P1_PHYADDRPOINTER_REG_22_ & n54789;
  assign n55298 = P1_P1_REIP_REG_22_ & n54807;
  assign n55299 = n54805 & ~n55293;
  assign n55300 = ~n54056 & n54802;
  assign n55301 = ~n55297 & ~n55298;
  assign n55302 = ~n55299 & n55301;
  assign n55303 = ~n55300 & n55302;
  assign n55304 = ~n55289 & ~n55294;
  assign n55305 = ~n55295 & n55304;
  assign n55306 = ~n55296 & n55305;
  assign n9066 = ~n55303 | ~n55306;
  assign n55308 = P1_P1_PHYADDRPOINTER_REG_22_ & n55285;
  assign n55309 = ~P1_P1_PHYADDRPOINTER_REG_23_ & n55308;
  assign n55310 = P1_P1_PHYADDRPOINTER_REG_23_ & ~n55308;
  assign n55311 = ~n55309 & ~n55310;
  assign n55312 = n54796 & ~n55311;
  assign n55313 = P1_P1_PHYADDRPOINTER_REG_22_ & n55290;
  assign n55314 = ~P1_P1_PHYADDRPOINTER_REG_23_ & n55313;
  assign n55315 = P1_P1_PHYADDRPOINTER_REG_23_ & ~n55313;
  assign n55316 = ~n55314 & ~n55315;
  assign n55317 = n54798 & ~n55316;
  assign n55318 = n54107 & n54793;
  assign n55319 = ~n54159 & n54791;
  assign n55320 = P1_P1_PHYADDRPOINTER_REG_23_ & n54789;
  assign n55321 = P1_P1_REIP_REG_23_ & n54807;
  assign n55322 = n54805 & ~n55316;
  assign n55323 = n54138 & n54802;
  assign n55324 = ~n55320 & ~n55321;
  assign n55325 = ~n55322 & n55324;
  assign n55326 = ~n55323 & n55325;
  assign n55327 = ~n55312 & ~n55317;
  assign n55328 = ~n55318 & n55327;
  assign n55329 = ~n55319 & n55328;
  assign n9071 = ~n55326 | ~n55329;
  assign n55331 = P1_P1_PHYADDRPOINTER_REG_23_ & n55308;
  assign n55332 = ~P1_P1_PHYADDRPOINTER_REG_24_ & n55331;
  assign n55333 = P1_P1_PHYADDRPOINTER_REG_24_ & ~n55331;
  assign n55334 = ~n55332 & ~n55333;
  assign n55335 = n54796 & ~n55334;
  assign n55336 = P1_P1_PHYADDRPOINTER_REG_23_ & n55313;
  assign n55337 = ~P1_P1_PHYADDRPOINTER_REG_24_ & n55336;
  assign n55338 = P1_P1_PHYADDRPOINTER_REG_24_ & ~n55336;
  assign n55339 = ~n55337 & ~n55338;
  assign n55340 = n54798 & ~n55339;
  assign n55341 = ~n54184 & n54793;
  assign n55342 = ~n54233 & n54791;
  assign n55343 = P1_P1_PHYADDRPOINTER_REG_24_ & n54789;
  assign n55344 = P1_P1_REIP_REG_24_ & n54807;
  assign n55345 = n54805 & ~n55339;
  assign n55346 = ~n54212 & n54802;
  assign n55347 = ~n55343 & ~n55344;
  assign n55348 = ~n55345 & n55347;
  assign n55349 = ~n55346 & n55348;
  assign n55350 = ~n55335 & ~n55340;
  assign n55351 = ~n55341 & n55350;
  assign n55352 = ~n55342 & n55351;
  assign n9076 = ~n55349 | ~n55352;
  assign n55354 = P1_P1_PHYADDRPOINTER_REG_24_ & n55331;
  assign n55355 = ~P1_P1_PHYADDRPOINTER_REG_25_ & n55354;
  assign n55356 = P1_P1_PHYADDRPOINTER_REG_25_ & ~n55354;
  assign n55357 = ~n55355 & ~n55356;
  assign n55358 = n54796 & ~n55357;
  assign n55359 = P1_P1_PHYADDRPOINTER_REG_24_ & n55336;
  assign n55360 = ~P1_P1_PHYADDRPOINTER_REG_25_ & n55359;
  assign n55361 = P1_P1_PHYADDRPOINTER_REG_25_ & ~n55359;
  assign n55362 = ~n55360 & ~n55361;
  assign n55363 = n54798 & ~n55362;
  assign n55364 = n54260 & n54793;
  assign n55365 = P1_P1_PHYADDRPOINTER_REG_25_ & n54789;
  assign n55366 = P1_P1_REIP_REG_25_ & n54807;
  assign n55367 = n54805 & ~n55362;
  assign n55368 = n54289 & n54802;
  assign n55369 = ~n55365 & ~n55366;
  assign n55370 = ~n55367 & n55369;
  assign n55371 = ~n55368 & n55370;
  assign n55372 = ~n54313 & n54791;
  assign n55373 = ~n55358 & ~n55363;
  assign n55374 = ~n55364 & n55373;
  assign n55375 = n55371 & n55374;
  assign n9081 = n55372 | ~n55375;
  assign n55377 = P1_P1_PHYADDRPOINTER_REG_25_ & n55354;
  assign n55378 = ~P1_P1_PHYADDRPOINTER_REG_26_ & n55377;
  assign n55379 = P1_P1_PHYADDRPOINTER_REG_26_ & ~n55377;
  assign n55380 = ~n55378 & ~n55379;
  assign n55381 = n54796 & ~n55380;
  assign n55382 = P1_P1_PHYADDRPOINTER_REG_25_ & n55359;
  assign n55383 = ~P1_P1_PHYADDRPOINTER_REG_26_ & n55382;
  assign n55384 = P1_P1_PHYADDRPOINTER_REG_26_ & ~n55382;
  assign n55385 = ~n55383 & ~n55384;
  assign n55386 = n54798 & ~n55385;
  assign n55387 = n54338 & n54793;
  assign n55388 = P1_P1_PHYADDRPOINTER_REG_26_ & n54789;
  assign n55389 = P1_P1_REIP_REG_26_ & n54807;
  assign n55390 = n54805 & ~n55385;
  assign n55391 = n54366 & n54802;
  assign n55392 = ~n55388 & ~n55389;
  assign n55393 = ~n55390 & n55392;
  assign n55394 = ~n55391 & n55393;
  assign n55395 = n54388 & n54791;
  assign n55396 = ~n55381 & ~n55386;
  assign n55397 = ~n55387 & n55396;
  assign n55398 = n55394 & n55397;
  assign n9086 = n55395 | ~n55398;
  assign n55400 = P1_P1_PHYADDRPOINTER_REG_26_ & n55377;
  assign n55401 = ~P1_P1_PHYADDRPOINTER_REG_27_ & n55400;
  assign n55402 = P1_P1_PHYADDRPOINTER_REG_27_ & ~n55400;
  assign n55403 = ~n55401 & ~n55402;
  assign n55404 = n54796 & ~n55403;
  assign n55405 = P1_P1_PHYADDRPOINTER_REG_26_ & n55382;
  assign n55406 = ~P1_P1_PHYADDRPOINTER_REG_27_ & n55405;
  assign n55407 = P1_P1_PHYADDRPOINTER_REG_27_ & ~n55405;
  assign n55408 = ~n55406 & ~n55407;
  assign n55409 = n54798 & ~n55408;
  assign n55410 = ~n54413 & n54793;
  assign n55411 = P1_P1_PHYADDRPOINTER_REG_27_ & n54789;
  assign n55412 = P1_P1_REIP_REG_27_ & n54807;
  assign n55413 = n54805 & ~n55408;
  assign n55414 = ~n54441 & n54802;
  assign n55415 = ~n55411 & ~n55412;
  assign n55416 = ~n55413 & n55415;
  assign n55417 = ~n55414 & n55416;
  assign n55418 = ~n54459 & n54791;
  assign n55419 = ~n55404 & ~n55409;
  assign n55420 = ~n55410 & n55419;
  assign n55421 = n55417 & n55420;
  assign n9091 = n55418 | ~n55421;
  assign n55423 = P1_P1_PHYADDRPOINTER_REG_27_ & n55400;
  assign n55424 = ~P1_P1_PHYADDRPOINTER_REG_28_ & n55423;
  assign n55425 = P1_P1_PHYADDRPOINTER_REG_28_ & ~n55423;
  assign n55426 = ~n55424 & ~n55425;
  assign n55427 = n54796 & ~n55426;
  assign n55428 = P1_P1_PHYADDRPOINTER_REG_27_ & n55405;
  assign n55429 = ~P1_P1_PHYADDRPOINTER_REG_28_ & n55428;
  assign n55430 = P1_P1_PHYADDRPOINTER_REG_28_ & ~n55428;
  assign n55431 = ~n55429 & ~n55430;
  assign n55432 = n54798 & ~n55431;
  assign n55433 = n54487 & n54793;
  assign n55434 = P1_P1_PHYADDRPOINTER_REG_28_ & n54789;
  assign n55435 = P1_P1_REIP_REG_28_ & n54807;
  assign n55436 = n54805 & ~n55431;
  assign n55437 = n54520 & n54802;
  assign n55438 = ~n55434 & ~n55435;
  assign n55439 = ~n55436 & n55438;
  assign n55440 = ~n55437 & n55439;
  assign n55441 = n54544 & n54791;
  assign n55442 = ~n55427 & ~n55432;
  assign n55443 = ~n55433 & n55442;
  assign n55444 = n55440 & n55443;
  assign n9096 = n55441 | ~n55444;
  assign n55446 = P1_P1_PHYADDRPOINTER_REG_28_ & n55423;
  assign n55447 = ~P1_P1_PHYADDRPOINTER_REG_29_ & n55446;
  assign n55448 = P1_P1_PHYADDRPOINTER_REG_29_ & ~n55446;
  assign n55449 = ~n55447 & ~n55448;
  assign n55450 = n54796 & ~n55449;
  assign n55451 = P1_P1_PHYADDRPOINTER_REG_28_ & n55428;
  assign n55452 = ~P1_P1_PHYADDRPOINTER_REG_29_ & n55451;
  assign n55453 = P1_P1_PHYADDRPOINTER_REG_29_ & ~n55451;
  assign n55454 = ~n55452 & ~n55453;
  assign n55455 = n54798 & ~n55454;
  assign n55456 = n54593 & n54793;
  assign n55457 = P1_P1_PHYADDRPOINTER_REG_29_ & n54789;
  assign n55458 = P1_P1_REIP_REG_29_ & n54807;
  assign n55459 = n54805 & ~n55454;
  assign n55460 = n54617 & n54802;
  assign n55461 = ~n55457 & ~n55458;
  assign n55462 = ~n55459 & n55461;
  assign n55463 = ~n55460 & n55462;
  assign n55464 = ~n54568 & n54791;
  assign n55465 = ~n55450 & ~n55455;
  assign n55466 = ~n55456 & n55465;
  assign n55467 = n55463 & n55466;
  assign n9101 = n55464 | ~n55467;
  assign n55469 = P1_P1_PHYADDRPOINTER_REG_29_ & n55446;
  assign n55470 = ~P1_P1_PHYADDRPOINTER_REG_30_ & n55469;
  assign n55471 = P1_P1_PHYADDRPOINTER_REG_30_ & ~n55469;
  assign n55472 = ~n55470 & ~n55471;
  assign n55473 = n54796 & ~n55472;
  assign n55474 = P1_P1_PHYADDRPOINTER_REG_29_ & n55451;
  assign n55475 = ~P1_P1_PHYADDRPOINTER_REG_30_ & n55474;
  assign n55476 = P1_P1_PHYADDRPOINTER_REG_30_ & ~n55474;
  assign n55477 = ~n55475 & ~n55476;
  assign n55478 = n54798 & ~n55477;
  assign n55479 = ~n54665 & n54793;
  assign n55480 = P1_P1_PHYADDRPOINTER_REG_30_ & n54789;
  assign n55481 = P1_P1_REIP_REG_30_ & n54807;
  assign n55482 = n54805 & ~n55477;
  assign n55483 = ~n54689 & n54802;
  assign n55484 = ~n55480 & ~n55481;
  assign n55485 = ~n55482 & n55484;
  assign n55486 = ~n55483 & n55485;
  assign n55487 = ~n54640 & n54791;
  assign n55488 = ~n55473 & ~n55478;
  assign n55489 = ~n55479 & n55488;
  assign n55490 = n55486 & n55489;
  assign n9106 = n55487 | ~n55490;
  assign n55492 = P1_P1_PHYADDRPOINTER_REG_30_ & n55469;
  assign n55493 = ~P1_P1_PHYADDRPOINTER_REG_31_ & n55492;
  assign n55494 = P1_P1_PHYADDRPOINTER_REG_31_ & ~n55492;
  assign n55495 = ~n55493 & ~n55494;
  assign n55496 = n54796 & ~n55495;
  assign n55497 = P1_P1_PHYADDRPOINTER_REG_30_ & n55474;
  assign n55498 = ~P1_P1_PHYADDRPOINTER_REG_31_ & n55497;
  assign n55499 = P1_P1_PHYADDRPOINTER_REG_31_ & ~n55497;
  assign n55500 = ~n55498 & ~n55499;
  assign n55501 = n54798 & ~n55500;
  assign n55502 = ~n54747 & n54793;
  assign n55503 = P1_P1_PHYADDRPOINTER_REG_31_ & n54789;
  assign n55504 = P1_P1_REIP_REG_31_ & n54807;
  assign n55505 = n54805 & ~n55500;
  assign n55506 = ~n54772 & n54802;
  assign n55507 = ~n55503 & ~n55504;
  assign n55508 = ~n55505 & n55507;
  assign n55509 = ~n55506 & n55508;
  assign n55510 = n54720 & n54791;
  assign n55511 = ~n55496 & ~n55501;
  assign n55512 = ~n55502 & n55511;
  assign n55513 = n55509 & n55512;
  assign n9111 = n55510 | ~n55513;
  assign n55515 = ~n43251 & n43707;
  assign n55516 = n43676 & n55515;
  assign n55517 = ~n43863 & ~n55516;
  assign n55518 = n43979 & ~n55517;
  assign n55519 = P1_P1_LWORD_REG_15_ & ~n55518;
  assign n55520 = n43592 & n55518;
  assign n55521 = P1_P1_EAX_REG_15_ & n55520;
  assign n55522 = P1_BUF1_REG_15_ & n12460;
  assign n55523 = ~n47110 & ~n47114;
  assign n55524 = n47110 & n47114;
  assign n55525 = ~n55523 & ~n55524;
  assign n55526 = n47200 & ~n55525;
  assign n55527 = ~n47115 & ~n47116;
  assign n55528 = ~n47200 & ~n55527;
  assign n55529 = ~n55526 & ~n55528;
  assign n55530 = ~n12460 & ~n55529;
  assign n55531 = ~n55522 & ~n55530;
  assign n55532 = ~n43592 & n55518;
  assign n55533 = ~n55531 & n55532;
  assign n55534 = ~n55519 & ~n55521;
  assign n9116 = n55533 | ~n55534;
  assign n55536 = P1_P1_LWORD_REG_14_ & ~n55518;
  assign n55537 = P1_P1_EAX_REG_14_ & n55520;
  assign n55538 = P1_BUF1_REG_14_ & n12460;
  assign n55539 = n47125 & ~n47198;
  assign n55540 = ~n47125 & n47198;
  assign n55541 = ~n55539 & ~n55540;
  assign n55542 = ~n47124 & n55541;
  assign n55543 = n47124 & n55540;
  assign n55544 = n47126 & ~n47198;
  assign n55545 = ~n55542 & ~n55543;
  assign n55546 = ~n55544 & n55545;
  assign n55547 = ~n12460 & ~n55546;
  assign n55548 = ~n55538 & ~n55547;
  assign n55549 = n55532 & ~n55548;
  assign n55550 = ~n55536 & ~n55537;
  assign n9121 = n55549 | ~n55550;
  assign n55552 = P1_P1_LWORD_REG_13_ & ~n55518;
  assign n55553 = P1_P1_EAX_REG_13_ & n55520;
  assign n55554 = P1_BUF1_REG_13_ & n12460;
  assign n55555 = ~n47128 & ~n47135;
  assign n55556 = n47128 & n47135;
  assign n55557 = ~n55555 & ~n55556;
  assign n55558 = n47196 & ~n55557;
  assign n55559 = ~n47196 & n55557;
  assign n55560 = ~n55558 & ~n55559;
  assign n55561 = ~n12460 & ~n55560;
  assign n55562 = ~n55554 & ~n55561;
  assign n55563 = n55532 & ~n55562;
  assign n55564 = ~n55552 & ~n55553;
  assign n9126 = n55563 | ~n55564;
  assign n55566 = P1_P1_LWORD_REG_12_ & ~n55518;
  assign n55567 = P1_P1_EAX_REG_12_ & n55520;
  assign n55568 = P1_BUF1_REG_12_ & n12460;
  assign n55569 = ~n47138 & n47194;
  assign n55570 = n47144 & n55569;
  assign n55571 = n47138 & ~n47194;
  assign n55572 = ~n55569 & ~n55571;
  assign n55573 = ~n47144 & n55572;
  assign n55574 = n47145 & ~n47194;
  assign n55575 = ~n55570 & ~n55573;
  assign n55576 = ~n55574 & n55575;
  assign n55577 = ~n12460 & ~n55576;
  assign n55578 = ~n55568 & ~n55577;
  assign n55579 = n55532 & ~n55578;
  assign n55580 = ~n55566 & ~n55567;
  assign n9131 = n55579 | ~n55580;
  assign n55582 = P1_P1_LWORD_REG_11_ & ~n55518;
  assign n55583 = P1_P1_EAX_REG_11_ & n55520;
  assign n55584 = P1_BUF1_REG_11_ & n12460;
  assign n55585 = ~n47147 & ~n47151;
  assign n55586 = n47147 & n47151;
  assign n55587 = ~n55585 & ~n55586;
  assign n55588 = n47192 & ~n55587;
  assign n55589 = ~n47152 & ~n47153;
  assign n55590 = ~n47192 & ~n55589;
  assign n55591 = ~n55588 & ~n55590;
  assign n55592 = ~n12460 & ~n55591;
  assign n55593 = ~n55584 & ~n55592;
  assign n55594 = n55532 & ~n55593;
  assign n55595 = ~n55582 & ~n55583;
  assign n9136 = n55594 | ~n55595;
  assign n55597 = P1_P1_LWORD_REG_10_ & ~n55518;
  assign n55598 = P1_P1_EAX_REG_10_ & n55520;
  assign n55599 = P1_BUF1_REG_10_ & n12460;
  assign n55600 = n47162 & ~n47190;
  assign n55601 = ~n47162 & n47190;
  assign n55602 = ~n55600 & ~n55601;
  assign n55603 = ~n47161 & n55602;
  assign n55604 = n47161 & n55601;
  assign n55605 = ~n55603 & ~n55604;
  assign n55606 = n47163 & ~n47190;
  assign n55607 = n55605 & ~n55606;
  assign n55608 = ~n12460 & ~n55607;
  assign n55609 = ~n55599 & ~n55608;
  assign n55610 = n55532 & ~n55609;
  assign n55611 = ~n55597 & ~n55598;
  assign n9141 = n55610 | ~n55611;
  assign n55613 = P1_P1_LWORD_REG_9_ & ~n55518;
  assign n55614 = P1_P1_EAX_REG_9_ & n55520;
  assign n55615 = P1_BUF1_REG_9_ & n12460;
  assign n55616 = ~n47174 & ~n47175;
  assign n55617 = n47188 & n55616;
  assign n55618 = ~n47188 & ~n55616;
  assign n55619 = ~n55617 & ~n55618;
  assign n55620 = ~n12460 & ~n55619;
  assign n55621 = ~n55615 & ~n55620;
  assign n55622 = n55532 & ~n55621;
  assign n55623 = ~n55613 & ~n55614;
  assign n9146 = n55622 | ~n55623;
  assign n55625 = P1_P1_LWORD_REG_8_ & ~n55518;
  assign n55626 = P1_P1_EAX_REG_8_ & n55520;
  assign n55627 = P1_BUF1_REG_8_ & n12460;
  assign n55628 = ~n47176 & ~n47185;
  assign n55629 = n47176 & n47185;
  assign n55630 = ~n55628 & ~n55629;
  assign n55631 = n47178 & ~n55630;
  assign n55632 = ~n47176 & n47185;
  assign n55633 = ~n47178 & n55632;
  assign n55634 = n47179 & ~n47185;
  assign n55635 = ~n55631 & ~n55633;
  assign n55636 = ~n55634 & n55635;
  assign n55637 = ~n12460 & ~n55636;
  assign n55638 = ~n55627 & ~n55637;
  assign n55639 = n55532 & ~n55638;
  assign n55640 = ~n55625 & ~n55626;
  assign n9151 = n55639 | ~n55640;
  assign n55642 = P1_P1_LWORD_REG_7_ & ~n55518;
  assign n55643 = P1_P1_EAX_REG_7_ & n55520;
  assign n55644 = ~n44368 & n55532;
  assign n55645 = ~n55642 & ~n55643;
  assign n9156 = n55644 | ~n55645;
  assign n55647 = P1_P1_LWORD_REG_6_ & ~n55518;
  assign n55648 = P1_P1_EAX_REG_6_ & n55520;
  assign n55649 = ~n50203 & n55532;
  assign n55650 = ~n55647 & ~n55648;
  assign n9161 = n55649 | ~n55650;
  assign n55652 = P1_P1_LWORD_REG_5_ & ~n55518;
  assign n55653 = P1_P1_EAX_REG_5_ & n55520;
  assign n55654 = ~n50250 & n55532;
  assign n55655 = ~n55652 & ~n55653;
  assign n9166 = n55654 | ~n55655;
  assign n55657 = ~n50294 & n55532;
  assign n55658 = P1_P1_EAX_REG_4_ & n55520;
  assign n55659 = P1_P1_LWORD_REG_4_ & ~n55518;
  assign n55660 = ~n55657 & ~n55658;
  assign n9171 = n55659 | ~n55660;
  assign n55662 = ~n50338 & n55532;
  assign n55663 = P1_P1_EAX_REG_3_ & n55520;
  assign n55664 = P1_P1_LWORD_REG_3_ & ~n55518;
  assign n55665 = ~n55662 & ~n55663;
  assign n9176 = n55664 | ~n55665;
  assign n55667 = ~n50380 & n55532;
  assign n55668 = P1_P1_EAX_REG_2_ & n55520;
  assign n55669 = P1_P1_LWORD_REG_2_ & ~n55518;
  assign n55670 = ~n55667 & ~n55668;
  assign n9181 = n55669 | ~n55670;
  assign n55672 = ~n50425 & n55532;
  assign n55673 = P1_P1_EAX_REG_1_ & n55520;
  assign n55674 = P1_P1_LWORD_REG_1_ & ~n55518;
  assign n55675 = ~n55672 & ~n55673;
  assign n9186 = n55674 | ~n55675;
  assign n55677 = ~n50458 & n55532;
  assign n55678 = P1_P1_EAX_REG_0_ & n55520;
  assign n55679 = P1_P1_LWORD_REG_0_ & ~n55518;
  assign n55680 = ~n55677 & ~n55678;
  assign n9191 = n55679 | ~n55680;
  assign n55682 = P1_P1_UWORD_REG_14_ & ~n55518;
  assign n55683 = P1_P1_EAX_REG_30_ & n55520;
  assign n55684 = ~n55682 & ~n55683;
  assign n9196 = n55549 | ~n55684;
  assign n55686 = P1_P1_UWORD_REG_13_ & ~n55518;
  assign n55687 = P1_P1_EAX_REG_29_ & n55520;
  assign n55688 = ~n55686 & ~n55687;
  assign n9201 = n55563 | ~n55688;
  assign n55690 = P1_P1_UWORD_REG_12_ & ~n55518;
  assign n55691 = P1_P1_EAX_REG_28_ & n55520;
  assign n55692 = ~n55690 & ~n55691;
  assign n9206 = n55579 | ~n55692;
  assign n55694 = P1_P1_UWORD_REG_11_ & ~n55518;
  assign n55695 = P1_P1_EAX_REG_27_ & n55520;
  assign n55696 = ~n55694 & ~n55695;
  assign n9211 = n55594 | ~n55696;
  assign n55698 = P1_P1_UWORD_REG_10_ & ~n55518;
  assign n55699 = P1_P1_EAX_REG_26_ & n55520;
  assign n55700 = ~n55698 & ~n55699;
  assign n9216 = n55610 | ~n55700;
  assign n55702 = P1_P1_UWORD_REG_9_ & ~n55518;
  assign n55703 = P1_P1_EAX_REG_25_ & n55520;
  assign n55704 = ~n55702 & ~n55703;
  assign n9221 = n55622 | ~n55704;
  assign n55706 = P1_P1_UWORD_REG_8_ & ~n55518;
  assign n55707 = P1_P1_EAX_REG_24_ & n55520;
  assign n55708 = ~n55706 & ~n55707;
  assign n9226 = n55639 | ~n55708;
  assign n55710 = P1_P1_UWORD_REG_7_ & ~n55518;
  assign n55711 = P1_P1_EAX_REG_23_ & n55520;
  assign n55712 = ~n55710 & ~n55711;
  assign n9231 = n55644 | ~n55712;
  assign n55714 = P1_P1_UWORD_REG_6_ & ~n55518;
  assign n55715 = P1_P1_EAX_REG_22_ & n55520;
  assign n55716 = ~n55714 & ~n55715;
  assign n9236 = n55649 | ~n55716;
  assign n55718 = P1_P1_UWORD_REG_5_ & ~n55518;
  assign n55719 = P1_P1_EAX_REG_21_ & n55520;
  assign n55720 = ~n55718 & ~n55719;
  assign n9241 = n55654 | ~n55720;
  assign n55722 = P1_P1_EAX_REG_20_ & n55520;
  assign n55723 = P1_P1_UWORD_REG_4_ & ~n55518;
  assign n55724 = ~n55657 & ~n55722;
  assign n9246 = n55723 | ~n55724;
  assign n55726 = P1_P1_EAX_REG_19_ & n55520;
  assign n55727 = P1_P1_UWORD_REG_3_ & ~n55518;
  assign n55728 = ~n55662 & ~n55726;
  assign n9251 = n55727 | ~n55728;
  assign n55730 = P1_P1_EAX_REG_18_ & n55520;
  assign n55731 = P1_P1_UWORD_REG_2_ & ~n55518;
  assign n55732 = ~n55667 & ~n55730;
  assign n9256 = n55731 | ~n55732;
  assign n55734 = P1_P1_EAX_REG_17_ & n55520;
  assign n55735 = P1_P1_UWORD_REG_1_ & ~n55518;
  assign n55736 = ~n55672 & ~n55734;
  assign n9261 = n55735 | ~n55736;
  assign n55738 = P1_P1_EAX_REG_16_ & n55520;
  assign n55739 = P1_P1_UWORD_REG_0_ & ~n55518;
  assign n55740 = ~n55677 & ~n55738;
  assign n9266 = n55739 | ~n55740;
  assign n55742 = ~P1_P1_STATE2_REG_0_ & n43336;
  assign n55743 = n43342 & n43979;
  assign n55744 = ~n43864 & n55743;
  assign n55745 = ~n55742 & ~n55744;
  assign n55746 = P1_P1_STATE2_REG_0_ & ~n55745;
  assign n55747 = P1_P1_EAX_REG_0_ & n55746;
  assign n55748 = ~P1_P1_STATE2_REG_0_ & ~n55745;
  assign n55749 = P1_P1_LWORD_REG_0_ & n55748;
  assign n55750 = P1_P1_DATAO_REG_0_ & n55745;
  assign n55751 = ~n55747 & ~n55749;
  assign n9271 = n55750 | ~n55751;
  assign n55753 = P1_P1_EAX_REG_1_ & n55746;
  assign n55754 = P1_P1_LWORD_REG_1_ & n55748;
  assign n55755 = P1_P1_DATAO_REG_1_ & n55745;
  assign n55756 = ~n55753 & ~n55754;
  assign n9276 = n55755 | ~n55756;
  assign n55758 = P1_P1_EAX_REG_2_ & n55746;
  assign n55759 = P1_P1_LWORD_REG_2_ & n55748;
  assign n55760 = P1_P1_DATAO_REG_2_ & n55745;
  assign n55761 = ~n55758 & ~n55759;
  assign n9281 = n55760 | ~n55761;
  assign n55763 = P1_P1_EAX_REG_3_ & n55746;
  assign n55764 = P1_P1_LWORD_REG_3_ & n55748;
  assign n55765 = P1_P1_DATAO_REG_3_ & n55745;
  assign n55766 = ~n55763 & ~n55764;
  assign n9286 = n55765 | ~n55766;
  assign n55768 = P1_P1_EAX_REG_4_ & n55746;
  assign n55769 = P1_P1_LWORD_REG_4_ & n55748;
  assign n55770 = P1_P1_DATAO_REG_4_ & n55745;
  assign n55771 = ~n55768 & ~n55769;
  assign n9291 = n55770 | ~n55771;
  assign n55773 = P1_P1_EAX_REG_5_ & n55746;
  assign n55774 = P1_P1_LWORD_REG_5_ & n55748;
  assign n55775 = P1_P1_DATAO_REG_5_ & n55745;
  assign n55776 = ~n55773 & ~n55774;
  assign n9296 = n55775 | ~n55776;
  assign n55778 = P1_P1_EAX_REG_6_ & n55746;
  assign n55779 = P1_P1_LWORD_REG_6_ & n55748;
  assign n55780 = P1_P1_DATAO_REG_6_ & n55745;
  assign n55781 = ~n55778 & ~n55779;
  assign n9301 = n55780 | ~n55781;
  assign n55783 = P1_P1_EAX_REG_7_ & n55746;
  assign n55784 = P1_P1_LWORD_REG_7_ & n55748;
  assign n55785 = P1_P1_DATAO_REG_7_ & n55745;
  assign n55786 = ~n55783 & ~n55784;
  assign n9306 = n55785 | ~n55786;
  assign n55788 = P1_P1_EAX_REG_8_ & n55746;
  assign n55789 = P1_P1_LWORD_REG_8_ & n55748;
  assign n55790 = P1_P1_DATAO_REG_8_ & n55745;
  assign n55791 = ~n55788 & ~n55789;
  assign n9311 = n55790 | ~n55791;
  assign n55793 = P1_P1_EAX_REG_9_ & n55746;
  assign n55794 = P1_P1_LWORD_REG_9_ & n55748;
  assign n55795 = P1_P1_DATAO_REG_9_ & n55745;
  assign n55796 = ~n55793 & ~n55794;
  assign n9316 = n55795 | ~n55796;
  assign n55798 = P1_P1_EAX_REG_10_ & n55746;
  assign n55799 = P1_P1_LWORD_REG_10_ & n55748;
  assign n55800 = P1_P1_DATAO_REG_10_ & n55745;
  assign n55801 = ~n55798 & ~n55799;
  assign n9321 = n55800 | ~n55801;
  assign n55803 = P1_P1_EAX_REG_11_ & n55746;
  assign n55804 = P1_P1_LWORD_REG_11_ & n55748;
  assign n55805 = P1_P1_DATAO_REG_11_ & n55745;
  assign n55806 = ~n55803 & ~n55804;
  assign n9326 = n55805 | ~n55806;
  assign n55808 = P1_P1_EAX_REG_12_ & n55746;
  assign n55809 = P1_P1_LWORD_REG_12_ & n55748;
  assign n55810 = P1_P1_DATAO_REG_12_ & n55745;
  assign n55811 = ~n55808 & ~n55809;
  assign n9331 = n55810 | ~n55811;
  assign n55813 = P1_P1_EAX_REG_13_ & n55746;
  assign n55814 = P1_P1_LWORD_REG_13_ & n55748;
  assign n55815 = P1_P1_DATAO_REG_13_ & n55745;
  assign n55816 = ~n55813 & ~n55814;
  assign n9336 = n55815 | ~n55816;
  assign n55818 = P1_P1_EAX_REG_14_ & n55746;
  assign n55819 = P1_P1_LWORD_REG_14_ & n55748;
  assign n55820 = P1_P1_DATAO_REG_14_ & n55745;
  assign n55821 = ~n55818 & ~n55819;
  assign n9341 = n55820 | ~n55821;
  assign n55823 = P1_P1_EAX_REG_15_ & n55746;
  assign n55824 = P1_P1_LWORD_REG_15_ & n55748;
  assign n55825 = P1_P1_DATAO_REG_15_ & n55745;
  assign n55826 = ~n55823 & ~n55824;
  assign n9346 = n55825 | ~n55826;
  assign n55828 = P1_P1_UWORD_REG_0_ & n55748;
  assign n55829 = P1_P1_DATAO_REG_16_ & n55745;
  assign n55830 = ~n55828 & ~n55829;
  assign n55831 = ~n43623 & n55746;
  assign n55832 = P1_P1_EAX_REG_16_ & n55831;
  assign n9351 = ~n55830 | n55832;
  assign n55834 = P1_P1_UWORD_REG_1_ & n55748;
  assign n55835 = P1_P1_DATAO_REG_17_ & n55745;
  assign n55836 = ~n55834 & ~n55835;
  assign n55837 = P1_P1_EAX_REG_17_ & n55831;
  assign n9356 = ~n55836 | n55837;
  assign n55839 = P1_P1_UWORD_REG_2_ & n55748;
  assign n55840 = P1_P1_DATAO_REG_18_ & n55745;
  assign n55841 = ~n55839 & ~n55840;
  assign n55842 = P1_P1_EAX_REG_18_ & n55831;
  assign n9361 = ~n55841 | n55842;
  assign n55844 = P1_P1_UWORD_REG_3_ & n55748;
  assign n55845 = P1_P1_DATAO_REG_19_ & n55745;
  assign n55846 = ~n55844 & ~n55845;
  assign n55847 = P1_P1_EAX_REG_19_ & n55831;
  assign n9366 = ~n55846 | n55847;
  assign n55849 = P1_P1_UWORD_REG_4_ & n55748;
  assign n55850 = P1_P1_DATAO_REG_20_ & n55745;
  assign n55851 = ~n55849 & ~n55850;
  assign n55852 = P1_P1_EAX_REG_20_ & n55831;
  assign n9371 = ~n55851 | n55852;
  assign n55854 = P1_P1_UWORD_REG_5_ & n55748;
  assign n55855 = P1_P1_DATAO_REG_21_ & n55745;
  assign n55856 = ~n55854 & ~n55855;
  assign n55857 = P1_P1_EAX_REG_21_ & n55831;
  assign n9376 = ~n55856 | n55857;
  assign n55859 = P1_P1_UWORD_REG_6_ & n55748;
  assign n55860 = P1_P1_DATAO_REG_22_ & n55745;
  assign n55861 = ~n55859 & ~n55860;
  assign n55862 = P1_P1_EAX_REG_22_ & n55831;
  assign n9381 = ~n55861 | n55862;
  assign n55864 = P1_P1_UWORD_REG_7_ & n55748;
  assign n55865 = P1_P1_DATAO_REG_23_ & n55745;
  assign n55866 = ~n55864 & ~n55865;
  assign n55867 = P1_P1_EAX_REG_23_ & n55831;
  assign n9386 = ~n55866 | n55867;
  assign n55869 = P1_P1_UWORD_REG_8_ & n55748;
  assign n55870 = P1_P1_DATAO_REG_24_ & n55745;
  assign n55871 = ~n55869 & ~n55870;
  assign n55872 = P1_P1_EAX_REG_24_ & n55831;
  assign n9391 = ~n55871 | n55872;
  assign n55874 = P1_P1_UWORD_REG_9_ & n55748;
  assign n55875 = P1_P1_DATAO_REG_25_ & n55745;
  assign n55876 = ~n55874 & ~n55875;
  assign n55877 = P1_P1_EAX_REG_25_ & n55831;
  assign n9396 = ~n55876 | n55877;
  assign n55879 = P1_P1_UWORD_REG_10_ & n55748;
  assign n55880 = P1_P1_DATAO_REG_26_ & n55745;
  assign n55881 = ~n55879 & ~n55880;
  assign n55882 = P1_P1_EAX_REG_26_ & n55831;
  assign n9401 = ~n55881 | n55882;
  assign n55884 = P1_P1_UWORD_REG_11_ & n55748;
  assign n55885 = P1_P1_DATAO_REG_27_ & n55745;
  assign n55886 = ~n55884 & ~n55885;
  assign n55887 = P1_P1_EAX_REG_27_ & n55831;
  assign n9406 = ~n55886 | n55887;
  assign n55889 = P1_P1_UWORD_REG_12_ & n55748;
  assign n55890 = P1_P1_DATAO_REG_28_ & n55745;
  assign n55891 = ~n55889 & ~n55890;
  assign n55892 = P1_P1_EAX_REG_28_ & n55831;
  assign n9411 = ~n55891 | n55892;
  assign n55894 = P1_P1_UWORD_REG_13_ & n55748;
  assign n55895 = P1_P1_DATAO_REG_29_ & n55745;
  assign n55896 = ~n55894 & ~n55895;
  assign n55897 = P1_P1_EAX_REG_29_ & n55831;
  assign n9416 = ~n55896 | n55897;
  assign n55899 = P1_P1_UWORD_REG_14_ & n55748;
  assign n55900 = P1_P1_DATAO_REG_30_ & n55745;
  assign n55901 = ~n55899 & ~n55900;
  assign n55902 = P1_P1_EAX_REG_30_ & n55831;
  assign n9421 = ~n55901 | n55902;
  assign n9426 = P1_P1_DATAO_REG_31_ & n55745;
  assign n55905 = n43858 & ~n43925;
  assign n55906 = n43979 & ~n55905;
  assign n55907 = n43712 & n55906;
  assign n55908 = ~n51995 & n55907;
  assign n55909 = ~n43495 & n55906;
  assign n55910 = ~n43712 & n55909;
  assign n55911 = ~n50458 & n55910;
  assign n55912 = P1_P1_EAX_REG_0_ & ~n55906;
  assign n55913 = n43495 & n55906;
  assign n55914 = ~P1_P1_EAX_REG_0_ & n55913;
  assign n55915 = ~n55912 & ~n55914;
  assign n55916 = ~n55908 & ~n55911;
  assign n9431 = ~n55915 | ~n55916;
  assign n55918 = ~n52118 & n55907;
  assign n55919 = ~n50425 & n55910;
  assign n55920 = P1_P1_EAX_REG_1_ & ~n55906;
  assign n55921 = P1_P1_EAX_REG_0_ & ~P1_P1_EAX_REG_1_;
  assign n55922 = ~P1_P1_EAX_REG_0_ & P1_P1_EAX_REG_1_;
  assign n55923 = ~n55921 & ~n55922;
  assign n55924 = n55913 & ~n55923;
  assign n55925 = ~n55920 & ~n55924;
  assign n55926 = ~n55918 & ~n55919;
  assign n9436 = ~n55925 | ~n55926;
  assign n55928 = ~n52233 & n55907;
  assign n55929 = ~n50380 & n55910;
  assign n55930 = P1_P1_EAX_REG_2_ & ~n55906;
  assign n55931 = P1_P1_EAX_REG_0_ & P1_P1_EAX_REG_1_;
  assign n55932 = ~P1_P1_EAX_REG_2_ & n55931;
  assign n55933 = P1_P1_EAX_REG_2_ & ~n55931;
  assign n55934 = ~n55932 & ~n55933;
  assign n55935 = n55913 & ~n55934;
  assign n55936 = ~n55930 & ~n55935;
  assign n55937 = ~n55928 & ~n55929;
  assign n9441 = ~n55936 | ~n55937;
  assign n55939 = ~n52355 & n55907;
  assign n55940 = ~n50338 & n55910;
  assign n55941 = P1_P1_EAX_REG_3_ & ~n55906;
  assign n55942 = P1_P1_EAX_REG_2_ & n55931;
  assign n55943 = ~P1_P1_EAX_REG_3_ & n55942;
  assign n55944 = P1_P1_EAX_REG_3_ & ~n55942;
  assign n55945 = ~n55943 & ~n55944;
  assign n55946 = n55913 & ~n55945;
  assign n55947 = ~n55941 & ~n55946;
  assign n55948 = ~n55939 & ~n55940;
  assign n9446 = ~n55947 | ~n55948;
  assign n55950 = ~n52484 & n55907;
  assign n55951 = ~n50294 & n55910;
  assign n55952 = P1_P1_EAX_REG_4_ & ~n55906;
  assign n55953 = P1_P1_EAX_REG_3_ & n55942;
  assign n55954 = ~P1_P1_EAX_REG_4_ & n55953;
  assign n55955 = P1_P1_EAX_REG_4_ & ~n55953;
  assign n55956 = ~n55954 & ~n55955;
  assign n55957 = n55913 & ~n55956;
  assign n55958 = ~n55952 & ~n55957;
  assign n55959 = ~n55950 & ~n55951;
  assign n9451 = ~n55958 | ~n55959;
  assign n55961 = ~n52625 & n55907;
  assign n55962 = ~n50250 & n55910;
  assign n55963 = P1_P1_EAX_REG_5_ & ~n55906;
  assign n55964 = P1_P1_EAX_REG_4_ & n55953;
  assign n55965 = ~P1_P1_EAX_REG_5_ & n55964;
  assign n55966 = P1_P1_EAX_REG_5_ & ~n55964;
  assign n55967 = ~n55965 & ~n55966;
  assign n55968 = n55913 & ~n55967;
  assign n55969 = ~n55963 & ~n55968;
  assign n55970 = ~n55961 & ~n55962;
  assign n9456 = ~n55969 | ~n55970;
  assign n55972 = ~n50203 & n55910;
  assign n55973 = P1_P1_EAX_REG_6_ & ~n55906;
  assign n55974 = P1_P1_EAX_REG_5_ & n55964;
  assign n55975 = ~P1_P1_EAX_REG_6_ & n55974;
  assign n55976 = P1_P1_EAX_REG_6_ & ~n55974;
  assign n55977 = ~n55975 & ~n55976;
  assign n55978 = n55913 & ~n55977;
  assign n55979 = ~n52759 & n55907;
  assign n55980 = ~n55973 & ~n55978;
  assign n55981 = ~n55979 & n55980;
  assign n9461 = n55972 | ~n55981;
  assign n55983 = ~n44368 & n55910;
  assign n55984 = P1_P1_EAX_REG_7_ & ~n55906;
  assign n55985 = P1_P1_EAX_REG_6_ & n55974;
  assign n55986 = ~P1_P1_EAX_REG_7_ & n55985;
  assign n55987 = P1_P1_EAX_REG_7_ & ~n55985;
  assign n55988 = ~n55986 & ~n55987;
  assign n55989 = n55913 & ~n55988;
  assign n55990 = ~n52029 & n55907;
  assign n55991 = ~n55984 & ~n55989;
  assign n55992 = ~n55990 & n55991;
  assign n9466 = n55983 | ~n55992;
  assign n55994 = ~n55638 & n55910;
  assign n55995 = P1_P1_EAX_REG_8_ & ~n55906;
  assign n55996 = P1_P1_EAX_REG_7_ & n55985;
  assign n55997 = ~P1_P1_EAX_REG_8_ & n55996;
  assign n55998 = P1_P1_EAX_REG_8_ & ~n55996;
  assign n55999 = ~n55997 & ~n55998;
  assign n56000 = n55913 & ~n55999;
  assign n56001 = ~n43872 & ~n43879;
  assign n56002 = ~n43823 & ~n56001;
  assign n56003 = n43353 & n56002;
  assign n56004 = P1_P1_INSTQUEUE_REG_15__0_ & n56003;
  assign n56005 = n43357 & n56002;
  assign n56006 = P1_P1_INSTQUEUE_REG_14__0_ & n56005;
  assign n56007 = n43344 & n56002;
  assign n56008 = P1_P1_INSTQUEUE_REG_13__0_ & n56007;
  assign n56009 = n43348 & n56002;
  assign n56010 = P1_P1_INSTQUEUE_REG_12__0_ & n56009;
  assign n56011 = ~n56004 & ~n56006;
  assign n56012 = ~n56008 & n56011;
  assign n56013 = ~n56010 & n56012;
  assign n56014 = n43823 & ~n56001;
  assign n56015 = n43353 & n56014;
  assign n56016 = P1_P1_INSTQUEUE_REG_11__0_ & n56015;
  assign n56017 = n43357 & n56014;
  assign n56018 = P1_P1_INSTQUEUE_REG_10__0_ & n56017;
  assign n56019 = n43344 & n56014;
  assign n56020 = P1_P1_INSTQUEUE_REG_9__0_ & n56019;
  assign n56021 = n43348 & n56014;
  assign n56022 = P1_P1_INSTQUEUE_REG_8__0_ & n56021;
  assign n56023 = ~n56016 & ~n56018;
  assign n56024 = ~n56020 & n56023;
  assign n56025 = ~n56022 & n56024;
  assign n56026 = ~n43823 & n56001;
  assign n56027 = n43353 & n56026;
  assign n56028 = P1_P1_INSTQUEUE_REG_7__0_ & n56027;
  assign n56029 = n43357 & n56026;
  assign n56030 = P1_P1_INSTQUEUE_REG_6__0_ & n56029;
  assign n56031 = n43344 & n56026;
  assign n56032 = P1_P1_INSTQUEUE_REG_5__0_ & n56031;
  assign n56033 = n43348 & n56026;
  assign n56034 = P1_P1_INSTQUEUE_REG_4__0_ & n56033;
  assign n56035 = ~n56028 & ~n56030;
  assign n56036 = ~n56032 & n56035;
  assign n56037 = ~n56034 & n56036;
  assign n56038 = n43823 & n56001;
  assign n56039 = n43353 & n56038;
  assign n56040 = P1_P1_INSTQUEUE_REG_3__0_ & n56039;
  assign n56041 = n43357 & n56038;
  assign n56042 = P1_P1_INSTQUEUE_REG_2__0_ & n56041;
  assign n56043 = n43344 & n56038;
  assign n56044 = P1_P1_INSTQUEUE_REG_1__0_ & n56043;
  assign n56045 = n43348 & n56038;
  assign n56046 = P1_P1_INSTQUEUE_REG_0__0_ & n56045;
  assign n56047 = ~n56040 & ~n56042;
  assign n56048 = ~n56044 & n56047;
  assign n56049 = ~n56046 & n56048;
  assign n56050 = n56013 & n56025;
  assign n56051 = n56037 & n56050;
  assign n56052 = n56049 & n56051;
  assign n56053 = n55907 & ~n56052;
  assign n56054 = ~n55995 & ~n56000;
  assign n56055 = ~n56053 & n56054;
  assign n9471 = n55994 | ~n56055;
  assign n56057 = ~n55621 & n55910;
  assign n56058 = P1_P1_EAX_REG_9_ & ~n55906;
  assign n56059 = P1_P1_EAX_REG_8_ & n55996;
  assign n56060 = ~P1_P1_EAX_REG_9_ & n56059;
  assign n56061 = P1_P1_EAX_REG_9_ & ~n56059;
  assign n56062 = ~n56060 & ~n56061;
  assign n56063 = n55913 & ~n56062;
  assign n56064 = P1_P1_INSTQUEUE_REG_15__1_ & n56003;
  assign n56065 = P1_P1_INSTQUEUE_REG_14__1_ & n56005;
  assign n56066 = P1_P1_INSTQUEUE_REG_13__1_ & n56007;
  assign n56067 = P1_P1_INSTQUEUE_REG_12__1_ & n56009;
  assign n56068 = ~n56064 & ~n56065;
  assign n56069 = ~n56066 & n56068;
  assign n56070 = ~n56067 & n56069;
  assign n56071 = P1_P1_INSTQUEUE_REG_11__1_ & n56015;
  assign n56072 = P1_P1_INSTQUEUE_REG_10__1_ & n56017;
  assign n56073 = P1_P1_INSTQUEUE_REG_9__1_ & n56019;
  assign n56074 = P1_P1_INSTQUEUE_REG_8__1_ & n56021;
  assign n56075 = ~n56071 & ~n56072;
  assign n56076 = ~n56073 & n56075;
  assign n56077 = ~n56074 & n56076;
  assign n56078 = P1_P1_INSTQUEUE_REG_7__1_ & n56027;
  assign n56079 = P1_P1_INSTQUEUE_REG_6__1_ & n56029;
  assign n56080 = P1_P1_INSTQUEUE_REG_5__1_ & n56031;
  assign n56081 = P1_P1_INSTQUEUE_REG_4__1_ & n56033;
  assign n56082 = ~n56078 & ~n56079;
  assign n56083 = ~n56080 & n56082;
  assign n56084 = ~n56081 & n56083;
  assign n56085 = P1_P1_INSTQUEUE_REG_3__1_ & n56039;
  assign n56086 = P1_P1_INSTQUEUE_REG_2__1_ & n56041;
  assign n56087 = P1_P1_INSTQUEUE_REG_1__1_ & n56043;
  assign n56088 = P1_P1_INSTQUEUE_REG_0__1_ & n56045;
  assign n56089 = ~n56085 & ~n56086;
  assign n56090 = ~n56087 & n56089;
  assign n56091 = ~n56088 & n56090;
  assign n56092 = n56070 & n56077;
  assign n56093 = n56084 & n56092;
  assign n56094 = n56091 & n56093;
  assign n56095 = n55907 & ~n56094;
  assign n56096 = ~n56058 & ~n56063;
  assign n56097 = ~n56095 & n56096;
  assign n9476 = n56057 | ~n56097;
  assign n56099 = ~n55609 & n55910;
  assign n56100 = P1_P1_EAX_REG_10_ & ~n55906;
  assign n56101 = P1_P1_EAX_REG_9_ & n56059;
  assign n56102 = ~P1_P1_EAX_REG_10_ & n56101;
  assign n56103 = P1_P1_EAX_REG_10_ & ~n56101;
  assign n56104 = ~n56102 & ~n56103;
  assign n56105 = n55913 & ~n56104;
  assign n56106 = P1_P1_INSTQUEUE_REG_15__2_ & n56003;
  assign n56107 = P1_P1_INSTQUEUE_REG_14__2_ & n56005;
  assign n56108 = P1_P1_INSTQUEUE_REG_13__2_ & n56007;
  assign n56109 = P1_P1_INSTQUEUE_REG_12__2_ & n56009;
  assign n56110 = ~n56106 & ~n56107;
  assign n56111 = ~n56108 & n56110;
  assign n56112 = ~n56109 & n56111;
  assign n56113 = P1_P1_INSTQUEUE_REG_11__2_ & n56015;
  assign n56114 = P1_P1_INSTQUEUE_REG_10__2_ & n56017;
  assign n56115 = P1_P1_INSTQUEUE_REG_9__2_ & n56019;
  assign n56116 = P1_P1_INSTQUEUE_REG_8__2_ & n56021;
  assign n56117 = ~n56113 & ~n56114;
  assign n56118 = ~n56115 & n56117;
  assign n56119 = ~n56116 & n56118;
  assign n56120 = P1_P1_INSTQUEUE_REG_7__2_ & n56027;
  assign n56121 = P1_P1_INSTQUEUE_REG_6__2_ & n56029;
  assign n56122 = P1_P1_INSTQUEUE_REG_5__2_ & n56031;
  assign n56123 = P1_P1_INSTQUEUE_REG_4__2_ & n56033;
  assign n56124 = ~n56120 & ~n56121;
  assign n56125 = ~n56122 & n56124;
  assign n56126 = ~n56123 & n56125;
  assign n56127 = P1_P1_INSTQUEUE_REG_3__2_ & n56039;
  assign n56128 = P1_P1_INSTQUEUE_REG_2__2_ & n56041;
  assign n56129 = P1_P1_INSTQUEUE_REG_1__2_ & n56043;
  assign n56130 = P1_P1_INSTQUEUE_REG_0__2_ & n56045;
  assign n56131 = ~n56127 & ~n56128;
  assign n56132 = ~n56129 & n56131;
  assign n56133 = ~n56130 & n56132;
  assign n56134 = n56112 & n56119;
  assign n56135 = n56126 & n56134;
  assign n56136 = n56133 & n56135;
  assign n56137 = n55907 & ~n56136;
  assign n56138 = ~n56100 & ~n56105;
  assign n56139 = ~n56137 & n56138;
  assign n9481 = n56099 | ~n56139;
  assign n56141 = ~n55593 & n55910;
  assign n56142 = P1_P1_EAX_REG_11_ & ~n55906;
  assign n56143 = P1_P1_EAX_REG_10_ & n56101;
  assign n56144 = ~P1_P1_EAX_REG_11_ & n56143;
  assign n56145 = P1_P1_EAX_REG_11_ & ~n56143;
  assign n56146 = ~n56144 & ~n56145;
  assign n56147 = n55913 & ~n56146;
  assign n56148 = P1_P1_INSTQUEUE_REG_15__3_ & n56003;
  assign n56149 = P1_P1_INSTQUEUE_REG_14__3_ & n56005;
  assign n56150 = P1_P1_INSTQUEUE_REG_13__3_ & n56007;
  assign n56151 = P1_P1_INSTQUEUE_REG_12__3_ & n56009;
  assign n56152 = ~n56148 & ~n56149;
  assign n56153 = ~n56150 & n56152;
  assign n56154 = ~n56151 & n56153;
  assign n56155 = P1_P1_INSTQUEUE_REG_11__3_ & n56015;
  assign n56156 = P1_P1_INSTQUEUE_REG_10__3_ & n56017;
  assign n56157 = P1_P1_INSTQUEUE_REG_9__3_ & n56019;
  assign n56158 = P1_P1_INSTQUEUE_REG_8__3_ & n56021;
  assign n56159 = ~n56155 & ~n56156;
  assign n56160 = ~n56157 & n56159;
  assign n56161 = ~n56158 & n56160;
  assign n56162 = P1_P1_INSTQUEUE_REG_7__3_ & n56027;
  assign n56163 = P1_P1_INSTQUEUE_REG_6__3_ & n56029;
  assign n56164 = P1_P1_INSTQUEUE_REG_5__3_ & n56031;
  assign n56165 = P1_P1_INSTQUEUE_REG_4__3_ & n56033;
  assign n56166 = ~n56162 & ~n56163;
  assign n56167 = ~n56164 & n56166;
  assign n56168 = ~n56165 & n56167;
  assign n56169 = P1_P1_INSTQUEUE_REG_3__3_ & n56039;
  assign n56170 = P1_P1_INSTQUEUE_REG_2__3_ & n56041;
  assign n56171 = P1_P1_INSTQUEUE_REG_1__3_ & n56043;
  assign n56172 = P1_P1_INSTQUEUE_REG_0__3_ & n56045;
  assign n56173 = ~n56169 & ~n56170;
  assign n56174 = ~n56171 & n56173;
  assign n56175 = ~n56172 & n56174;
  assign n56176 = n56154 & n56161;
  assign n56177 = n56168 & n56176;
  assign n56178 = n56175 & n56177;
  assign n56179 = n55907 & ~n56178;
  assign n56180 = ~n56142 & ~n56147;
  assign n56181 = ~n56179 & n56180;
  assign n9486 = n56141 | ~n56181;
  assign n56183 = ~n55578 & n55910;
  assign n56184 = P1_P1_EAX_REG_12_ & ~n55906;
  assign n56185 = P1_P1_EAX_REG_11_ & n56143;
  assign n56186 = ~P1_P1_EAX_REG_12_ & n56185;
  assign n56187 = P1_P1_EAX_REG_12_ & ~n56185;
  assign n56188 = ~n56186 & ~n56187;
  assign n56189 = n55913 & ~n56188;
  assign n56190 = P1_P1_INSTQUEUE_REG_15__4_ & n56003;
  assign n56191 = P1_P1_INSTQUEUE_REG_14__4_ & n56005;
  assign n56192 = P1_P1_INSTQUEUE_REG_13__4_ & n56007;
  assign n56193 = P1_P1_INSTQUEUE_REG_12__4_ & n56009;
  assign n56194 = ~n56190 & ~n56191;
  assign n56195 = ~n56192 & n56194;
  assign n56196 = ~n56193 & n56195;
  assign n56197 = P1_P1_INSTQUEUE_REG_11__4_ & n56015;
  assign n56198 = P1_P1_INSTQUEUE_REG_10__4_ & n56017;
  assign n56199 = P1_P1_INSTQUEUE_REG_9__4_ & n56019;
  assign n56200 = P1_P1_INSTQUEUE_REG_8__4_ & n56021;
  assign n56201 = ~n56197 & ~n56198;
  assign n56202 = ~n56199 & n56201;
  assign n56203 = ~n56200 & n56202;
  assign n56204 = P1_P1_INSTQUEUE_REG_7__4_ & n56027;
  assign n56205 = P1_P1_INSTQUEUE_REG_6__4_ & n56029;
  assign n56206 = P1_P1_INSTQUEUE_REG_5__4_ & n56031;
  assign n56207 = P1_P1_INSTQUEUE_REG_4__4_ & n56033;
  assign n56208 = ~n56204 & ~n56205;
  assign n56209 = ~n56206 & n56208;
  assign n56210 = ~n56207 & n56209;
  assign n56211 = P1_P1_INSTQUEUE_REG_3__4_ & n56039;
  assign n56212 = P1_P1_INSTQUEUE_REG_2__4_ & n56041;
  assign n56213 = P1_P1_INSTQUEUE_REG_1__4_ & n56043;
  assign n56214 = P1_P1_INSTQUEUE_REG_0__4_ & n56045;
  assign n56215 = ~n56211 & ~n56212;
  assign n56216 = ~n56213 & n56215;
  assign n56217 = ~n56214 & n56216;
  assign n56218 = n56196 & n56203;
  assign n56219 = n56210 & n56218;
  assign n56220 = n56217 & n56219;
  assign n56221 = n55907 & ~n56220;
  assign n56222 = ~n56184 & ~n56189;
  assign n56223 = ~n56221 & n56222;
  assign n9491 = n56183 | ~n56223;
  assign n56225 = ~n55562 & n55910;
  assign n56226 = P1_P1_EAX_REG_13_ & ~n55906;
  assign n56227 = P1_P1_EAX_REG_12_ & n56185;
  assign n56228 = ~P1_P1_EAX_REG_13_ & n56227;
  assign n56229 = P1_P1_EAX_REG_13_ & ~n56227;
  assign n56230 = ~n56228 & ~n56229;
  assign n56231 = n55913 & ~n56230;
  assign n56232 = P1_P1_INSTQUEUE_REG_15__5_ & n56003;
  assign n56233 = P1_P1_INSTQUEUE_REG_14__5_ & n56005;
  assign n56234 = P1_P1_INSTQUEUE_REG_13__5_ & n56007;
  assign n56235 = P1_P1_INSTQUEUE_REG_12__5_ & n56009;
  assign n56236 = ~n56232 & ~n56233;
  assign n56237 = ~n56234 & n56236;
  assign n56238 = ~n56235 & n56237;
  assign n56239 = P1_P1_INSTQUEUE_REG_11__5_ & n56015;
  assign n56240 = P1_P1_INSTQUEUE_REG_10__5_ & n56017;
  assign n56241 = P1_P1_INSTQUEUE_REG_9__5_ & n56019;
  assign n56242 = P1_P1_INSTQUEUE_REG_8__5_ & n56021;
  assign n56243 = ~n56239 & ~n56240;
  assign n56244 = ~n56241 & n56243;
  assign n56245 = ~n56242 & n56244;
  assign n56246 = P1_P1_INSTQUEUE_REG_7__5_ & n56027;
  assign n56247 = P1_P1_INSTQUEUE_REG_6__5_ & n56029;
  assign n56248 = P1_P1_INSTQUEUE_REG_5__5_ & n56031;
  assign n56249 = P1_P1_INSTQUEUE_REG_4__5_ & n56033;
  assign n56250 = ~n56246 & ~n56247;
  assign n56251 = ~n56248 & n56250;
  assign n56252 = ~n56249 & n56251;
  assign n56253 = P1_P1_INSTQUEUE_REG_3__5_ & n56039;
  assign n56254 = P1_P1_INSTQUEUE_REG_2__5_ & n56041;
  assign n56255 = P1_P1_INSTQUEUE_REG_1__5_ & n56043;
  assign n56256 = P1_P1_INSTQUEUE_REG_0__5_ & n56045;
  assign n56257 = ~n56253 & ~n56254;
  assign n56258 = ~n56255 & n56257;
  assign n56259 = ~n56256 & n56258;
  assign n56260 = n56238 & n56245;
  assign n56261 = n56252 & n56260;
  assign n56262 = n56259 & n56261;
  assign n56263 = n55907 & ~n56262;
  assign n56264 = ~n56226 & ~n56231;
  assign n56265 = ~n56263 & n56264;
  assign n9496 = n56225 | ~n56265;
  assign n56267 = ~n55548 & n55910;
  assign n56268 = P1_P1_EAX_REG_14_ & ~n55906;
  assign n56269 = P1_P1_EAX_REG_13_ & n56227;
  assign n56270 = ~P1_P1_EAX_REG_14_ & n56269;
  assign n56271 = P1_P1_EAX_REG_14_ & ~n56269;
  assign n56272 = ~n56270 & ~n56271;
  assign n56273 = n55913 & ~n56272;
  assign n56274 = P1_P1_INSTQUEUE_REG_15__6_ & n56003;
  assign n56275 = P1_P1_INSTQUEUE_REG_14__6_ & n56005;
  assign n56276 = P1_P1_INSTQUEUE_REG_13__6_ & n56007;
  assign n56277 = P1_P1_INSTQUEUE_REG_12__6_ & n56009;
  assign n56278 = ~n56274 & ~n56275;
  assign n56279 = ~n56276 & n56278;
  assign n56280 = ~n56277 & n56279;
  assign n56281 = P1_P1_INSTQUEUE_REG_11__6_ & n56015;
  assign n56282 = P1_P1_INSTQUEUE_REG_10__6_ & n56017;
  assign n56283 = P1_P1_INSTQUEUE_REG_9__6_ & n56019;
  assign n56284 = P1_P1_INSTQUEUE_REG_8__6_ & n56021;
  assign n56285 = ~n56281 & ~n56282;
  assign n56286 = ~n56283 & n56285;
  assign n56287 = ~n56284 & n56286;
  assign n56288 = P1_P1_INSTQUEUE_REG_7__6_ & n56027;
  assign n56289 = P1_P1_INSTQUEUE_REG_6__6_ & n56029;
  assign n56290 = P1_P1_INSTQUEUE_REG_5__6_ & n56031;
  assign n56291 = P1_P1_INSTQUEUE_REG_4__6_ & n56033;
  assign n56292 = ~n56288 & ~n56289;
  assign n56293 = ~n56290 & n56292;
  assign n56294 = ~n56291 & n56293;
  assign n56295 = P1_P1_INSTQUEUE_REG_3__6_ & n56039;
  assign n56296 = P1_P1_INSTQUEUE_REG_2__6_ & n56041;
  assign n56297 = P1_P1_INSTQUEUE_REG_1__6_ & n56043;
  assign n56298 = P1_P1_INSTQUEUE_REG_0__6_ & n56045;
  assign n56299 = ~n56295 & ~n56296;
  assign n56300 = ~n56297 & n56299;
  assign n56301 = ~n56298 & n56300;
  assign n56302 = n56280 & n56287;
  assign n56303 = n56294 & n56302;
  assign n56304 = n56301 & n56303;
  assign n56305 = n55907 & ~n56304;
  assign n56306 = ~n56268 & ~n56273;
  assign n56307 = ~n56305 & n56306;
  assign n9501 = n56267 | ~n56307;
  assign n56309 = ~n55531 & n55910;
  assign n56310 = P1_P1_EAX_REG_15_ & ~n55906;
  assign n56311 = P1_P1_EAX_REG_14_ & n56269;
  assign n56312 = ~P1_P1_EAX_REG_15_ & n56311;
  assign n56313 = P1_P1_EAX_REG_15_ & ~n56311;
  assign n56314 = ~n56312 & ~n56313;
  assign n56315 = n55913 & ~n56314;
  assign n56316 = P1_P1_INSTQUEUE_REG_15__7_ & n56003;
  assign n56317 = P1_P1_INSTQUEUE_REG_14__7_ & n56005;
  assign n56318 = P1_P1_INSTQUEUE_REG_13__7_ & n56007;
  assign n56319 = P1_P1_INSTQUEUE_REG_12__7_ & n56009;
  assign n56320 = ~n56316 & ~n56317;
  assign n56321 = ~n56318 & n56320;
  assign n56322 = ~n56319 & n56321;
  assign n56323 = P1_P1_INSTQUEUE_REG_11__7_ & n56015;
  assign n56324 = P1_P1_INSTQUEUE_REG_10__7_ & n56017;
  assign n56325 = P1_P1_INSTQUEUE_REG_9__7_ & n56019;
  assign n56326 = P1_P1_INSTQUEUE_REG_8__7_ & n56021;
  assign n56327 = ~n56323 & ~n56324;
  assign n56328 = ~n56325 & n56327;
  assign n56329 = ~n56326 & n56328;
  assign n56330 = P1_P1_INSTQUEUE_REG_7__7_ & n56027;
  assign n56331 = P1_P1_INSTQUEUE_REG_6__7_ & n56029;
  assign n56332 = P1_P1_INSTQUEUE_REG_5__7_ & n56031;
  assign n56333 = P1_P1_INSTQUEUE_REG_4__7_ & n56033;
  assign n56334 = ~n56330 & ~n56331;
  assign n56335 = ~n56332 & n56334;
  assign n56336 = ~n56333 & n56335;
  assign n56337 = P1_P1_INSTQUEUE_REG_3__7_ & n56039;
  assign n56338 = P1_P1_INSTQUEUE_REG_2__7_ & n56041;
  assign n56339 = P1_P1_INSTQUEUE_REG_1__7_ & n56043;
  assign n56340 = P1_P1_INSTQUEUE_REG_0__7_ & n56045;
  assign n56341 = ~n56337 & ~n56338;
  assign n56342 = ~n56339 & n56341;
  assign n56343 = ~n56340 & n56342;
  assign n56344 = n56322 & n56329;
  assign n56345 = n56336 & n56344;
  assign n56346 = n56343 & n56345;
  assign n56347 = n55907 & ~n56346;
  assign n56348 = ~n56310 & ~n56315;
  assign n56349 = ~n56347 & n56348;
  assign n9506 = n56309 | ~n56349;
  assign n56351 = P1_P1_INSTQUEUERD_ADDR_REG_2_ & ~n43357;
  assign n56352 = ~P1_P1_INSTQUEUERD_ADDR_REG_3_ & n56351;
  assign n56353 = P1_P1_INSTQUEUERD_ADDR_REG_3_ & ~n56351;
  assign n56354 = ~n56352 & ~n56353;
  assign n56355 = ~n43358 & ~n56351;
  assign n56356 = n56354 & n56355;
  assign n56357 = n51945 & n56356;
  assign n56358 = P1_P1_INSTQUEUE_REG_7__0_ & n56357;
  assign n56359 = n51942 & n56356;
  assign n56360 = P1_P1_INSTQUEUE_REG_6__0_ & n56359;
  assign n56361 = n51951 & n56356;
  assign n56362 = P1_P1_INSTQUEUE_REG_5__0_ & n56361;
  assign n56363 = n51948 & n56356;
  assign n56364 = P1_P1_INSTQUEUE_REG_4__0_ & n56363;
  assign n56365 = ~n56358 & ~n56360;
  assign n56366 = ~n56362 & n56365;
  assign n56367 = ~n56364 & n56366;
  assign n56368 = n56354 & ~n56355;
  assign n56369 = n51945 & n56368;
  assign n56370 = P1_P1_INSTQUEUE_REG_3__0_ & n56369;
  assign n56371 = n51942 & n56368;
  assign n56372 = P1_P1_INSTQUEUE_REG_2__0_ & n56371;
  assign n56373 = n51951 & n56368;
  assign n56374 = P1_P1_INSTQUEUE_REG_1__0_ & n56373;
  assign n56375 = n51948 & n56368;
  assign n56376 = P1_P1_INSTQUEUE_REG_0__0_ & n56375;
  assign n56377 = ~n56370 & ~n56372;
  assign n56378 = ~n56374 & n56377;
  assign n56379 = ~n56376 & n56378;
  assign n56380 = ~n56354 & n56355;
  assign n56381 = n51945 & n56380;
  assign n56382 = P1_P1_INSTQUEUE_REG_15__0_ & n56381;
  assign n56383 = n51942 & n56380;
  assign n56384 = P1_P1_INSTQUEUE_REG_14__0_ & n56383;
  assign n56385 = n51951 & n56380;
  assign n56386 = P1_P1_INSTQUEUE_REG_13__0_ & n56385;
  assign n56387 = n51948 & n56380;
  assign n56388 = P1_P1_INSTQUEUE_REG_12__0_ & n56387;
  assign n56389 = ~n56382 & ~n56384;
  assign n56390 = ~n56386 & n56389;
  assign n56391 = ~n56388 & n56390;
  assign n56392 = ~n56354 & ~n56355;
  assign n56393 = n51945 & n56392;
  assign n56394 = P1_P1_INSTQUEUE_REG_11__0_ & n56393;
  assign n56395 = n51942 & n56392;
  assign n56396 = P1_P1_INSTQUEUE_REG_10__0_ & n56395;
  assign n56397 = n51951 & n56392;
  assign n56398 = P1_P1_INSTQUEUE_REG_9__0_ & n56397;
  assign n56399 = n51948 & n56392;
  assign n56400 = P1_P1_INSTQUEUE_REG_8__0_ & n56399;
  assign n56401 = ~n56394 & ~n56396;
  assign n56402 = ~n56398 & n56401;
  assign n56403 = ~n56400 & n56402;
  assign n56404 = n56367 & n56379;
  assign n56405 = n56391 & n56404;
  assign n56406 = n56403 & n56405;
  assign n56407 = n55907 & ~n56406;
  assign n56408 = n43401 & n55909;
  assign n56409 = ~n50458 & n56408;
  assign n56410 = P1_P1_EAX_REG_16_ & ~n55906;
  assign n56411 = P1_P1_EAX_REG_15_ & n56311;
  assign n56412 = ~P1_P1_EAX_REG_16_ & n56411;
  assign n56413 = P1_P1_EAX_REG_16_ & ~n56411;
  assign n56414 = ~n56412 & ~n56413;
  assign n56415 = n55913 & ~n56414;
  assign n56416 = ~n56410 & ~n56415;
  assign n56417 = ~n43432 & n55909;
  assign n56418 = ~n50473 & n56417;
  assign n56419 = ~n56407 & ~n56409;
  assign n56420 = n56416 & n56419;
  assign n9511 = n56418 | ~n56420;
  assign n56422 = P1_P1_INSTQUEUE_REG_7__1_ & n56357;
  assign n56423 = P1_P1_INSTQUEUE_REG_6__1_ & n56359;
  assign n56424 = P1_P1_INSTQUEUE_REG_5__1_ & n56361;
  assign n56425 = P1_P1_INSTQUEUE_REG_4__1_ & n56363;
  assign n56426 = ~n56422 & ~n56423;
  assign n56427 = ~n56424 & n56426;
  assign n56428 = ~n56425 & n56427;
  assign n56429 = P1_P1_INSTQUEUE_REG_3__1_ & n56369;
  assign n56430 = P1_P1_INSTQUEUE_REG_2__1_ & n56371;
  assign n56431 = P1_P1_INSTQUEUE_REG_1__1_ & n56373;
  assign n56432 = P1_P1_INSTQUEUE_REG_0__1_ & n56375;
  assign n56433 = ~n56429 & ~n56430;
  assign n56434 = ~n56431 & n56433;
  assign n56435 = ~n56432 & n56434;
  assign n56436 = P1_P1_INSTQUEUE_REG_15__1_ & n56381;
  assign n56437 = P1_P1_INSTQUEUE_REG_14__1_ & n56383;
  assign n56438 = P1_P1_INSTQUEUE_REG_13__1_ & n56385;
  assign n56439 = P1_P1_INSTQUEUE_REG_12__1_ & n56387;
  assign n56440 = ~n56436 & ~n56437;
  assign n56441 = ~n56438 & n56440;
  assign n56442 = ~n56439 & n56441;
  assign n56443 = P1_P1_INSTQUEUE_REG_11__1_ & n56393;
  assign n56444 = P1_P1_INSTQUEUE_REG_10__1_ & n56395;
  assign n56445 = P1_P1_INSTQUEUE_REG_9__1_ & n56397;
  assign n56446 = P1_P1_INSTQUEUE_REG_8__1_ & n56399;
  assign n56447 = ~n56443 & ~n56444;
  assign n56448 = ~n56445 & n56447;
  assign n56449 = ~n56446 & n56448;
  assign n56450 = n56428 & n56435;
  assign n56451 = n56442 & n56450;
  assign n56452 = n56449 & n56451;
  assign n56453 = n55907 & ~n56452;
  assign n56454 = ~n50425 & n56408;
  assign n56455 = P1_P1_EAX_REG_17_ & ~n55906;
  assign n56456 = P1_P1_EAX_REG_16_ & n56411;
  assign n56457 = ~P1_P1_EAX_REG_17_ & n56456;
  assign n56458 = P1_P1_EAX_REG_17_ & ~n56456;
  assign n56459 = ~n56457 & ~n56458;
  assign n56460 = n55913 & ~n56459;
  assign n56461 = ~n56455 & ~n56460;
  assign n56462 = ~n50436 & n56417;
  assign n56463 = ~n56453 & ~n56454;
  assign n56464 = n56461 & n56463;
  assign n9516 = n56462 | ~n56464;
  assign n56466 = P1_P1_INSTQUEUE_REG_7__2_ & n56357;
  assign n56467 = P1_P1_INSTQUEUE_REG_6__2_ & n56359;
  assign n56468 = P1_P1_INSTQUEUE_REG_5__2_ & n56361;
  assign n56469 = P1_P1_INSTQUEUE_REG_4__2_ & n56363;
  assign n56470 = ~n56466 & ~n56467;
  assign n56471 = ~n56468 & n56470;
  assign n56472 = ~n56469 & n56471;
  assign n56473 = P1_P1_INSTQUEUE_REG_3__2_ & n56369;
  assign n56474 = P1_P1_INSTQUEUE_REG_2__2_ & n56371;
  assign n56475 = P1_P1_INSTQUEUE_REG_1__2_ & n56373;
  assign n56476 = P1_P1_INSTQUEUE_REG_0__2_ & n56375;
  assign n56477 = ~n56473 & ~n56474;
  assign n56478 = ~n56475 & n56477;
  assign n56479 = ~n56476 & n56478;
  assign n56480 = P1_P1_INSTQUEUE_REG_15__2_ & n56381;
  assign n56481 = P1_P1_INSTQUEUE_REG_14__2_ & n56383;
  assign n56482 = P1_P1_INSTQUEUE_REG_13__2_ & n56385;
  assign n56483 = P1_P1_INSTQUEUE_REG_12__2_ & n56387;
  assign n56484 = ~n56480 & ~n56481;
  assign n56485 = ~n56482 & n56484;
  assign n56486 = ~n56483 & n56485;
  assign n56487 = P1_P1_INSTQUEUE_REG_11__2_ & n56393;
  assign n56488 = P1_P1_INSTQUEUE_REG_10__2_ & n56395;
  assign n56489 = P1_P1_INSTQUEUE_REG_9__2_ & n56397;
  assign n56490 = P1_P1_INSTQUEUE_REG_8__2_ & n56399;
  assign n56491 = ~n56487 & ~n56488;
  assign n56492 = ~n56489 & n56491;
  assign n56493 = ~n56490 & n56492;
  assign n56494 = n56472 & n56479;
  assign n56495 = n56486 & n56494;
  assign n56496 = n56493 & n56495;
  assign n56497 = n55907 & ~n56496;
  assign n56498 = ~n50380 & n56408;
  assign n56499 = P1_P1_EAX_REG_18_ & ~n55906;
  assign n56500 = P1_P1_EAX_REG_17_ & n56456;
  assign n56501 = ~P1_P1_EAX_REG_18_ & n56500;
  assign n56502 = P1_P1_EAX_REG_18_ & ~n56500;
  assign n56503 = ~n56501 & ~n56502;
  assign n56504 = n55913 & ~n56503;
  assign n56505 = ~n56499 & ~n56504;
  assign n56506 = ~n50396 & n56417;
  assign n56507 = ~n56497 & ~n56498;
  assign n56508 = n56505 & n56507;
  assign n9521 = n56506 | ~n56508;
  assign n56510 = P1_P1_INSTQUEUE_REG_7__3_ & n56357;
  assign n56511 = P1_P1_INSTQUEUE_REG_6__3_ & n56359;
  assign n56512 = P1_P1_INSTQUEUE_REG_5__3_ & n56361;
  assign n56513 = P1_P1_INSTQUEUE_REG_4__3_ & n56363;
  assign n56514 = ~n56510 & ~n56511;
  assign n56515 = ~n56512 & n56514;
  assign n56516 = ~n56513 & n56515;
  assign n56517 = P1_P1_INSTQUEUE_REG_3__3_ & n56369;
  assign n56518 = P1_P1_INSTQUEUE_REG_2__3_ & n56371;
  assign n56519 = P1_P1_INSTQUEUE_REG_1__3_ & n56373;
  assign n56520 = P1_P1_INSTQUEUE_REG_0__3_ & n56375;
  assign n56521 = ~n56517 & ~n56518;
  assign n56522 = ~n56519 & n56521;
  assign n56523 = ~n56520 & n56522;
  assign n56524 = P1_P1_INSTQUEUE_REG_15__3_ & n56381;
  assign n56525 = P1_P1_INSTQUEUE_REG_14__3_ & n56383;
  assign n56526 = P1_P1_INSTQUEUE_REG_13__3_ & n56385;
  assign n56527 = P1_P1_INSTQUEUE_REG_12__3_ & n56387;
  assign n56528 = ~n56524 & ~n56525;
  assign n56529 = ~n56526 & n56528;
  assign n56530 = ~n56527 & n56529;
  assign n56531 = P1_P1_INSTQUEUE_REG_11__3_ & n56393;
  assign n56532 = P1_P1_INSTQUEUE_REG_10__3_ & n56395;
  assign n56533 = P1_P1_INSTQUEUE_REG_9__3_ & n56397;
  assign n56534 = P1_P1_INSTQUEUE_REG_8__3_ & n56399;
  assign n56535 = ~n56531 & ~n56532;
  assign n56536 = ~n56533 & n56535;
  assign n56537 = ~n56534 & n56536;
  assign n56538 = n56516 & n56523;
  assign n56539 = n56530 & n56538;
  assign n56540 = n56537 & n56539;
  assign n56541 = n55907 & ~n56540;
  assign n56542 = ~n50338 & n56408;
  assign n56543 = P1_P1_EAX_REG_19_ & ~n55906;
  assign n56544 = P1_P1_EAX_REG_18_ & n56500;
  assign n56545 = ~P1_P1_EAX_REG_19_ & n56544;
  assign n56546 = P1_P1_EAX_REG_19_ & ~n56544;
  assign n56547 = ~n56545 & ~n56546;
  assign n56548 = n55913 & ~n56547;
  assign n56549 = ~n56543 & ~n56548;
  assign n56550 = ~n50352 & n56417;
  assign n56551 = ~n56541 & ~n56542;
  assign n56552 = n56549 & n56551;
  assign n9526 = n56550 | ~n56552;
  assign n56554 = P1_P1_INSTQUEUE_REG_7__4_ & n56357;
  assign n56555 = P1_P1_INSTQUEUE_REG_6__4_ & n56359;
  assign n56556 = P1_P1_INSTQUEUE_REG_5__4_ & n56361;
  assign n56557 = P1_P1_INSTQUEUE_REG_4__4_ & n56363;
  assign n56558 = ~n56554 & ~n56555;
  assign n56559 = ~n56556 & n56558;
  assign n56560 = ~n56557 & n56559;
  assign n56561 = P1_P1_INSTQUEUE_REG_3__4_ & n56369;
  assign n56562 = P1_P1_INSTQUEUE_REG_2__4_ & n56371;
  assign n56563 = P1_P1_INSTQUEUE_REG_1__4_ & n56373;
  assign n56564 = P1_P1_INSTQUEUE_REG_0__4_ & n56375;
  assign n56565 = ~n56561 & ~n56562;
  assign n56566 = ~n56563 & n56565;
  assign n56567 = ~n56564 & n56566;
  assign n56568 = P1_P1_INSTQUEUE_REG_15__4_ & n56381;
  assign n56569 = P1_P1_INSTQUEUE_REG_14__4_ & n56383;
  assign n56570 = P1_P1_INSTQUEUE_REG_13__4_ & n56385;
  assign n56571 = P1_P1_INSTQUEUE_REG_12__4_ & n56387;
  assign n56572 = ~n56568 & ~n56569;
  assign n56573 = ~n56570 & n56572;
  assign n56574 = ~n56571 & n56573;
  assign n56575 = P1_P1_INSTQUEUE_REG_11__4_ & n56393;
  assign n56576 = P1_P1_INSTQUEUE_REG_10__4_ & n56395;
  assign n56577 = P1_P1_INSTQUEUE_REG_9__4_ & n56397;
  assign n56578 = P1_P1_INSTQUEUE_REG_8__4_ & n56399;
  assign n56579 = ~n56575 & ~n56576;
  assign n56580 = ~n56577 & n56579;
  assign n56581 = ~n56578 & n56580;
  assign n56582 = n56560 & n56567;
  assign n56583 = n56574 & n56582;
  assign n56584 = n56581 & n56583;
  assign n56585 = n55907 & ~n56584;
  assign n56586 = ~n50294 & n56408;
  assign n56587 = P1_P1_EAX_REG_20_ & ~n55906;
  assign n56588 = P1_P1_EAX_REG_19_ & n56544;
  assign n56589 = ~P1_P1_EAX_REG_20_ & n56588;
  assign n56590 = P1_P1_EAX_REG_20_ & ~n56588;
  assign n56591 = ~n56589 & ~n56590;
  assign n56592 = n55913 & ~n56591;
  assign n56593 = ~n56587 & ~n56592;
  assign n56594 = ~n50309 & n56417;
  assign n56595 = ~n56585 & ~n56586;
  assign n56596 = n56593 & n56595;
  assign n9531 = n56594 | ~n56596;
  assign n56598 = P1_P1_INSTQUEUE_REG_7__5_ & n56357;
  assign n56599 = P1_P1_INSTQUEUE_REG_6__5_ & n56359;
  assign n56600 = P1_P1_INSTQUEUE_REG_5__5_ & n56361;
  assign n56601 = P1_P1_INSTQUEUE_REG_4__5_ & n56363;
  assign n56602 = ~n56598 & ~n56599;
  assign n56603 = ~n56600 & n56602;
  assign n56604 = ~n56601 & n56603;
  assign n56605 = P1_P1_INSTQUEUE_REG_3__5_ & n56369;
  assign n56606 = P1_P1_INSTQUEUE_REG_2__5_ & n56371;
  assign n56607 = P1_P1_INSTQUEUE_REG_1__5_ & n56373;
  assign n56608 = P1_P1_INSTQUEUE_REG_0__5_ & n56375;
  assign n56609 = ~n56605 & ~n56606;
  assign n56610 = ~n56607 & n56609;
  assign n56611 = ~n56608 & n56610;
  assign n56612 = P1_P1_INSTQUEUE_REG_15__5_ & n56381;
  assign n56613 = P1_P1_INSTQUEUE_REG_14__5_ & n56383;
  assign n56614 = P1_P1_INSTQUEUE_REG_13__5_ & n56385;
  assign n56615 = P1_P1_INSTQUEUE_REG_12__5_ & n56387;
  assign n56616 = ~n56612 & ~n56613;
  assign n56617 = ~n56614 & n56616;
  assign n56618 = ~n56615 & n56617;
  assign n56619 = P1_P1_INSTQUEUE_REG_11__5_ & n56393;
  assign n56620 = P1_P1_INSTQUEUE_REG_10__5_ & n56395;
  assign n56621 = P1_P1_INSTQUEUE_REG_9__5_ & n56397;
  assign n56622 = P1_P1_INSTQUEUE_REG_8__5_ & n56399;
  assign n56623 = ~n56619 & ~n56620;
  assign n56624 = ~n56621 & n56623;
  assign n56625 = ~n56622 & n56624;
  assign n56626 = n56604 & n56611;
  assign n56627 = n56618 & n56626;
  assign n56628 = n56625 & n56627;
  assign n56629 = n55907 & ~n56628;
  assign n56630 = ~n50250 & n56408;
  assign n56631 = P1_P1_EAX_REG_21_ & ~n55906;
  assign n56632 = P1_P1_EAX_REG_20_ & n56588;
  assign n56633 = ~P1_P1_EAX_REG_21_ & n56632;
  assign n56634 = P1_P1_EAX_REG_21_ & ~n56632;
  assign n56635 = ~n56633 & ~n56634;
  assign n56636 = n55913 & ~n56635;
  assign n56637 = ~n56631 & ~n56636;
  assign n56638 = ~n50263 & n56417;
  assign n56639 = ~n56629 & ~n56630;
  assign n56640 = n56637 & n56639;
  assign n9536 = n56638 | ~n56640;
  assign n56642 = P1_P1_EAX_REG_22_ & ~n55906;
  assign n56643 = P1_P1_EAX_REG_21_ & n56632;
  assign n56644 = ~P1_P1_EAX_REG_22_ & n56643;
  assign n56645 = P1_P1_EAX_REG_22_ & ~n56643;
  assign n56646 = ~n56644 & ~n56645;
  assign n56647 = n55913 & ~n56646;
  assign n56648 = P1_P1_INSTQUEUE_REG_7__6_ & n56357;
  assign n56649 = P1_P1_INSTQUEUE_REG_6__6_ & n56359;
  assign n56650 = P1_P1_INSTQUEUE_REG_5__6_ & n56361;
  assign n56651 = P1_P1_INSTQUEUE_REG_4__6_ & n56363;
  assign n56652 = ~n56648 & ~n56649;
  assign n56653 = ~n56650 & n56652;
  assign n56654 = ~n56651 & n56653;
  assign n56655 = P1_P1_INSTQUEUE_REG_3__6_ & n56369;
  assign n56656 = P1_P1_INSTQUEUE_REG_2__6_ & n56371;
  assign n56657 = P1_P1_INSTQUEUE_REG_1__6_ & n56373;
  assign n56658 = P1_P1_INSTQUEUE_REG_0__6_ & n56375;
  assign n56659 = ~n56655 & ~n56656;
  assign n56660 = ~n56657 & n56659;
  assign n56661 = ~n56658 & n56660;
  assign n56662 = P1_P1_INSTQUEUE_REG_15__6_ & n56381;
  assign n56663 = P1_P1_INSTQUEUE_REG_14__6_ & n56383;
  assign n56664 = P1_P1_INSTQUEUE_REG_13__6_ & n56385;
  assign n56665 = P1_P1_INSTQUEUE_REG_12__6_ & n56387;
  assign n56666 = ~n56662 & ~n56663;
  assign n56667 = ~n56664 & n56666;
  assign n56668 = ~n56665 & n56667;
  assign n56669 = P1_P1_INSTQUEUE_REG_11__6_ & n56393;
  assign n56670 = P1_P1_INSTQUEUE_REG_10__6_ & n56395;
  assign n56671 = P1_P1_INSTQUEUE_REG_9__6_ & n56397;
  assign n56672 = P1_P1_INSTQUEUE_REG_8__6_ & n56399;
  assign n56673 = ~n56669 & ~n56670;
  assign n56674 = ~n56671 & n56673;
  assign n56675 = ~n56672 & n56674;
  assign n56676 = n56654 & n56661;
  assign n56677 = n56668 & n56676;
  assign n56678 = n56675 & n56677;
  assign n56679 = n55907 & ~n56678;
  assign n56680 = ~n56642 & ~n56647;
  assign n56681 = ~n56679 & n56680;
  assign n56682 = ~n50203 & n56408;
  assign n56683 = ~n50219 & n56417;
  assign n56684 = n56681 & ~n56682;
  assign n9541 = n56683 | ~n56684;
  assign n56686 = P1_P1_EAX_REG_23_ & ~n55906;
  assign n56687 = P1_P1_EAX_REG_22_ & n56643;
  assign n56688 = ~P1_P1_EAX_REG_23_ & n56687;
  assign n56689 = P1_P1_EAX_REG_23_ & ~n56687;
  assign n56690 = ~n56688 & ~n56689;
  assign n56691 = n55913 & ~n56690;
  assign n56692 = P1_P1_INSTQUEUERD_ADDR_REG_3_ & ~P1_P1_INSTQUEUERD_ADDR_REG_2_;
  assign n56693 = ~n43374 & ~n56692;
  assign n56694 = n43345 & n56693;
  assign n56695 = P1_P1_INSTQUEUE_REG_7__0_ & n56694;
  assign n56696 = n43349 & n56693;
  assign n56697 = P1_P1_INSTQUEUE_REG_6__0_ & n56696;
  assign n56698 = n43354 & n56693;
  assign n56699 = P1_P1_INSTQUEUE_REG_5__0_ & n56698;
  assign n56700 = n43358 & n56693;
  assign n56701 = P1_P1_INSTQUEUE_REG_4__0_ & n56700;
  assign n56702 = ~n56695 & ~n56697;
  assign n56703 = ~n56699 & n56702;
  assign n56704 = ~n56701 & n56703;
  assign n56705 = P1_P1_INSTQUEUERD_ADDR_REG_2_ & n56693;
  assign n56706 = n43344 & n56705;
  assign n56707 = P1_P1_INSTQUEUE_REG_3__0_ & n56706;
  assign n56708 = n43348 & n56705;
  assign n56709 = P1_P1_INSTQUEUE_REG_2__0_ & n56708;
  assign n56710 = n43353 & n56705;
  assign n56711 = P1_P1_INSTQUEUE_REG_1__0_ & n56710;
  assign n56712 = n43357 & n56705;
  assign n56713 = P1_P1_INSTQUEUE_REG_0__0_ & n56712;
  assign n56714 = ~n56707 & ~n56709;
  assign n56715 = ~n56711 & n56714;
  assign n56716 = ~n56713 & n56715;
  assign n56717 = n43345 & ~n56693;
  assign n56718 = P1_P1_INSTQUEUE_REG_15__0_ & n56717;
  assign n56719 = n43349 & ~n56693;
  assign n56720 = P1_P1_INSTQUEUE_REG_14__0_ & n56719;
  assign n56721 = n43354 & ~n56693;
  assign n56722 = P1_P1_INSTQUEUE_REG_13__0_ & n56721;
  assign n56723 = n43358 & ~n56693;
  assign n56724 = P1_P1_INSTQUEUE_REG_12__0_ & n56723;
  assign n56725 = ~n56718 & ~n56720;
  assign n56726 = ~n56722 & n56725;
  assign n56727 = ~n56724 & n56726;
  assign n56728 = P1_P1_INSTQUEUERD_ADDR_REG_2_ & ~n56693;
  assign n56729 = n43344 & n56728;
  assign n56730 = P1_P1_INSTQUEUE_REG_11__0_ & n56729;
  assign n56731 = n43348 & n56728;
  assign n56732 = P1_P1_INSTQUEUE_REG_10__0_ & n56731;
  assign n56733 = n43353 & n56728;
  assign n56734 = P1_P1_INSTQUEUE_REG_9__0_ & n56733;
  assign n56735 = n43357 & n56728;
  assign n56736 = P1_P1_INSTQUEUE_REG_8__0_ & n56735;
  assign n56737 = ~n56730 & ~n56732;
  assign n56738 = ~n56734 & n56737;
  assign n56739 = ~n56736 & n56738;
  assign n56740 = n56704 & n56716;
  assign n56741 = n56727 & n56740;
  assign n56742 = n56739 & n56741;
  assign n56743 = P1_P1_INSTQUEUE_REG_7__7_ & n56357;
  assign n56744 = P1_P1_INSTQUEUE_REG_6__7_ & n56359;
  assign n56745 = P1_P1_INSTQUEUE_REG_5__7_ & n56361;
  assign n56746 = P1_P1_INSTQUEUE_REG_4__7_ & n56363;
  assign n56747 = ~n56743 & ~n56744;
  assign n56748 = ~n56745 & n56747;
  assign n56749 = ~n56746 & n56748;
  assign n56750 = P1_P1_INSTQUEUE_REG_3__7_ & n56369;
  assign n56751 = P1_P1_INSTQUEUE_REG_2__7_ & n56371;
  assign n56752 = P1_P1_INSTQUEUE_REG_1__7_ & n56373;
  assign n56753 = P1_P1_INSTQUEUE_REG_0__7_ & n56375;
  assign n56754 = ~n56750 & ~n56751;
  assign n56755 = ~n56752 & n56754;
  assign n56756 = ~n56753 & n56755;
  assign n56757 = P1_P1_INSTQUEUE_REG_15__7_ & n56381;
  assign n56758 = P1_P1_INSTQUEUE_REG_14__7_ & n56383;
  assign n56759 = P1_P1_INSTQUEUE_REG_13__7_ & n56385;
  assign n56760 = P1_P1_INSTQUEUE_REG_12__7_ & n56387;
  assign n56761 = ~n56757 & ~n56758;
  assign n56762 = ~n56759 & n56761;
  assign n56763 = ~n56760 & n56762;
  assign n56764 = P1_P1_INSTQUEUE_REG_11__7_ & n56393;
  assign n56765 = P1_P1_INSTQUEUE_REG_10__7_ & n56395;
  assign n56766 = P1_P1_INSTQUEUE_REG_9__7_ & n56397;
  assign n56767 = P1_P1_INSTQUEUE_REG_8__7_ & n56399;
  assign n56768 = ~n56764 & ~n56765;
  assign n56769 = ~n56766 & n56768;
  assign n56770 = ~n56767 & n56769;
  assign n56771 = n56749 & n56756;
  assign n56772 = n56763 & n56771;
  assign n56773 = n56770 & n56772;
  assign n56774 = ~n56742 & n56773;
  assign n56775 = n56742 & ~n56773;
  assign n56776 = ~n56774 & ~n56775;
  assign n56777 = n55907 & ~n56776;
  assign n56778 = ~n56686 & ~n56691;
  assign n56779 = ~n56777 & n56778;
  assign n56780 = ~n44368 & n56408;
  assign n56781 = ~n47259 & n56417;
  assign n56782 = n56779 & ~n56780;
  assign n9546 = n56781 | ~n56782;
  assign n56784 = P1_P1_EAX_REG_24_ & ~n55906;
  assign n56785 = P1_P1_EAX_REG_23_ & n56687;
  assign n56786 = ~P1_P1_EAX_REG_24_ & n56785;
  assign n56787 = P1_P1_EAX_REG_24_ & ~n56785;
  assign n56788 = ~n56786 & ~n56787;
  assign n56789 = n55913 & ~n56788;
  assign n56790 = ~n56742 & ~n56773;
  assign n56791 = P1_P1_INSTQUEUE_REG_7__1_ & n56694;
  assign n56792 = P1_P1_INSTQUEUE_REG_6__1_ & n56696;
  assign n56793 = P1_P1_INSTQUEUE_REG_5__1_ & n56698;
  assign n56794 = P1_P1_INSTQUEUE_REG_4__1_ & n56700;
  assign n56795 = ~n56791 & ~n56792;
  assign n56796 = ~n56793 & n56795;
  assign n56797 = ~n56794 & n56796;
  assign n56798 = P1_P1_INSTQUEUE_REG_3__1_ & n56706;
  assign n56799 = P1_P1_INSTQUEUE_REG_2__1_ & n56708;
  assign n56800 = P1_P1_INSTQUEUE_REG_1__1_ & n56710;
  assign n56801 = P1_P1_INSTQUEUE_REG_0__1_ & n56712;
  assign n56802 = ~n56798 & ~n56799;
  assign n56803 = ~n56800 & n56802;
  assign n56804 = ~n56801 & n56803;
  assign n56805 = P1_P1_INSTQUEUE_REG_15__1_ & n56717;
  assign n56806 = P1_P1_INSTQUEUE_REG_14__1_ & n56719;
  assign n56807 = P1_P1_INSTQUEUE_REG_13__1_ & n56721;
  assign n56808 = P1_P1_INSTQUEUE_REG_12__1_ & n56723;
  assign n56809 = ~n56805 & ~n56806;
  assign n56810 = ~n56807 & n56809;
  assign n56811 = ~n56808 & n56810;
  assign n56812 = P1_P1_INSTQUEUE_REG_11__1_ & n56729;
  assign n56813 = P1_P1_INSTQUEUE_REG_10__1_ & n56731;
  assign n56814 = P1_P1_INSTQUEUE_REG_9__1_ & n56733;
  assign n56815 = P1_P1_INSTQUEUE_REG_8__1_ & n56735;
  assign n56816 = ~n56812 & ~n56813;
  assign n56817 = ~n56814 & n56816;
  assign n56818 = ~n56815 & n56817;
  assign n56819 = n56797 & n56804;
  assign n56820 = n56811 & n56819;
  assign n56821 = n56818 & n56820;
  assign n56822 = n56790 & n56821;
  assign n56823 = ~n56790 & ~n56821;
  assign n56824 = ~n56822 & ~n56823;
  assign n56825 = n55907 & ~n56824;
  assign n56826 = ~n56784 & ~n56789;
  assign n56827 = ~n56825 & n56826;
  assign n56828 = ~n55638 & n56408;
  assign n56829 = ~n50487 & n56417;
  assign n56830 = n56827 & ~n56828;
  assign n9551 = n56829 | ~n56830;
  assign n56832 = P1_P1_EAX_REG_25_ & ~n55906;
  assign n56833 = P1_P1_EAX_REG_24_ & n56785;
  assign n56834 = ~P1_P1_EAX_REG_25_ & n56833;
  assign n56835 = P1_P1_EAX_REG_25_ & ~n56833;
  assign n56836 = ~n56834 & ~n56835;
  assign n56837 = n55913 & ~n56836;
  assign n56838 = n56790 & ~n56821;
  assign n56839 = P1_P1_INSTQUEUE_REG_7__2_ & n56694;
  assign n56840 = P1_P1_INSTQUEUE_REG_6__2_ & n56696;
  assign n56841 = P1_P1_INSTQUEUE_REG_5__2_ & n56698;
  assign n56842 = P1_P1_INSTQUEUE_REG_4__2_ & n56700;
  assign n56843 = ~n56839 & ~n56840;
  assign n56844 = ~n56841 & n56843;
  assign n56845 = ~n56842 & n56844;
  assign n56846 = P1_P1_INSTQUEUE_REG_3__2_ & n56706;
  assign n56847 = P1_P1_INSTQUEUE_REG_2__2_ & n56708;
  assign n56848 = P1_P1_INSTQUEUE_REG_1__2_ & n56710;
  assign n56849 = P1_P1_INSTQUEUE_REG_0__2_ & n56712;
  assign n56850 = ~n56846 & ~n56847;
  assign n56851 = ~n56848 & n56850;
  assign n56852 = ~n56849 & n56851;
  assign n56853 = P1_P1_INSTQUEUE_REG_15__2_ & n56717;
  assign n56854 = P1_P1_INSTQUEUE_REG_14__2_ & n56719;
  assign n56855 = P1_P1_INSTQUEUE_REG_13__2_ & n56721;
  assign n56856 = P1_P1_INSTQUEUE_REG_12__2_ & n56723;
  assign n56857 = ~n56853 & ~n56854;
  assign n56858 = ~n56855 & n56857;
  assign n56859 = ~n56856 & n56858;
  assign n56860 = P1_P1_INSTQUEUE_REG_11__2_ & n56729;
  assign n56861 = P1_P1_INSTQUEUE_REG_10__2_ & n56731;
  assign n56862 = P1_P1_INSTQUEUE_REG_9__2_ & n56733;
  assign n56863 = P1_P1_INSTQUEUE_REG_8__2_ & n56735;
  assign n56864 = ~n56860 & ~n56861;
  assign n56865 = ~n56862 & n56864;
  assign n56866 = ~n56863 & n56865;
  assign n56867 = n56845 & n56852;
  assign n56868 = n56859 & n56867;
  assign n56869 = n56866 & n56868;
  assign n56870 = n56838 & n56869;
  assign n56871 = ~n56838 & ~n56869;
  assign n56872 = ~n56870 & ~n56871;
  assign n56873 = n55907 & ~n56872;
  assign n56874 = ~n56832 & ~n56837;
  assign n56875 = ~n56873 & n56874;
  assign n56876 = ~n55621 & n56408;
  assign n56877 = ~n50448 & n56417;
  assign n56878 = n56875 & ~n56876;
  assign n9556 = n56877 | ~n56878;
  assign n56880 = P1_P1_EAX_REG_26_ & ~n55906;
  assign n56881 = P1_P1_EAX_REG_25_ & n56833;
  assign n56882 = ~P1_P1_EAX_REG_26_ & n56881;
  assign n56883 = P1_P1_EAX_REG_26_ & ~n56881;
  assign n56884 = ~n56882 & ~n56883;
  assign n56885 = n55913 & ~n56884;
  assign n56886 = n56838 & ~n56869;
  assign n56887 = P1_P1_INSTQUEUE_REG_7__3_ & n56694;
  assign n56888 = P1_P1_INSTQUEUE_REG_6__3_ & n56696;
  assign n56889 = P1_P1_INSTQUEUE_REG_5__3_ & n56698;
  assign n56890 = P1_P1_INSTQUEUE_REG_4__3_ & n56700;
  assign n56891 = ~n56887 & ~n56888;
  assign n56892 = ~n56889 & n56891;
  assign n56893 = ~n56890 & n56892;
  assign n56894 = P1_P1_INSTQUEUE_REG_3__3_ & n56706;
  assign n56895 = P1_P1_INSTQUEUE_REG_2__3_ & n56708;
  assign n56896 = P1_P1_INSTQUEUE_REG_1__3_ & n56710;
  assign n56897 = P1_P1_INSTQUEUE_REG_0__3_ & n56712;
  assign n56898 = ~n56894 & ~n56895;
  assign n56899 = ~n56896 & n56898;
  assign n56900 = ~n56897 & n56899;
  assign n56901 = P1_P1_INSTQUEUE_REG_15__3_ & n56717;
  assign n56902 = P1_P1_INSTQUEUE_REG_14__3_ & n56719;
  assign n56903 = P1_P1_INSTQUEUE_REG_13__3_ & n56721;
  assign n56904 = P1_P1_INSTQUEUE_REG_12__3_ & n56723;
  assign n56905 = ~n56901 & ~n56902;
  assign n56906 = ~n56903 & n56905;
  assign n56907 = ~n56904 & n56906;
  assign n56908 = P1_P1_INSTQUEUE_REG_11__3_ & n56729;
  assign n56909 = P1_P1_INSTQUEUE_REG_10__3_ & n56731;
  assign n56910 = P1_P1_INSTQUEUE_REG_9__3_ & n56733;
  assign n56911 = P1_P1_INSTQUEUE_REG_8__3_ & n56735;
  assign n56912 = ~n56908 & ~n56909;
  assign n56913 = ~n56910 & n56912;
  assign n56914 = ~n56911 & n56913;
  assign n56915 = n56893 & n56900;
  assign n56916 = n56907 & n56915;
  assign n56917 = n56914 & n56916;
  assign n56918 = n56886 & n56917;
  assign n56919 = ~n56886 & ~n56917;
  assign n56920 = ~n56918 & ~n56919;
  assign n56921 = n55907 & ~n56920;
  assign n56922 = ~n56880 & ~n56885;
  assign n56923 = ~n56921 & n56922;
  assign n56924 = ~n55609 & n56408;
  assign n56925 = ~n50410 & n56417;
  assign n56926 = n56923 & ~n56924;
  assign n9561 = n56925 | ~n56926;
  assign n56928 = P1_P1_EAX_REG_27_ & ~n55906;
  assign n56929 = P1_P1_EAX_REG_26_ & n56881;
  assign n56930 = ~P1_P1_EAX_REG_27_ & n56929;
  assign n56931 = P1_P1_EAX_REG_27_ & ~n56929;
  assign n56932 = ~n56930 & ~n56931;
  assign n56933 = n55913 & ~n56932;
  assign n56934 = n56886 & ~n56917;
  assign n56935 = P1_P1_INSTQUEUE_REG_7__4_ & n56694;
  assign n56936 = P1_P1_INSTQUEUE_REG_6__4_ & n56696;
  assign n56937 = P1_P1_INSTQUEUE_REG_5__4_ & n56698;
  assign n56938 = P1_P1_INSTQUEUE_REG_4__4_ & n56700;
  assign n56939 = ~n56935 & ~n56936;
  assign n56940 = ~n56937 & n56939;
  assign n56941 = ~n56938 & n56940;
  assign n56942 = P1_P1_INSTQUEUE_REG_3__4_ & n56706;
  assign n56943 = P1_P1_INSTQUEUE_REG_2__4_ & n56708;
  assign n56944 = P1_P1_INSTQUEUE_REG_1__4_ & n56710;
  assign n56945 = P1_P1_INSTQUEUE_REG_0__4_ & n56712;
  assign n56946 = ~n56942 & ~n56943;
  assign n56947 = ~n56944 & n56946;
  assign n56948 = ~n56945 & n56947;
  assign n56949 = P1_P1_INSTQUEUE_REG_15__4_ & n56717;
  assign n56950 = P1_P1_INSTQUEUE_REG_14__4_ & n56719;
  assign n56951 = P1_P1_INSTQUEUE_REG_13__4_ & n56721;
  assign n56952 = P1_P1_INSTQUEUE_REG_12__4_ & n56723;
  assign n56953 = ~n56949 & ~n56950;
  assign n56954 = ~n56951 & n56953;
  assign n56955 = ~n56952 & n56954;
  assign n56956 = P1_P1_INSTQUEUE_REG_11__4_ & n56729;
  assign n56957 = P1_P1_INSTQUEUE_REG_10__4_ & n56731;
  assign n56958 = P1_P1_INSTQUEUE_REG_9__4_ & n56733;
  assign n56959 = P1_P1_INSTQUEUE_REG_8__4_ & n56735;
  assign n56960 = ~n56956 & ~n56957;
  assign n56961 = ~n56958 & n56960;
  assign n56962 = ~n56959 & n56961;
  assign n56963 = n56941 & n56948;
  assign n56964 = n56955 & n56963;
  assign n56965 = n56962 & n56964;
  assign n56966 = n56934 & n56965;
  assign n56967 = ~n56934 & ~n56965;
  assign n56968 = ~n56966 & ~n56967;
  assign n56969 = n55907 & ~n56968;
  assign n56970 = ~n56928 & ~n56933;
  assign n56971 = ~n56969 & n56970;
  assign n56972 = ~n55593 & n56408;
  assign n56973 = ~n50362 & n56417;
  assign n56974 = n56971 & ~n56972;
  assign n9566 = n56973 | ~n56974;
  assign n56976 = P1_P1_EAX_REG_28_ & ~n55906;
  assign n56977 = P1_P1_EAX_REG_27_ & n56929;
  assign n56978 = ~P1_P1_EAX_REG_28_ & n56977;
  assign n56979 = P1_P1_EAX_REG_28_ & ~n56977;
  assign n56980 = ~n56978 & ~n56979;
  assign n56981 = n55913 & ~n56980;
  assign n56982 = n56934 & ~n56965;
  assign n56983 = P1_P1_INSTQUEUE_REG_7__5_ & n56694;
  assign n56984 = P1_P1_INSTQUEUE_REG_6__5_ & n56696;
  assign n56985 = P1_P1_INSTQUEUE_REG_5__5_ & n56698;
  assign n56986 = P1_P1_INSTQUEUE_REG_4__5_ & n56700;
  assign n56987 = ~n56983 & ~n56984;
  assign n56988 = ~n56985 & n56987;
  assign n56989 = ~n56986 & n56988;
  assign n56990 = P1_P1_INSTQUEUE_REG_3__5_ & n56706;
  assign n56991 = P1_P1_INSTQUEUE_REG_2__5_ & n56708;
  assign n56992 = P1_P1_INSTQUEUE_REG_1__5_ & n56710;
  assign n56993 = P1_P1_INSTQUEUE_REG_0__5_ & n56712;
  assign n56994 = ~n56990 & ~n56991;
  assign n56995 = ~n56992 & n56994;
  assign n56996 = ~n56993 & n56995;
  assign n56997 = P1_P1_INSTQUEUE_REG_15__5_ & n56717;
  assign n56998 = P1_P1_INSTQUEUE_REG_14__5_ & n56719;
  assign n56999 = P1_P1_INSTQUEUE_REG_13__5_ & n56721;
  assign n57000 = P1_P1_INSTQUEUE_REG_12__5_ & n56723;
  assign n57001 = ~n56997 & ~n56998;
  assign n57002 = ~n56999 & n57001;
  assign n57003 = ~n57000 & n57002;
  assign n57004 = P1_P1_INSTQUEUE_REG_11__5_ & n56729;
  assign n57005 = P1_P1_INSTQUEUE_REG_10__5_ & n56731;
  assign n57006 = P1_P1_INSTQUEUE_REG_9__5_ & n56733;
  assign n57007 = P1_P1_INSTQUEUE_REG_8__5_ & n56735;
  assign n57008 = ~n57004 & ~n57005;
  assign n57009 = ~n57006 & n57008;
  assign n57010 = ~n57007 & n57009;
  assign n57011 = n56989 & n56996;
  assign n57012 = n57003 & n57011;
  assign n57013 = n57010 & n57012;
  assign n57014 = n56982 & n57013;
  assign n57015 = ~n56982 & ~n57013;
  assign n57016 = ~n57014 & ~n57015;
  assign n57017 = n55907 & ~n57016;
  assign n57018 = ~n56976 & ~n56981;
  assign n57019 = ~n57017 & n57018;
  assign n57020 = ~n55578 & n56408;
  assign n57021 = ~n50321 & n56417;
  assign n57022 = n57019 & ~n57020;
  assign n9571 = n57021 | ~n57022;
  assign n57024 = P1_P1_EAX_REG_29_ & ~n55906;
  assign n57025 = P1_P1_EAX_REG_28_ & n56977;
  assign n57026 = ~P1_P1_EAX_REG_29_ & n57025;
  assign n57027 = P1_P1_EAX_REG_29_ & ~n57025;
  assign n57028 = ~n57026 & ~n57027;
  assign n57029 = n55913 & ~n57028;
  assign n57030 = n56982 & ~n57013;
  assign n57031 = P1_P1_INSTQUEUE_REG_7__6_ & n56694;
  assign n57032 = P1_P1_INSTQUEUE_REG_6__6_ & n56696;
  assign n57033 = P1_P1_INSTQUEUE_REG_5__6_ & n56698;
  assign n57034 = P1_P1_INSTQUEUE_REG_4__6_ & n56700;
  assign n57035 = ~n57031 & ~n57032;
  assign n57036 = ~n57033 & n57035;
  assign n57037 = ~n57034 & n57036;
  assign n57038 = P1_P1_INSTQUEUE_REG_3__6_ & n56706;
  assign n57039 = P1_P1_INSTQUEUE_REG_2__6_ & n56708;
  assign n57040 = P1_P1_INSTQUEUE_REG_1__6_ & n56710;
  assign n57041 = P1_P1_INSTQUEUE_REG_0__6_ & n56712;
  assign n57042 = ~n57038 & ~n57039;
  assign n57043 = ~n57040 & n57042;
  assign n57044 = ~n57041 & n57043;
  assign n57045 = P1_P1_INSTQUEUE_REG_15__6_ & n56717;
  assign n57046 = P1_P1_INSTQUEUE_REG_14__6_ & n56719;
  assign n57047 = P1_P1_INSTQUEUE_REG_13__6_ & n56721;
  assign n57048 = P1_P1_INSTQUEUE_REG_12__6_ & n56723;
  assign n57049 = ~n57045 & ~n57046;
  assign n57050 = ~n57047 & n57049;
  assign n57051 = ~n57048 & n57050;
  assign n57052 = P1_P1_INSTQUEUE_REG_11__6_ & n56729;
  assign n57053 = P1_P1_INSTQUEUE_REG_10__6_ & n56731;
  assign n57054 = P1_P1_INSTQUEUE_REG_9__6_ & n56733;
  assign n57055 = P1_P1_INSTQUEUE_REG_8__6_ & n56735;
  assign n57056 = ~n57052 & ~n57053;
  assign n57057 = ~n57054 & n57056;
  assign n57058 = ~n57055 & n57057;
  assign n57059 = n57037 & n57044;
  assign n57060 = n57051 & n57059;
  assign n57061 = n57058 & n57060;
  assign n57062 = n57030 & n57061;
  assign n57063 = ~n57030 & ~n57061;
  assign n57064 = ~n57062 & ~n57063;
  assign n57065 = n55907 & ~n57064;
  assign n57066 = ~n57024 & ~n57029;
  assign n57067 = ~n57065 & n57066;
  assign n57068 = ~n55562 & n56408;
  assign n57069 = ~n50275 & n56417;
  assign n57070 = n57067 & ~n57068;
  assign n9576 = n57069 | ~n57070;
  assign n57072 = P1_P1_EAX_REG_30_ & ~n55906;
  assign n57073 = P1_P1_EAX_REG_29_ & n57025;
  assign n57074 = ~P1_P1_EAX_REG_30_ & n57073;
  assign n57075 = P1_P1_EAX_REG_30_ & ~n57073;
  assign n57076 = ~n57074 & ~n57075;
  assign n57077 = n55913 & ~n57076;
  assign n57078 = n57030 & ~n57061;
  assign n57079 = P1_P1_INSTQUEUE_REG_7__7_ & n56694;
  assign n57080 = P1_P1_INSTQUEUE_REG_6__7_ & n56696;
  assign n57081 = P1_P1_INSTQUEUE_REG_5__7_ & n56698;
  assign n57082 = P1_P1_INSTQUEUE_REG_4__7_ & n56700;
  assign n57083 = ~n57079 & ~n57080;
  assign n57084 = ~n57081 & n57083;
  assign n57085 = ~n57082 & n57084;
  assign n57086 = P1_P1_INSTQUEUE_REG_3__7_ & n56706;
  assign n57087 = P1_P1_INSTQUEUE_REG_2__7_ & n56708;
  assign n57088 = P1_P1_INSTQUEUE_REG_1__7_ & n56710;
  assign n57089 = P1_P1_INSTQUEUE_REG_0__7_ & n56712;
  assign n57090 = ~n57086 & ~n57087;
  assign n57091 = ~n57088 & n57090;
  assign n57092 = ~n57089 & n57091;
  assign n57093 = P1_P1_INSTQUEUE_REG_15__7_ & n56717;
  assign n57094 = P1_P1_INSTQUEUE_REG_14__7_ & n56719;
  assign n57095 = P1_P1_INSTQUEUE_REG_13__7_ & n56721;
  assign n57096 = P1_P1_INSTQUEUE_REG_12__7_ & n56723;
  assign n57097 = ~n57093 & ~n57094;
  assign n57098 = ~n57095 & n57097;
  assign n57099 = ~n57096 & n57098;
  assign n57100 = P1_P1_INSTQUEUE_REG_11__7_ & n56729;
  assign n57101 = P1_P1_INSTQUEUE_REG_10__7_ & n56731;
  assign n57102 = P1_P1_INSTQUEUE_REG_9__7_ & n56733;
  assign n57103 = P1_P1_INSTQUEUE_REG_8__7_ & n56735;
  assign n57104 = ~n57100 & ~n57101;
  assign n57105 = ~n57102 & n57104;
  assign n57106 = ~n57103 & n57105;
  assign n57107 = n57085 & n57092;
  assign n57108 = n57099 & n57107;
  assign n57109 = n57106 & n57108;
  assign n57110 = n57078 & n57109;
  assign n57111 = ~n57078 & ~n57109;
  assign n57112 = ~n57110 & ~n57111;
  assign n57113 = n55907 & ~n57112;
  assign n57114 = ~n57072 & ~n57077;
  assign n57115 = ~n57113 & n57114;
  assign n57116 = ~n55548 & n56408;
  assign n57117 = ~n50233 & n56417;
  assign n57118 = n57115 & ~n57116;
  assign n9581 = n57117 | ~n57118;
  assign n57120 = P1_P1_EAX_REG_30_ & n57073;
  assign n57121 = ~P1_P1_EAX_REG_31_ & n57120;
  assign n57122 = P1_P1_EAX_REG_31_ & ~n57120;
  assign n57123 = ~n57121 & ~n57122;
  assign n57124 = n55913 & ~n57123;
  assign n57125 = P1_P1_EAX_REG_31_ & ~n55906;
  assign n57126 = ~n57124 & ~n57125;
  assign n57127 = ~n50186 & n56417;
  assign n9586 = ~n57126 | n57127;
  assign n57129 = ~n43765 & ~n43859;
  assign n57130 = n43979 & ~n57129;
  assign n57131 = n43495 & n57130;
  assign n57132 = ~P1_P1_EBX_REG_0_ & n57131;
  assign n57133 = ~n43495 & n57130;
  assign n57134 = P1_P1_INSTQUEUE_REG_0__0_ & n57133;
  assign n57135 = P1_P1_EBX_REG_0_ & ~n57130;
  assign n57136 = ~n57132 & ~n57134;
  assign n9591 = n57135 | ~n57136;
  assign n57138 = ~P1_P1_EBX_REG_0_ & P1_P1_EBX_REG_1_;
  assign n57139 = P1_P1_EBX_REG_0_ & ~P1_P1_EBX_REG_1_;
  assign n57140 = ~n57138 & ~n57139;
  assign n57141 = n57131 & ~n57140;
  assign n57142 = P1_P1_INSTQUEUE_REG_0__1_ & n57133;
  assign n57143 = P1_P1_EBX_REG_1_ & ~n57130;
  assign n57144 = ~n57141 & ~n57142;
  assign n9596 = n57143 | ~n57144;
  assign n57146 = P1_P1_EBX_REG_0_ & P1_P1_EBX_REG_1_;
  assign n57147 = ~P1_P1_EBX_REG_2_ & n57146;
  assign n57148 = P1_P1_EBX_REG_2_ & ~n57146;
  assign n57149 = ~n57147 & ~n57148;
  assign n57150 = n57131 & ~n57149;
  assign n57151 = P1_P1_INSTQUEUE_REG_0__2_ & n57133;
  assign n57152 = P1_P1_EBX_REG_2_ & ~n57130;
  assign n57153 = ~n57150 & ~n57151;
  assign n9601 = n57152 | ~n57153;
  assign n57155 = P1_P1_EBX_REG_0_ & P1_P1_EBX_REG_2_;
  assign n57156 = P1_P1_EBX_REG_1_ & n57155;
  assign n57157 = P1_P1_EBX_REG_3_ & ~n57156;
  assign n57158 = ~P1_P1_EBX_REG_3_ & n57156;
  assign n57159 = ~n57157 & ~n57158;
  assign n57160 = n57131 & ~n57159;
  assign n57161 = P1_P1_INSTQUEUE_REG_0__3_ & n57133;
  assign n57162 = P1_P1_EBX_REG_3_ & ~n57130;
  assign n57163 = ~n57160 & ~n57161;
  assign n9606 = n57162 | ~n57163;
  assign n57165 = P1_P1_EBX_REG_3_ & n57156;
  assign n57166 = ~P1_P1_EBX_REG_4_ & n57165;
  assign n57167 = P1_P1_EBX_REG_4_ & ~n57165;
  assign n57168 = ~n57166 & ~n57167;
  assign n57169 = n57131 & ~n57168;
  assign n57170 = P1_P1_INSTQUEUE_REG_0__4_ & n57133;
  assign n57171 = P1_P1_EBX_REG_4_ & ~n57130;
  assign n57172 = ~n57169 & ~n57170;
  assign n9611 = n57171 | ~n57172;
  assign n57174 = P1_P1_EBX_REG_3_ & P1_P1_EBX_REG_4_;
  assign n57175 = n57156 & n57174;
  assign n57176 = P1_P1_EBX_REG_5_ & ~n57175;
  assign n57177 = ~P1_P1_EBX_REG_5_ & n57175;
  assign n57178 = ~n57176 & ~n57177;
  assign n57179 = n57131 & ~n57178;
  assign n57180 = P1_P1_INSTQUEUE_REG_0__5_ & n57133;
  assign n57181 = P1_P1_EBX_REG_5_ & ~n57130;
  assign n57182 = ~n57179 & ~n57180;
  assign n9616 = n57181 | ~n57182;
  assign n57184 = P1_P1_EBX_REG_5_ & n57175;
  assign n57185 = ~P1_P1_EBX_REG_6_ & n57184;
  assign n57186 = P1_P1_EBX_REG_6_ & ~n57184;
  assign n57187 = ~n57185 & ~n57186;
  assign n57188 = n57131 & ~n57187;
  assign n57189 = P1_P1_INSTQUEUE_REG_0__6_ & n57133;
  assign n57190 = P1_P1_EBX_REG_6_ & ~n57130;
  assign n57191 = ~n57188 & ~n57189;
  assign n9621 = n57190 | ~n57191;
  assign n57193 = P1_P1_EBX_REG_5_ & P1_P1_EBX_REG_6_;
  assign n57194 = n57175 & n57193;
  assign n57195 = P1_P1_EBX_REG_7_ & ~n57194;
  assign n57196 = ~P1_P1_EBX_REG_7_ & n57194;
  assign n57197 = ~n57195 & ~n57196;
  assign n57198 = n57131 & ~n57197;
  assign n57199 = P1_P1_INSTQUEUE_REG_0__7_ & n57133;
  assign n57200 = P1_P1_EBX_REG_7_ & ~n57130;
  assign n57201 = ~n57198 & ~n57199;
  assign n9626 = n57200 | ~n57201;
  assign n57203 = P1_P1_EBX_REG_7_ & n57194;
  assign n57204 = ~P1_P1_EBX_REG_8_ & n57203;
  assign n57205 = P1_P1_EBX_REG_8_ & ~n57203;
  assign n57206 = ~n57204 & ~n57205;
  assign n57207 = n57131 & ~n57206;
  assign n57208 = ~n56052 & n57133;
  assign n57209 = P1_P1_EBX_REG_8_ & ~n57130;
  assign n57210 = ~n57207 & ~n57208;
  assign n9631 = n57209 | ~n57210;
  assign n57212 = P1_P1_EBX_REG_7_ & P1_P1_EBX_REG_8_;
  assign n57213 = n57194 & n57212;
  assign n57214 = P1_P1_EBX_REG_9_ & ~n57213;
  assign n57215 = ~P1_P1_EBX_REG_9_ & n57213;
  assign n57216 = ~n57214 & ~n57215;
  assign n57217 = n57131 & ~n57216;
  assign n57218 = ~n56094 & n57133;
  assign n57219 = P1_P1_EBX_REG_9_ & ~n57130;
  assign n57220 = ~n57217 & ~n57218;
  assign n9636 = n57219 | ~n57220;
  assign n57222 = P1_P1_EBX_REG_9_ & n57213;
  assign n57223 = ~P1_P1_EBX_REG_10_ & n57222;
  assign n57224 = P1_P1_EBX_REG_10_ & ~n57222;
  assign n57225 = ~n57223 & ~n57224;
  assign n57226 = n57131 & ~n57225;
  assign n57227 = ~n56136 & n57133;
  assign n57228 = P1_P1_EBX_REG_10_ & ~n57130;
  assign n57229 = ~n57226 & ~n57227;
  assign n9641 = n57228 | ~n57229;
  assign n57231 = P1_P1_EBX_REG_9_ & P1_P1_EBX_REG_10_;
  assign n57232 = n57213 & n57231;
  assign n57233 = P1_P1_EBX_REG_11_ & ~n57232;
  assign n57234 = ~P1_P1_EBX_REG_11_ & n57232;
  assign n57235 = ~n57233 & ~n57234;
  assign n57236 = n57131 & ~n57235;
  assign n57237 = ~n56178 & n57133;
  assign n57238 = P1_P1_EBX_REG_11_ & ~n57130;
  assign n57239 = ~n57236 & ~n57237;
  assign n9646 = n57238 | ~n57239;
  assign n57241 = P1_P1_EBX_REG_11_ & n57232;
  assign n57242 = ~P1_P1_EBX_REG_12_ & n57241;
  assign n57243 = P1_P1_EBX_REG_12_ & ~n57241;
  assign n57244 = ~n57242 & ~n57243;
  assign n57245 = n57131 & ~n57244;
  assign n57246 = ~n56220 & n57133;
  assign n57247 = P1_P1_EBX_REG_12_ & ~n57130;
  assign n57248 = ~n57245 & ~n57246;
  assign n9651 = n57247 | ~n57248;
  assign n57250 = P1_P1_EBX_REG_11_ & P1_P1_EBX_REG_12_;
  assign n57251 = n57232 & n57250;
  assign n57252 = P1_P1_EBX_REG_13_ & ~n57251;
  assign n57253 = ~P1_P1_EBX_REG_13_ & n57251;
  assign n57254 = ~n57252 & ~n57253;
  assign n57255 = n57131 & ~n57254;
  assign n57256 = ~n56262 & n57133;
  assign n57257 = P1_P1_EBX_REG_13_ & ~n57130;
  assign n57258 = ~n57255 & ~n57256;
  assign n9656 = n57257 | ~n57258;
  assign n57260 = P1_P1_EBX_REG_13_ & n57251;
  assign n57261 = ~P1_P1_EBX_REG_14_ & n57260;
  assign n57262 = P1_P1_EBX_REG_14_ & ~n57260;
  assign n57263 = ~n57261 & ~n57262;
  assign n57264 = n57131 & ~n57263;
  assign n57265 = ~n56304 & n57133;
  assign n57266 = P1_P1_EBX_REG_14_ & ~n57130;
  assign n57267 = ~n57264 & ~n57265;
  assign n9661 = n57266 | ~n57267;
  assign n57269 = P1_P1_EBX_REG_13_ & P1_P1_EBX_REG_14_;
  assign n57270 = n57251 & n57269;
  assign n57271 = P1_P1_EBX_REG_15_ & ~n57270;
  assign n57272 = ~P1_P1_EBX_REG_15_ & n57270;
  assign n57273 = ~n57271 & ~n57272;
  assign n57274 = n57131 & ~n57273;
  assign n57275 = ~n56346 & n57133;
  assign n57276 = P1_P1_EBX_REG_15_ & ~n57130;
  assign n57277 = ~n57274 & ~n57275;
  assign n9666 = n57276 | ~n57277;
  assign n57279 = P1_P1_EBX_REG_15_ & n57270;
  assign n57280 = ~P1_P1_EBX_REG_16_ & n57279;
  assign n57281 = P1_P1_EBX_REG_16_ & ~n57279;
  assign n57282 = ~n57280 & ~n57281;
  assign n57283 = n57131 & ~n57282;
  assign n57284 = ~n56406 & n57133;
  assign n57285 = P1_P1_EBX_REG_16_ & ~n57130;
  assign n57286 = ~n57283 & ~n57284;
  assign n9671 = n57285 | ~n57286;
  assign n57288 = P1_P1_EBX_REG_15_ & P1_P1_EBX_REG_16_;
  assign n57289 = n57270 & n57288;
  assign n57290 = P1_P1_EBX_REG_17_ & ~n57289;
  assign n57291 = ~P1_P1_EBX_REG_17_ & n57289;
  assign n57292 = ~n57290 & ~n57291;
  assign n57293 = n57131 & ~n57292;
  assign n57294 = ~n56452 & n57133;
  assign n57295 = P1_P1_EBX_REG_17_ & ~n57130;
  assign n57296 = ~n57293 & ~n57294;
  assign n9676 = n57295 | ~n57296;
  assign n57298 = P1_P1_EBX_REG_17_ & n57289;
  assign n57299 = ~P1_P1_EBX_REG_18_ & n57298;
  assign n57300 = P1_P1_EBX_REG_18_ & ~n57298;
  assign n57301 = ~n57299 & ~n57300;
  assign n57302 = n57131 & ~n57301;
  assign n57303 = ~n56496 & n57133;
  assign n57304 = P1_P1_EBX_REG_18_ & ~n57130;
  assign n57305 = ~n57302 & ~n57303;
  assign n9681 = n57304 | ~n57305;
  assign n57307 = P1_P1_EBX_REG_19_ & ~n57130;
  assign n57308 = ~n56540 & n57133;
  assign n57309 = P1_P1_EBX_REG_17_ & P1_P1_EBX_REG_18_;
  assign n57310 = n57289 & n57309;
  assign n57311 = P1_P1_EBX_REG_19_ & ~n57310;
  assign n57312 = ~P1_P1_EBX_REG_19_ & n57310;
  assign n57313 = ~n57311 & ~n57312;
  assign n57314 = n57131 & ~n57313;
  assign n57315 = ~n57307 & ~n57308;
  assign n9686 = n57314 | ~n57315;
  assign n57317 = P1_P1_EBX_REG_20_ & ~n57130;
  assign n57318 = ~n56584 & n57133;
  assign n57319 = P1_P1_EBX_REG_19_ & n57310;
  assign n57320 = ~P1_P1_EBX_REG_20_ & n57319;
  assign n57321 = P1_P1_EBX_REG_20_ & ~n57319;
  assign n57322 = ~n57320 & ~n57321;
  assign n57323 = n57131 & ~n57322;
  assign n57324 = ~n57317 & ~n57318;
  assign n9691 = n57323 | ~n57324;
  assign n57326 = P1_P1_EBX_REG_21_ & ~n57130;
  assign n57327 = ~n56628 & n57133;
  assign n57328 = P1_P1_EBX_REG_19_ & P1_P1_EBX_REG_20_;
  assign n57329 = n57310 & n57328;
  assign n57330 = P1_P1_EBX_REG_21_ & ~n57329;
  assign n57331 = ~P1_P1_EBX_REG_21_ & n57329;
  assign n57332 = ~n57330 & ~n57331;
  assign n57333 = n57131 & ~n57332;
  assign n57334 = ~n57326 & ~n57327;
  assign n9696 = n57333 | ~n57334;
  assign n57336 = P1_P1_EBX_REG_22_ & ~n57130;
  assign n57337 = ~n56678 & n57133;
  assign n57338 = P1_P1_EBX_REG_21_ & n57329;
  assign n57339 = ~P1_P1_EBX_REG_22_ & n57338;
  assign n57340 = P1_P1_EBX_REG_22_ & ~n57338;
  assign n57341 = ~n57339 & ~n57340;
  assign n57342 = n57131 & ~n57341;
  assign n57343 = ~n57336 & ~n57337;
  assign n9701 = n57342 | ~n57343;
  assign n57345 = P1_P1_EBX_REG_23_ & ~n57130;
  assign n57346 = ~n56776 & n57133;
  assign n57347 = P1_P1_EBX_REG_21_ & P1_P1_EBX_REG_22_;
  assign n57348 = n57329 & n57347;
  assign n57349 = P1_P1_EBX_REG_23_ & ~n57348;
  assign n57350 = ~P1_P1_EBX_REG_23_ & n57348;
  assign n57351 = ~n57349 & ~n57350;
  assign n57352 = n57131 & ~n57351;
  assign n57353 = ~n57345 & ~n57346;
  assign n9706 = n57352 | ~n57353;
  assign n57355 = P1_P1_EBX_REG_24_ & ~n57130;
  assign n57356 = ~n56824 & n57133;
  assign n57357 = P1_P1_EBX_REG_23_ & n57348;
  assign n57358 = ~P1_P1_EBX_REG_24_ & n57357;
  assign n57359 = P1_P1_EBX_REG_24_ & ~n57357;
  assign n57360 = ~n57358 & ~n57359;
  assign n57361 = n57131 & ~n57360;
  assign n57362 = ~n57355 & ~n57356;
  assign n9711 = n57361 | ~n57362;
  assign n57364 = P1_P1_EBX_REG_25_ & ~n57130;
  assign n57365 = ~n56872 & n57133;
  assign n57366 = P1_P1_EBX_REG_23_ & P1_P1_EBX_REG_24_;
  assign n57367 = n57348 & n57366;
  assign n57368 = P1_P1_EBX_REG_25_ & ~n57367;
  assign n57369 = ~P1_P1_EBX_REG_25_ & n57367;
  assign n57370 = ~n57368 & ~n57369;
  assign n57371 = n57131 & ~n57370;
  assign n57372 = ~n57364 & ~n57365;
  assign n9716 = n57371 | ~n57372;
  assign n57374 = P1_P1_EBX_REG_26_ & ~n57130;
  assign n57375 = ~n56920 & n57133;
  assign n57376 = P1_P1_EBX_REG_25_ & n57367;
  assign n57377 = ~P1_P1_EBX_REG_26_ & n57376;
  assign n57378 = P1_P1_EBX_REG_26_ & ~n57376;
  assign n57379 = ~n57377 & ~n57378;
  assign n57380 = n57131 & ~n57379;
  assign n57381 = ~n57374 & ~n57375;
  assign n9721 = n57380 | ~n57381;
  assign n57383 = P1_P1_EBX_REG_27_ & ~n57130;
  assign n57384 = ~n56968 & n57133;
  assign n57385 = P1_P1_EBX_REG_25_ & P1_P1_EBX_REG_26_;
  assign n57386 = n57367 & n57385;
  assign n57387 = P1_P1_EBX_REG_27_ & ~n57386;
  assign n57388 = ~P1_P1_EBX_REG_27_ & n57386;
  assign n57389 = ~n57387 & ~n57388;
  assign n57390 = n57131 & ~n57389;
  assign n57391 = ~n57383 & ~n57384;
  assign n9726 = n57390 | ~n57391;
  assign n57393 = P1_P1_EBX_REG_28_ & ~n57130;
  assign n57394 = ~n57016 & n57133;
  assign n57395 = P1_P1_EBX_REG_27_ & n57386;
  assign n57396 = ~P1_P1_EBX_REG_28_ & n57395;
  assign n57397 = P1_P1_EBX_REG_28_ & ~n57395;
  assign n57398 = ~n57396 & ~n57397;
  assign n57399 = n57131 & ~n57398;
  assign n57400 = ~n57393 & ~n57394;
  assign n9731 = n57399 | ~n57400;
  assign n57402 = P1_P1_EBX_REG_29_ & ~n57130;
  assign n57403 = ~n57064 & n57133;
  assign n57404 = P1_P1_EBX_REG_27_ & P1_P1_EBX_REG_28_;
  assign n57405 = n57386 & n57404;
  assign n57406 = P1_P1_EBX_REG_29_ & ~n57405;
  assign n57407 = ~P1_P1_EBX_REG_29_ & n57405;
  assign n57408 = ~n57406 & ~n57407;
  assign n57409 = n57131 & ~n57408;
  assign n57410 = ~n57402 & ~n57403;
  assign n9736 = n57409 | ~n57410;
  assign n57412 = P1_P1_EBX_REG_30_ & ~n57130;
  assign n57413 = ~n57112 & n57133;
  assign n57414 = P1_P1_EBX_REG_29_ & n57405;
  assign n57415 = ~P1_P1_EBX_REG_30_ & n57414;
  assign n57416 = P1_P1_EBX_REG_30_ & ~n57414;
  assign n57417 = ~n57415 & ~n57416;
  assign n57418 = n57131 & ~n57417;
  assign n57419 = ~n57412 & ~n57413;
  assign n9741 = n57418 | ~n57419;
  assign n57421 = P1_P1_EBX_REG_31_ & ~n57130;
  assign n57422 = P1_P1_EBX_REG_30_ & n57414;
  assign n57423 = ~P1_P1_EBX_REG_31_ & n57422;
  assign n57424 = P1_P1_EBX_REG_31_ & ~n57422;
  assign n57425 = ~n57423 & ~n57424;
  assign n57426 = n57131 & ~n57425;
  assign n9746 = n57421 | n57426;
  assign n57428 = ~n43990 & ~n44029;
  assign n57429 = ~n51899 & n57428;
  assign n57430 = n43856 & n43864;
  assign n57431 = n43979 & ~n57430;
  assign n57432 = n57429 & ~n57431;
  assign n57433 = P1_P1_STATE2_REG_2_ & ~n57432;
  assign n57434 = n43706 & n57433;
  assign n57435 = ~n43339 & n57434;
  assign n57436 = ~P1_P1_EBX_REG_31_ & n57435;
  assign n57437 = n43624 & n57433;
  assign n57438 = ~n43342 & n57437;
  assign n57439 = n43342 & n57437;
  assign n57440 = ~n43339 & n57439;
  assign n57441 = ~n57436 & ~n57438;
  assign n57442 = ~n57440 & n57441;
  assign n57443 = P1_P1_EBX_REG_0_ & ~n57442;
  assign n57444 = n43339 & n57439;
  assign n57445 = P1_P1_REIP_REG_0_ & n57444;
  assign n57446 = P1_P1_EBX_REG_31_ & n57435;
  assign n57447 = P1_P1_EBX_REG_0_ & n57446;
  assign n57448 = n43701 & n57433;
  assign n57449 = ~P1_P1_INSTQUEUERD_ADDR_REG_0_ & n57448;
  assign n57450 = n43697 & n57433;
  assign n57451 = ~P1_P1_INSTQUEUERD_ADDR_REG_0_ & n57450;
  assign n57452 = ~n57449 & ~n57451;
  assign n57453 = ~n57445 & ~n57447;
  assign n57454 = n57452 & n57453;
  assign n57455 = n43339 & n57434;
  assign n57456 = P1_P1_REIP_REG_0_ & n57455;
  assign n57457 = P1_P1_STATE2_REG_1_ & ~n57432;
  assign n57458 = n55500 & n57457;
  assign n57459 = P1_P1_PHYADDRPOINTER_REG_0_ & n57458;
  assign n57460 = P1_P1_REIP_REG_0_ & n57432;
  assign n57461 = P1_P1_STATE2_REG_3_ & ~n57432;
  assign n57462 = P1_P1_PHYADDRPOINTER_REG_0_ & n57461;
  assign n57463 = ~n57460 & ~n57462;
  assign n57464 = ~n55500 & n57457;
  assign n57465 = P1_P1_PHYADDRPOINTER_REG_0_ & n57464;
  assign n57466 = n57463 & ~n57465;
  assign n57467 = ~n57443 & n57454;
  assign n57468 = ~n57456 & n57467;
  assign n57469 = ~n57459 & n57468;
  assign n9751 = ~n57466 | ~n57469;
  assign n57471 = P1_P1_EBX_REG_1_ & ~n57442;
  assign n57472 = ~P1_P1_REIP_REG_1_ & n57444;
  assign n57473 = ~n57140 & n57446;
  assign n57474 = ~n43348 & ~n43353;
  assign n57475 = n57448 & ~n57474;
  assign n57476 = n57450 & ~n57474;
  assign n57477 = ~n57475 & ~n57476;
  assign n57478 = ~n57472 & ~n57473;
  assign n57479 = n57477 & n57478;
  assign n57480 = ~P1_P1_REIP_REG_1_ & n57455;
  assign n57481 = ~P1_P1_PHYADDRPOINTER_REG_1_ & n57458;
  assign n57482 = P1_P1_REIP_REG_1_ & n57432;
  assign n57483 = P1_P1_PHYADDRPOINTER_REG_1_ & n57461;
  assign n57484 = ~n57482 & ~n57483;
  assign n57485 = P1_P1_PHYADDRPOINTER_REG_0_ & P1_P1_PHYADDRPOINTER_REG_1_;
  assign n57486 = ~P1_P1_PHYADDRPOINTER_REG_0_ & ~P1_P1_PHYADDRPOINTER_REG_1_;
  assign n57487 = ~n57485 & ~n57486;
  assign n57488 = n57464 & ~n57487;
  assign n57489 = n57484 & ~n57488;
  assign n57490 = ~n57471 & n57479;
  assign n57491 = ~n57480 & n57490;
  assign n57492 = ~n57481 & n57491;
  assign n9756 = ~n57489 | ~n57492;
  assign n57494 = P1_P1_EBX_REG_2_ & ~n57442;
  assign n57495 = P1_P1_REIP_REG_1_ & ~P1_P1_REIP_REG_2_;
  assign n57496 = ~P1_P1_REIP_REG_1_ & P1_P1_REIP_REG_2_;
  assign n57497 = ~n57495 & ~n57496;
  assign n57498 = n57444 & ~n57497;
  assign n57499 = ~P1_P1_EBX_REG_0_ & ~P1_P1_EBX_REG_1_;
  assign n57500 = P1_P1_EBX_REG_2_ & ~n57499;
  assign n57501 = ~P1_P1_EBX_REG_2_ & n57499;
  assign n57502 = ~n57500 & ~n57501;
  assign n57503 = n57446 & n57502;
  assign n57504 = ~n43826 & n57448;
  assign n57505 = ~n43826 & n57450;
  assign n57506 = ~n57504 & ~n57505;
  assign n57507 = ~n57498 & ~n57503;
  assign n57508 = n57506 & n57507;
  assign n57509 = n57455 & ~n57497;
  assign n57510 = ~n54836 & n57458;
  assign n57511 = P1_P1_REIP_REG_2_ & n57432;
  assign n57512 = P1_P1_PHYADDRPOINTER_REG_2_ & n57461;
  assign n57513 = ~n57511 & ~n57512;
  assign n57514 = ~P1_P1_PHYADDRPOINTER_REG_0_ & P1_P1_PHYADDRPOINTER_REG_1_;
  assign n57515 = ~n54836 & ~n57514;
  assign n57516 = n54836 & n57514;
  assign n57517 = ~n57515 & ~n57516;
  assign n57518 = n57464 & n57517;
  assign n57519 = n57513 & ~n57518;
  assign n57520 = ~n57494 & n57508;
  assign n57521 = ~n57509 & n57520;
  assign n57522 = ~n57510 & n57521;
  assign n9761 = ~n57519 | ~n57522;
  assign n57524 = P1_P1_EBX_REG_3_ & ~n57442;
  assign n57525 = P1_P1_REIP_REG_1_ & P1_P1_REIP_REG_2_;
  assign n57526 = ~P1_P1_REIP_REG_3_ & n57525;
  assign n57527 = P1_P1_REIP_REG_3_ & ~n57525;
  assign n57528 = ~n57526 & ~n57527;
  assign n57529 = n57444 & ~n57528;
  assign n57530 = ~P1_P1_EBX_REG_3_ & n57501;
  assign n57531 = P1_P1_EBX_REG_3_ & ~n57501;
  assign n57532 = ~n57530 & ~n57531;
  assign n57533 = n57446 & n57532;
  assign n57534 = ~P1_P1_INSTQUEUERD_ADDR_REG_3_ & n43874;
  assign n57535 = ~n43875 & ~n57534;
  assign n57536 = n57448 & ~n57535;
  assign n57537 = n57450 & ~n57535;
  assign n57538 = ~n57536 & ~n57537;
  assign n57539 = ~n57529 & ~n57533;
  assign n57540 = n57538 & n57539;
  assign n57541 = n57455 & ~n57528;
  assign n57542 = ~n54858 & n57458;
  assign n57543 = P1_P1_REIP_REG_3_ & n57432;
  assign n57544 = P1_P1_PHYADDRPOINTER_REG_3_ & n57461;
  assign n57545 = ~n57543 & ~n57544;
  assign n57546 = n54858 & n57516;
  assign n57547 = ~n54858 & ~n57516;
  assign n57548 = ~n57546 & ~n57547;
  assign n57549 = n57464 & n57548;
  assign n57550 = n57545 & ~n57549;
  assign n57551 = ~n57524 & n57540;
  assign n57552 = ~n57541 & n57551;
  assign n57553 = ~n57542 & n57552;
  assign n9766 = ~n57550 | ~n57553;
  assign n57555 = P1_P1_INSTQUEUERD_ADDR_REG_3_ & n43874;
  assign n57556 = ~P1_P1_INSTQUEUERD_ADDR_REG_4_ & n57555;
  assign n57557 = P1_P1_INSTQUEUERD_ADDR_REG_4_ & ~n57555;
  assign n57558 = ~n57556 & ~n57557;
  assign n57559 = n57450 & ~n57558;
  assign n57560 = n57448 & ~n57558;
  assign n57561 = ~n57559 & ~n57560;
  assign n57562 = P1_P1_EBX_REG_4_ & ~n57442;
  assign n57563 = P1_P1_EBX_REG_4_ & ~n57530;
  assign n57564 = ~P1_P1_EBX_REG_3_ & ~P1_P1_EBX_REG_4_;
  assign n57565 = n57501 & n57564;
  assign n57566 = ~n57563 & ~n57565;
  assign n57567 = n57446 & n57566;
  assign n57568 = n51898 & ~n57432;
  assign n57569 = P1_P1_REIP_REG_3_ & n57525;
  assign n57570 = ~P1_P1_REIP_REG_4_ & n57569;
  assign n57571 = P1_P1_REIP_REG_4_ & ~n57569;
  assign n57572 = ~n57570 & ~n57571;
  assign n57573 = n57444 & ~n57572;
  assign n57574 = ~n57567 & ~n57568;
  assign n57575 = ~n57573 & n57574;
  assign n57576 = n57455 & ~n57572;
  assign n57577 = ~n54879 & n57458;
  assign n57578 = n57561 & ~n57562;
  assign n57579 = n57575 & n57578;
  assign n57580 = ~n57576 & n57579;
  assign n57581 = ~n57577 & n57580;
  assign n57582 = P1_P1_REIP_REG_4_ & n57432;
  assign n57583 = P1_P1_PHYADDRPOINTER_REG_4_ & n57461;
  assign n57584 = ~n57582 & ~n57583;
  assign n57585 = ~n54879 & ~n57546;
  assign n57586 = n54858 & n54879;
  assign n57587 = n57516 & n57586;
  assign n57588 = ~n57585 & ~n57587;
  assign n57589 = n57464 & n57588;
  assign n57590 = n57584 & ~n57589;
  assign n9771 = ~n57581 | ~n57590;
  assign n57592 = P1_P1_INSTQUEUERD_ADDR_REG_4_ & n57555;
  assign n57593 = n57450 & n57592;
  assign n57594 = n57448 & n57592;
  assign n57595 = ~n57593 & ~n57594;
  assign n57596 = P1_P1_EBX_REG_5_ & ~n57442;
  assign n57597 = ~P1_P1_EBX_REG_5_ & n57565;
  assign n57598 = P1_P1_EBX_REG_5_ & ~n57565;
  assign n57599 = ~n57597 & ~n57598;
  assign n57600 = n57446 & n57599;
  assign n57601 = P1_P1_REIP_REG_4_ & n57569;
  assign n57602 = ~P1_P1_REIP_REG_5_ & n57601;
  assign n57603 = P1_P1_REIP_REG_5_ & ~n57601;
  assign n57604 = ~n57602 & ~n57603;
  assign n57605 = n57444 & ~n57604;
  assign n57606 = ~n57568 & ~n57600;
  assign n57607 = ~n57605 & n57606;
  assign n57608 = n57455 & ~n57604;
  assign n57609 = ~n54902 & n57458;
  assign n57610 = n57595 & ~n57596;
  assign n57611 = n57607 & n57610;
  assign n57612 = ~n57608 & n57611;
  assign n57613 = ~n57609 & n57612;
  assign n57614 = P1_P1_REIP_REG_5_ & n57432;
  assign n57615 = P1_P1_PHYADDRPOINTER_REG_5_ & n57461;
  assign n57616 = ~n57614 & ~n57615;
  assign n57617 = n54902 & n57587;
  assign n57618 = ~n54902 & ~n57587;
  assign n57619 = ~n57617 & ~n57618;
  assign n57620 = n57464 & n57619;
  assign n57621 = n57616 & ~n57620;
  assign n9776 = ~n57613 | ~n57621;
  assign n57623 = P1_P1_REIP_REG_5_ & n57601;
  assign n57624 = ~P1_P1_REIP_REG_6_ & n57623;
  assign n57625 = P1_P1_REIP_REG_6_ & ~n57623;
  assign n57626 = ~n57624 & ~n57625;
  assign n57627 = n57455 & ~n57626;
  assign n57628 = P1_P1_EBX_REG_6_ & ~n57442;
  assign n57629 = P1_P1_EBX_REG_6_ & ~n57597;
  assign n57630 = ~P1_P1_EBX_REG_5_ & ~P1_P1_EBX_REG_6_;
  assign n57631 = n57565 & n57630;
  assign n57632 = ~n57629 & ~n57631;
  assign n57633 = n57446 & n57632;
  assign n57634 = n57444 & ~n57626;
  assign n57635 = ~n57568 & ~n57633;
  assign n57636 = ~n57634 & n57635;
  assign n57637 = ~n54925 & ~n57617;
  assign n57638 = n54902 & n54925;
  assign n57639 = n57587 & n57638;
  assign n57640 = ~n57637 & ~n57639;
  assign n57641 = n57464 & n57640;
  assign n57642 = P1_P1_REIP_REG_6_ & n57432;
  assign n57643 = P1_P1_PHYADDRPOINTER_REG_6_ & n57461;
  assign n57644 = ~n57642 & ~n57643;
  assign n57645 = ~n54925 & n57458;
  assign n57646 = n57644 & ~n57645;
  assign n57647 = ~n57627 & ~n57628;
  assign n57648 = n57636 & n57647;
  assign n57649 = ~n57641 & n57648;
  assign n9781 = ~n57646 | ~n57649;
  assign n57651 = P1_P1_REIP_REG_6_ & n57623;
  assign n57652 = ~P1_P1_REIP_REG_7_ & n57651;
  assign n57653 = P1_P1_REIP_REG_7_ & ~n57651;
  assign n57654 = ~n57652 & ~n57653;
  assign n57655 = n57455 & ~n57654;
  assign n57656 = P1_P1_EBX_REG_7_ & ~n57442;
  assign n57657 = ~P1_P1_EBX_REG_7_ & n57631;
  assign n57658 = P1_P1_EBX_REG_7_ & ~n57631;
  assign n57659 = ~n57657 & ~n57658;
  assign n57660 = n57446 & n57659;
  assign n57661 = n57444 & ~n57654;
  assign n57662 = ~n57568 & ~n57660;
  assign n57663 = ~n57661 & n57662;
  assign n57664 = n54948 & n57639;
  assign n57665 = ~n54948 & ~n57639;
  assign n57666 = ~n57664 & ~n57665;
  assign n57667 = n57464 & n57666;
  assign n57668 = P1_P1_REIP_REG_7_ & n57432;
  assign n57669 = P1_P1_PHYADDRPOINTER_REG_7_ & n57461;
  assign n57670 = ~n57668 & ~n57669;
  assign n57671 = ~n54948 & n57458;
  assign n57672 = n57670 & ~n57671;
  assign n57673 = ~n57655 & ~n57656;
  assign n57674 = n57663 & n57673;
  assign n57675 = ~n57667 & n57674;
  assign n9786 = ~n57672 | ~n57675;
  assign n57677 = P1_P1_REIP_REG_7_ & n57651;
  assign n57678 = ~P1_P1_REIP_REG_8_ & n57677;
  assign n57679 = P1_P1_REIP_REG_8_ & ~n57677;
  assign n57680 = ~n57678 & ~n57679;
  assign n57681 = n57455 & ~n57680;
  assign n57682 = P1_P1_EBX_REG_8_ & ~n57442;
  assign n57683 = P1_P1_EBX_REG_8_ & ~n57657;
  assign n57684 = ~P1_P1_EBX_REG_7_ & ~P1_P1_EBX_REG_8_;
  assign n57685 = n57631 & n57684;
  assign n57686 = ~n57683 & ~n57685;
  assign n57687 = n57446 & n57686;
  assign n57688 = n57444 & ~n57680;
  assign n57689 = ~n57568 & ~n57687;
  assign n57690 = ~n57688 & n57689;
  assign n57691 = ~n54971 & ~n57664;
  assign n57692 = n54948 & n54971;
  assign n57693 = n57639 & n57692;
  assign n57694 = ~n57691 & ~n57693;
  assign n57695 = n57464 & n57694;
  assign n57696 = P1_P1_REIP_REG_8_ & n57432;
  assign n57697 = P1_P1_PHYADDRPOINTER_REG_8_ & n57461;
  assign n57698 = ~n57696 & ~n57697;
  assign n57699 = ~n54971 & n57458;
  assign n57700 = n57698 & ~n57699;
  assign n57701 = ~n57681 & ~n57682;
  assign n57702 = n57690 & n57701;
  assign n57703 = ~n57695 & n57702;
  assign n9791 = ~n57700 | ~n57703;
  assign n57705 = P1_P1_REIP_REG_8_ & n57677;
  assign n57706 = ~P1_P1_REIP_REG_9_ & n57705;
  assign n57707 = P1_P1_REIP_REG_9_ & ~n57705;
  assign n57708 = ~n57706 & ~n57707;
  assign n57709 = n57455 & ~n57708;
  assign n57710 = P1_P1_EBX_REG_9_ & ~n57442;
  assign n57711 = ~P1_P1_EBX_REG_9_ & n57685;
  assign n57712 = P1_P1_EBX_REG_9_ & ~n57685;
  assign n57713 = ~n57711 & ~n57712;
  assign n57714 = n57446 & n57713;
  assign n57715 = n57444 & ~n57708;
  assign n57716 = ~n57568 & ~n57714;
  assign n57717 = ~n57715 & n57716;
  assign n57718 = n54994 & n57693;
  assign n57719 = ~n54994 & ~n57693;
  assign n57720 = ~n57718 & ~n57719;
  assign n57721 = n57464 & n57720;
  assign n57722 = P1_P1_REIP_REG_9_ & n57432;
  assign n57723 = P1_P1_PHYADDRPOINTER_REG_9_ & n57461;
  assign n57724 = ~n57722 & ~n57723;
  assign n57725 = ~n54994 & n57458;
  assign n57726 = n57724 & ~n57725;
  assign n57727 = ~n57709 & ~n57710;
  assign n57728 = n57717 & n57727;
  assign n57729 = ~n57721 & n57728;
  assign n9796 = ~n57726 | ~n57729;
  assign n57731 = P1_P1_REIP_REG_9_ & n57705;
  assign n57732 = ~P1_P1_REIP_REG_10_ & n57731;
  assign n57733 = P1_P1_REIP_REG_10_ & ~n57731;
  assign n57734 = ~n57732 & ~n57733;
  assign n57735 = n57455 & ~n57734;
  assign n57736 = P1_P1_EBX_REG_10_ & ~n57442;
  assign n57737 = P1_P1_EBX_REG_10_ & ~n57711;
  assign n57738 = ~P1_P1_EBX_REG_9_ & ~P1_P1_EBX_REG_10_;
  assign n57739 = n57685 & n57738;
  assign n57740 = ~n57737 & ~n57739;
  assign n57741 = n57446 & n57740;
  assign n57742 = n57444 & ~n57734;
  assign n57743 = ~n57568 & ~n57741;
  assign n57744 = ~n57742 & n57743;
  assign n57745 = ~n55017 & ~n57718;
  assign n57746 = n54994 & n55017;
  assign n57747 = n57693 & n57746;
  assign n57748 = ~n57745 & ~n57747;
  assign n57749 = n57464 & n57748;
  assign n57750 = P1_P1_REIP_REG_10_ & n57432;
  assign n57751 = P1_P1_PHYADDRPOINTER_REG_10_ & n57461;
  assign n57752 = ~n57750 & ~n57751;
  assign n57753 = ~n55017 & n57458;
  assign n57754 = n57752 & ~n57753;
  assign n57755 = ~n57735 & ~n57736;
  assign n57756 = n57744 & n57755;
  assign n57757 = ~n57749 & n57756;
  assign n9801 = ~n57754 | ~n57757;
  assign n57759 = P1_P1_REIP_REG_10_ & n57731;
  assign n57760 = ~P1_P1_REIP_REG_11_ & n57759;
  assign n57761 = P1_P1_REIP_REG_11_ & ~n57759;
  assign n57762 = ~n57760 & ~n57761;
  assign n57763 = n57455 & ~n57762;
  assign n57764 = P1_P1_EBX_REG_11_ & ~n57442;
  assign n57765 = ~P1_P1_EBX_REG_11_ & n57739;
  assign n57766 = P1_P1_EBX_REG_11_ & ~n57739;
  assign n57767 = ~n57765 & ~n57766;
  assign n57768 = n57446 & n57767;
  assign n57769 = n57444 & ~n57762;
  assign n57770 = ~n57568 & ~n57768;
  assign n57771 = ~n57769 & n57770;
  assign n57772 = n55040 & n57747;
  assign n57773 = ~n55040 & ~n57747;
  assign n57774 = ~n57772 & ~n57773;
  assign n57775 = n57464 & n57774;
  assign n57776 = P1_P1_REIP_REG_11_ & n57432;
  assign n57777 = P1_P1_PHYADDRPOINTER_REG_11_ & n57461;
  assign n57778 = ~n57776 & ~n57777;
  assign n57779 = ~n55040 & n57458;
  assign n57780 = n57778 & ~n57779;
  assign n57781 = ~n57763 & ~n57764;
  assign n57782 = n57771 & n57781;
  assign n57783 = ~n57775 & n57782;
  assign n9806 = ~n57780 | ~n57783;
  assign n57785 = P1_P1_REIP_REG_11_ & n57759;
  assign n57786 = ~P1_P1_REIP_REG_12_ & n57785;
  assign n57787 = P1_P1_REIP_REG_12_ & ~n57785;
  assign n57788 = ~n57786 & ~n57787;
  assign n57789 = n57455 & ~n57788;
  assign n57790 = P1_P1_EBX_REG_12_ & ~n57442;
  assign n57791 = P1_P1_EBX_REG_12_ & ~n57765;
  assign n57792 = ~P1_P1_EBX_REG_11_ & ~P1_P1_EBX_REG_12_;
  assign n57793 = n57739 & n57792;
  assign n57794 = ~n57791 & ~n57793;
  assign n57795 = n57446 & n57794;
  assign n57796 = n57444 & ~n57788;
  assign n57797 = ~n57568 & ~n57795;
  assign n57798 = ~n57796 & n57797;
  assign n57799 = ~n55063 & ~n57772;
  assign n57800 = n55040 & n55063;
  assign n57801 = n57747 & n57800;
  assign n57802 = ~n57799 & ~n57801;
  assign n57803 = n57464 & n57802;
  assign n57804 = P1_P1_REIP_REG_12_ & n57432;
  assign n57805 = P1_P1_PHYADDRPOINTER_REG_12_ & n57461;
  assign n57806 = ~n57804 & ~n57805;
  assign n57807 = ~n55063 & n57458;
  assign n57808 = n57806 & ~n57807;
  assign n57809 = ~n57789 & ~n57790;
  assign n57810 = n57798 & n57809;
  assign n57811 = ~n57803 & n57810;
  assign n9811 = ~n57808 | ~n57811;
  assign n57813 = P1_P1_REIP_REG_12_ & n57785;
  assign n57814 = ~P1_P1_REIP_REG_13_ & n57813;
  assign n57815 = P1_P1_REIP_REG_13_ & ~n57813;
  assign n57816 = ~n57814 & ~n57815;
  assign n57817 = n57455 & ~n57816;
  assign n57818 = P1_P1_EBX_REG_13_ & ~n57442;
  assign n57819 = ~P1_P1_EBX_REG_13_ & n57793;
  assign n57820 = P1_P1_EBX_REG_13_ & ~n57793;
  assign n57821 = ~n57819 & ~n57820;
  assign n57822 = n57446 & n57821;
  assign n57823 = n57444 & ~n57816;
  assign n57824 = ~n57568 & ~n57822;
  assign n57825 = ~n57823 & n57824;
  assign n57826 = n55086 & n57801;
  assign n57827 = ~n55086 & ~n57801;
  assign n57828 = ~n57826 & ~n57827;
  assign n57829 = n57464 & n57828;
  assign n57830 = P1_P1_REIP_REG_13_ & n57432;
  assign n57831 = P1_P1_PHYADDRPOINTER_REG_13_ & n57461;
  assign n57832 = ~n57830 & ~n57831;
  assign n57833 = ~n55086 & n57458;
  assign n57834 = n57832 & ~n57833;
  assign n57835 = ~n57817 & ~n57818;
  assign n57836 = n57825 & n57835;
  assign n57837 = ~n57829 & n57836;
  assign n9816 = ~n57834 | ~n57837;
  assign n57839 = P1_P1_REIP_REG_13_ & n57813;
  assign n57840 = ~P1_P1_REIP_REG_14_ & n57839;
  assign n57841 = P1_P1_REIP_REG_14_ & ~n57839;
  assign n57842 = ~n57840 & ~n57841;
  assign n57843 = n57455 & ~n57842;
  assign n57844 = P1_P1_EBX_REG_14_ & ~n57442;
  assign n57845 = P1_P1_EBX_REG_14_ & ~n57819;
  assign n57846 = ~P1_P1_EBX_REG_13_ & ~P1_P1_EBX_REG_14_;
  assign n57847 = n57793 & n57846;
  assign n57848 = ~n57845 & ~n57847;
  assign n57849 = n57446 & n57848;
  assign n57850 = n57444 & ~n57842;
  assign n57851 = ~n57568 & ~n57849;
  assign n57852 = ~n57850 & n57851;
  assign n57853 = ~n55109 & ~n57826;
  assign n57854 = n55086 & n55109;
  assign n57855 = n57801 & n57854;
  assign n57856 = ~n57853 & ~n57855;
  assign n57857 = n57464 & n57856;
  assign n57858 = P1_P1_REIP_REG_14_ & n57432;
  assign n57859 = P1_P1_PHYADDRPOINTER_REG_14_ & n57461;
  assign n57860 = ~n57858 & ~n57859;
  assign n57861 = ~n55109 & n57458;
  assign n57862 = n57860 & ~n57861;
  assign n57863 = ~n57843 & ~n57844;
  assign n57864 = n57852 & n57863;
  assign n57865 = ~n57857 & n57864;
  assign n9821 = ~n57862 | ~n57865;
  assign n57867 = P1_P1_REIP_REG_14_ & n57839;
  assign n57868 = ~P1_P1_REIP_REG_15_ & n57867;
  assign n57869 = P1_P1_REIP_REG_15_ & ~n57867;
  assign n57870 = ~n57868 & ~n57869;
  assign n57871 = n57455 & ~n57870;
  assign n57872 = P1_P1_EBX_REG_15_ & ~n57442;
  assign n57873 = ~P1_P1_EBX_REG_15_ & n57847;
  assign n57874 = P1_P1_EBX_REG_15_ & ~n57847;
  assign n57875 = ~n57873 & ~n57874;
  assign n57876 = n57446 & n57875;
  assign n57877 = n57444 & ~n57870;
  assign n57878 = ~n57568 & ~n57876;
  assign n57879 = ~n57877 & n57878;
  assign n57880 = n55132 & n57855;
  assign n57881 = ~n55132 & ~n57855;
  assign n57882 = ~n57880 & ~n57881;
  assign n57883 = n57464 & n57882;
  assign n57884 = P1_P1_REIP_REG_15_ & n57432;
  assign n57885 = P1_P1_PHYADDRPOINTER_REG_15_ & n57461;
  assign n57886 = ~n57884 & ~n57885;
  assign n57887 = ~n55132 & n57458;
  assign n57888 = n57886 & ~n57887;
  assign n57889 = ~n57871 & ~n57872;
  assign n57890 = n57879 & n57889;
  assign n57891 = ~n57883 & n57890;
  assign n9826 = ~n57888 | ~n57891;
  assign n57893 = P1_P1_REIP_REG_15_ & n57867;
  assign n57894 = ~P1_P1_REIP_REG_16_ & n57893;
  assign n57895 = P1_P1_REIP_REG_16_ & ~n57893;
  assign n57896 = ~n57894 & ~n57895;
  assign n57897 = n57455 & ~n57896;
  assign n57898 = P1_P1_EBX_REG_16_ & ~n57442;
  assign n57899 = P1_P1_EBX_REG_16_ & ~n57873;
  assign n57900 = ~P1_P1_EBX_REG_15_ & ~P1_P1_EBX_REG_16_;
  assign n57901 = n57847 & n57900;
  assign n57902 = ~n57899 & ~n57901;
  assign n57903 = n57446 & n57902;
  assign n57904 = n57444 & ~n57896;
  assign n57905 = ~n57568 & ~n57903;
  assign n57906 = ~n57904 & n57905;
  assign n57907 = ~n55155 & ~n57880;
  assign n57908 = n55132 & n55155;
  assign n57909 = n57855 & n57908;
  assign n57910 = ~n57907 & ~n57909;
  assign n57911 = n57464 & n57910;
  assign n57912 = P1_P1_REIP_REG_16_ & n57432;
  assign n57913 = P1_P1_PHYADDRPOINTER_REG_16_ & n57461;
  assign n57914 = ~n57912 & ~n57913;
  assign n57915 = ~n55155 & n57458;
  assign n57916 = n57914 & ~n57915;
  assign n57917 = ~n57897 & ~n57898;
  assign n57918 = n57906 & n57917;
  assign n57919 = ~n57911 & n57918;
  assign n9831 = ~n57916 | ~n57919;
  assign n57921 = P1_P1_REIP_REG_16_ & n57893;
  assign n57922 = ~P1_P1_REIP_REG_17_ & n57921;
  assign n57923 = P1_P1_REIP_REG_17_ & ~n57921;
  assign n57924 = ~n57922 & ~n57923;
  assign n57925 = n57455 & ~n57924;
  assign n57926 = P1_P1_EBX_REG_17_ & ~n57442;
  assign n57927 = ~P1_P1_EBX_REG_17_ & n57901;
  assign n57928 = P1_P1_EBX_REG_17_ & ~n57901;
  assign n57929 = ~n57927 & ~n57928;
  assign n57930 = n57446 & n57929;
  assign n57931 = n57444 & ~n57924;
  assign n57932 = ~n57568 & ~n57930;
  assign n57933 = ~n57931 & n57932;
  assign n57934 = n55178 & n57909;
  assign n57935 = ~n55178 & ~n57909;
  assign n57936 = ~n57934 & ~n57935;
  assign n57937 = n57464 & n57936;
  assign n57938 = P1_P1_REIP_REG_17_ & n57432;
  assign n57939 = P1_P1_PHYADDRPOINTER_REG_17_ & n57461;
  assign n57940 = ~n57938 & ~n57939;
  assign n57941 = ~n55178 & n57458;
  assign n57942 = n57940 & ~n57941;
  assign n57943 = ~n57925 & ~n57926;
  assign n57944 = n57933 & n57943;
  assign n57945 = ~n57937 & n57944;
  assign n9836 = ~n57942 | ~n57945;
  assign n57947 = P1_P1_REIP_REG_17_ & n57921;
  assign n57948 = ~P1_P1_REIP_REG_18_ & n57947;
  assign n57949 = P1_P1_REIP_REG_18_ & ~n57947;
  assign n57950 = ~n57948 & ~n57949;
  assign n57951 = n57455 & ~n57950;
  assign n57952 = P1_P1_EBX_REG_18_ & ~n57442;
  assign n57953 = P1_P1_EBX_REG_18_ & ~n57927;
  assign n57954 = ~P1_P1_EBX_REG_17_ & ~P1_P1_EBX_REG_18_;
  assign n57955 = n57901 & n57954;
  assign n57956 = ~n57953 & ~n57955;
  assign n57957 = n57446 & n57956;
  assign n57958 = n57444 & ~n57950;
  assign n57959 = ~n57568 & ~n57957;
  assign n57960 = ~n57958 & n57959;
  assign n57961 = ~n55201 & ~n57934;
  assign n57962 = n55178 & n55201;
  assign n57963 = n57909 & n57962;
  assign n57964 = ~n57961 & ~n57963;
  assign n57965 = n57464 & n57964;
  assign n57966 = P1_P1_REIP_REG_18_ & n57432;
  assign n57967 = P1_P1_PHYADDRPOINTER_REG_18_ & n57461;
  assign n57968 = ~n57966 & ~n57967;
  assign n57969 = ~n55201 & n57458;
  assign n57970 = n57968 & ~n57969;
  assign n57971 = ~n57951 & ~n57952;
  assign n57972 = n57960 & n57971;
  assign n57973 = ~n57965 & n57972;
  assign n9841 = ~n57970 | ~n57973;
  assign n57975 = P1_P1_REIP_REG_18_ & n57947;
  assign n57976 = ~P1_P1_REIP_REG_19_ & n57975;
  assign n57977 = P1_P1_REIP_REG_19_ & ~n57975;
  assign n57978 = ~n57976 & ~n57977;
  assign n57979 = n57455 & ~n57978;
  assign n57980 = P1_P1_EBX_REG_19_ & ~n57442;
  assign n57981 = ~P1_P1_EBX_REG_19_ & n57955;
  assign n57982 = P1_P1_EBX_REG_19_ & ~n57955;
  assign n57983 = ~n57981 & ~n57982;
  assign n57984 = n57446 & n57983;
  assign n57985 = n57444 & ~n57978;
  assign n57986 = ~n57568 & ~n57984;
  assign n57987 = ~n57985 & n57986;
  assign n57988 = n55224 & n57963;
  assign n57989 = ~n55224 & ~n57963;
  assign n57990 = ~n57988 & ~n57989;
  assign n57991 = n57464 & n57990;
  assign n57992 = P1_P1_REIP_REG_19_ & n57432;
  assign n57993 = P1_P1_PHYADDRPOINTER_REG_19_ & n57461;
  assign n57994 = ~n57992 & ~n57993;
  assign n57995 = ~n55224 & n57458;
  assign n57996 = n57994 & ~n57995;
  assign n57997 = ~n57979 & ~n57980;
  assign n57998 = n57987 & n57997;
  assign n57999 = ~n57991 & n57998;
  assign n9846 = ~n57996 | ~n57999;
  assign n58001 = P1_P1_REIP_REG_19_ & n57975;
  assign n58002 = ~P1_P1_REIP_REG_20_ & n58001;
  assign n58003 = P1_P1_REIP_REG_20_ & ~n58001;
  assign n58004 = ~n58002 & ~n58003;
  assign n58005 = n57444 & ~n58004;
  assign n58006 = P1_P1_EBX_REG_20_ & ~n57981;
  assign n58007 = ~P1_P1_EBX_REG_19_ & ~P1_P1_EBX_REG_20_;
  assign n58008 = n57955 & n58007;
  assign n58009 = ~n58006 & ~n58008;
  assign n58010 = n57446 & n58009;
  assign n58011 = n57455 & ~n58004;
  assign n58012 = ~n58005 & ~n58010;
  assign n58013 = ~n58011 & n58012;
  assign n58014 = P1_P1_EBX_REG_20_ & ~n57442;
  assign n58015 = ~n55247 & ~n57988;
  assign n58016 = n55224 & n55247;
  assign n58017 = n57963 & n58016;
  assign n58018 = ~n58015 & ~n58017;
  assign n58019 = n57464 & n58018;
  assign n58020 = P1_P1_REIP_REG_20_ & n57432;
  assign n58021 = P1_P1_PHYADDRPOINTER_REG_20_ & n57461;
  assign n58022 = ~n58020 & ~n58021;
  assign n58023 = ~n55247 & n57458;
  assign n58024 = n58022 & ~n58023;
  assign n58025 = n58013 & ~n58014;
  assign n58026 = ~n58019 & n58025;
  assign n9851 = ~n58024 | ~n58026;
  assign n58028 = P1_P1_REIP_REG_20_ & n58001;
  assign n58029 = ~P1_P1_REIP_REG_21_ & n58028;
  assign n58030 = P1_P1_REIP_REG_21_ & ~n58028;
  assign n58031 = ~n58029 & ~n58030;
  assign n58032 = n57444 & ~n58031;
  assign n58033 = ~P1_P1_EBX_REG_21_ & n58008;
  assign n58034 = P1_P1_EBX_REG_21_ & ~n58008;
  assign n58035 = ~n58033 & ~n58034;
  assign n58036 = n57446 & n58035;
  assign n58037 = n57455 & ~n58031;
  assign n58038 = ~n58032 & ~n58036;
  assign n58039 = ~n58037 & n58038;
  assign n58040 = P1_P1_EBX_REG_21_ & ~n57442;
  assign n58041 = n55270 & n58017;
  assign n58042 = ~n55270 & ~n58017;
  assign n58043 = ~n58041 & ~n58042;
  assign n58044 = n57464 & n58043;
  assign n58045 = P1_P1_REIP_REG_21_ & n57432;
  assign n58046 = P1_P1_PHYADDRPOINTER_REG_21_ & n57461;
  assign n58047 = ~n58045 & ~n58046;
  assign n58048 = ~n55270 & n57458;
  assign n58049 = n58047 & ~n58048;
  assign n58050 = n58039 & ~n58040;
  assign n58051 = ~n58044 & n58050;
  assign n9856 = ~n58049 | ~n58051;
  assign n58053 = P1_P1_REIP_REG_21_ & n58028;
  assign n58054 = ~P1_P1_REIP_REG_22_ & n58053;
  assign n58055 = P1_P1_REIP_REG_22_ & ~n58053;
  assign n58056 = ~n58054 & ~n58055;
  assign n58057 = n57444 & ~n58056;
  assign n58058 = P1_P1_EBX_REG_22_ & ~n58033;
  assign n58059 = ~P1_P1_EBX_REG_21_ & ~P1_P1_EBX_REG_22_;
  assign n58060 = n58008 & n58059;
  assign n58061 = ~n58058 & ~n58060;
  assign n58062 = n57446 & n58061;
  assign n58063 = n57455 & ~n58056;
  assign n58064 = ~n58057 & ~n58062;
  assign n58065 = ~n58063 & n58064;
  assign n58066 = P1_P1_EBX_REG_22_ & ~n57442;
  assign n58067 = ~n55293 & ~n58041;
  assign n58068 = n55270 & n55293;
  assign n58069 = n58017 & n58068;
  assign n58070 = ~n58067 & ~n58069;
  assign n58071 = n57464 & n58070;
  assign n58072 = P1_P1_REIP_REG_22_ & n57432;
  assign n58073 = P1_P1_PHYADDRPOINTER_REG_22_ & n57461;
  assign n58074 = ~n58072 & ~n58073;
  assign n58075 = ~n55293 & n57458;
  assign n58076 = n58074 & ~n58075;
  assign n58077 = n58065 & ~n58066;
  assign n58078 = ~n58071 & n58077;
  assign n9861 = ~n58076 | ~n58078;
  assign n58080 = P1_P1_REIP_REG_22_ & n58053;
  assign n58081 = ~P1_P1_REIP_REG_23_ & n58080;
  assign n58082 = P1_P1_REIP_REG_23_ & ~n58080;
  assign n58083 = ~n58081 & ~n58082;
  assign n58084 = n57444 & ~n58083;
  assign n58085 = ~P1_P1_EBX_REG_23_ & n58060;
  assign n58086 = P1_P1_EBX_REG_23_ & ~n58060;
  assign n58087 = ~n58085 & ~n58086;
  assign n58088 = n57446 & n58087;
  assign n58089 = n57455 & ~n58083;
  assign n58090 = ~n58084 & ~n58088;
  assign n58091 = ~n58089 & n58090;
  assign n58092 = P1_P1_EBX_REG_23_ & ~n57442;
  assign n58093 = n55316 & n58069;
  assign n58094 = ~n55316 & ~n58069;
  assign n58095 = ~n58093 & ~n58094;
  assign n58096 = n57464 & n58095;
  assign n58097 = P1_P1_REIP_REG_23_ & n57432;
  assign n58098 = P1_P1_PHYADDRPOINTER_REG_23_ & n57461;
  assign n58099 = ~n58097 & ~n58098;
  assign n58100 = ~n55316 & n57458;
  assign n58101 = n58099 & ~n58100;
  assign n58102 = n58091 & ~n58092;
  assign n58103 = ~n58096 & n58102;
  assign n9866 = ~n58101 | ~n58103;
  assign n58105 = P1_P1_REIP_REG_23_ & n58080;
  assign n58106 = ~P1_P1_REIP_REG_24_ & n58105;
  assign n58107 = P1_P1_REIP_REG_24_ & ~n58105;
  assign n58108 = ~n58106 & ~n58107;
  assign n58109 = n57455 & ~n58108;
  assign n58110 = P1_P1_EBX_REG_24_ & ~n57442;
  assign n58111 = n57444 & ~n58108;
  assign n58112 = P1_P1_EBX_REG_24_ & ~n58085;
  assign n58113 = ~P1_P1_EBX_REG_23_ & ~P1_P1_EBX_REG_24_;
  assign n58114 = n58060 & n58113;
  assign n58115 = ~n58112 & ~n58114;
  assign n58116 = n57446 & n58115;
  assign n58117 = ~n58111 & ~n58116;
  assign n58118 = ~n55339 & ~n58093;
  assign n58119 = n55316 & n55339;
  assign n58120 = n58069 & n58119;
  assign n58121 = ~n58118 & ~n58120;
  assign n58122 = n57464 & n58121;
  assign n58123 = P1_P1_REIP_REG_24_ & n57432;
  assign n58124 = P1_P1_PHYADDRPOINTER_REG_24_ & n57461;
  assign n58125 = ~n58123 & ~n58124;
  assign n58126 = ~n55339 & n57458;
  assign n58127 = n58125 & ~n58126;
  assign n58128 = ~n58109 & ~n58110;
  assign n58129 = n58117 & n58128;
  assign n58130 = ~n58122 & n58129;
  assign n9871 = ~n58127 | ~n58130;
  assign n58132 = P1_P1_REIP_REG_24_ & n58105;
  assign n58133 = ~P1_P1_REIP_REG_25_ & n58132;
  assign n58134 = P1_P1_REIP_REG_25_ & ~n58132;
  assign n58135 = ~n58133 & ~n58134;
  assign n58136 = n57455 & ~n58135;
  assign n58137 = P1_P1_EBX_REG_25_ & ~n57442;
  assign n58138 = n57444 & ~n58135;
  assign n58139 = ~P1_P1_EBX_REG_25_ & n58114;
  assign n58140 = P1_P1_EBX_REG_25_ & ~n58114;
  assign n58141 = ~n58139 & ~n58140;
  assign n58142 = n57446 & n58141;
  assign n58143 = ~n58138 & ~n58142;
  assign n58144 = n55362 & n58120;
  assign n58145 = ~n55362 & ~n58120;
  assign n58146 = ~n58144 & ~n58145;
  assign n58147 = n57464 & n58146;
  assign n58148 = P1_P1_REIP_REG_25_ & n57432;
  assign n58149 = P1_P1_PHYADDRPOINTER_REG_25_ & n57461;
  assign n58150 = ~n58148 & ~n58149;
  assign n58151 = ~n55362 & n57458;
  assign n58152 = n58150 & ~n58151;
  assign n58153 = ~n58136 & ~n58137;
  assign n58154 = n58143 & n58153;
  assign n58155 = ~n58147 & n58154;
  assign n9876 = ~n58152 | ~n58155;
  assign n58157 = P1_P1_REIP_REG_25_ & n58132;
  assign n58158 = ~P1_P1_REIP_REG_26_ & n58157;
  assign n58159 = P1_P1_REIP_REG_26_ & ~n58157;
  assign n58160 = ~n58158 & ~n58159;
  assign n58161 = n57455 & ~n58160;
  assign n58162 = P1_P1_EBX_REG_26_ & ~n57442;
  assign n58163 = n57444 & ~n58160;
  assign n58164 = P1_P1_EBX_REG_26_ & ~n58139;
  assign n58165 = ~P1_P1_EBX_REG_25_ & ~P1_P1_EBX_REG_26_;
  assign n58166 = n58114 & n58165;
  assign n58167 = ~n58164 & ~n58166;
  assign n58168 = n57446 & n58167;
  assign n58169 = ~n58163 & ~n58168;
  assign n58170 = ~n55385 & ~n58144;
  assign n58171 = n55362 & n55385;
  assign n58172 = n58120 & n58171;
  assign n58173 = ~n58170 & ~n58172;
  assign n58174 = n57464 & n58173;
  assign n58175 = P1_P1_REIP_REG_26_ & n57432;
  assign n58176 = P1_P1_PHYADDRPOINTER_REG_26_ & n57461;
  assign n58177 = ~n58175 & ~n58176;
  assign n58178 = ~n55385 & n57458;
  assign n58179 = n58177 & ~n58178;
  assign n58180 = ~n58161 & ~n58162;
  assign n58181 = n58169 & n58180;
  assign n58182 = ~n58174 & n58181;
  assign n9881 = ~n58179 | ~n58182;
  assign n58184 = P1_P1_REIP_REG_26_ & n58157;
  assign n58185 = ~P1_P1_REIP_REG_27_ & n58184;
  assign n58186 = P1_P1_REIP_REG_27_ & ~n58184;
  assign n58187 = ~n58185 & ~n58186;
  assign n58188 = n57455 & ~n58187;
  assign n58189 = P1_P1_EBX_REG_27_ & ~n57442;
  assign n58190 = n57444 & ~n58187;
  assign n58191 = ~P1_P1_EBX_REG_27_ & n58166;
  assign n58192 = P1_P1_EBX_REG_27_ & ~n58166;
  assign n58193 = ~n58191 & ~n58192;
  assign n58194 = n57446 & n58193;
  assign n58195 = ~n58190 & ~n58194;
  assign n58196 = n55408 & n58172;
  assign n58197 = ~n55408 & ~n58172;
  assign n58198 = ~n58196 & ~n58197;
  assign n58199 = n57464 & n58198;
  assign n58200 = P1_P1_REIP_REG_27_ & n57432;
  assign n58201 = P1_P1_PHYADDRPOINTER_REG_27_ & n57461;
  assign n58202 = ~n58200 & ~n58201;
  assign n58203 = ~n55408 & n57458;
  assign n58204 = n58202 & ~n58203;
  assign n58205 = ~n58188 & ~n58189;
  assign n58206 = n58195 & n58205;
  assign n58207 = ~n58199 & n58206;
  assign n9886 = ~n58204 | ~n58207;
  assign n58209 = P1_P1_REIP_REG_27_ & n58184;
  assign n58210 = ~P1_P1_REIP_REG_28_ & n58209;
  assign n58211 = P1_P1_REIP_REG_28_ & ~n58209;
  assign n58212 = ~n58210 & ~n58211;
  assign n58213 = n57455 & ~n58212;
  assign n58214 = P1_P1_EBX_REG_28_ & ~n57442;
  assign n58215 = n57444 & ~n58212;
  assign n58216 = P1_P1_EBX_REG_28_ & ~n58191;
  assign n58217 = ~P1_P1_EBX_REG_27_ & ~P1_P1_EBX_REG_28_;
  assign n58218 = n58166 & n58217;
  assign n58219 = ~n58216 & ~n58218;
  assign n58220 = n57446 & n58219;
  assign n58221 = ~n55431 & ~n58196;
  assign n58222 = n55408 & n55431;
  assign n58223 = n58172 & n58222;
  assign n58224 = ~n58221 & ~n58223;
  assign n58225 = n57464 & n58224;
  assign n58226 = ~n58213 & ~n58214;
  assign n58227 = ~n58215 & n58226;
  assign n58228 = ~n58220 & n58227;
  assign n58229 = ~n58225 & n58228;
  assign n58230 = P1_P1_REIP_REG_28_ & n57432;
  assign n58231 = P1_P1_PHYADDRPOINTER_REG_28_ & n57461;
  assign n58232 = ~n58230 & ~n58231;
  assign n58233 = ~n55431 & n57458;
  assign n58234 = n58232 & ~n58233;
  assign n9891 = ~n58229 | ~n58234;
  assign n58236 = P1_P1_REIP_REG_28_ & n58209;
  assign n58237 = ~P1_P1_REIP_REG_29_ & n58236;
  assign n58238 = P1_P1_REIP_REG_29_ & ~n58236;
  assign n58239 = ~n58237 & ~n58238;
  assign n58240 = n57455 & ~n58239;
  assign n58241 = P1_P1_EBX_REG_29_ & ~n57442;
  assign n58242 = n57444 & ~n58239;
  assign n58243 = P1_P1_EBX_REG_29_ & ~n58218;
  assign n58244 = ~P1_P1_EBX_REG_29_ & n58218;
  assign n58245 = ~n58243 & ~n58244;
  assign n58246 = n57446 & n58245;
  assign n58247 = ~n58242 & ~n58246;
  assign n58248 = ~n55454 & ~n58223;
  assign n58249 = n55454 & n58223;
  assign n58250 = ~n58248 & ~n58249;
  assign n58251 = n57464 & n58250;
  assign n58252 = P1_P1_REIP_REG_29_ & n57432;
  assign n58253 = P1_P1_PHYADDRPOINTER_REG_29_ & n57461;
  assign n58254 = ~n58252 & ~n58253;
  assign n58255 = ~n55454 & n57458;
  assign n58256 = n58254 & ~n58255;
  assign n58257 = ~n58240 & ~n58241;
  assign n58258 = n58247 & n58257;
  assign n58259 = ~n58251 & n58258;
  assign n9896 = ~n58256 | ~n58259;
  assign n58261 = P1_P1_REIP_REG_29_ & n58236;
  assign n58262 = ~P1_P1_REIP_REG_30_ & n58261;
  assign n58263 = P1_P1_REIP_REG_30_ & ~n58261;
  assign n58264 = ~n58262 & ~n58263;
  assign n58265 = n57455 & ~n58264;
  assign n58266 = P1_P1_EBX_REG_30_ & ~n57442;
  assign n58267 = n57444 & ~n58264;
  assign n58268 = ~P1_P1_EBX_REG_30_ & n58244;
  assign n58269 = P1_P1_EBX_REG_30_ & ~n58244;
  assign n58270 = ~n58268 & ~n58269;
  assign n58271 = n57446 & n58270;
  assign n58272 = P1_P1_REIP_REG_30_ & n57432;
  assign n58273 = P1_P1_PHYADDRPOINTER_REG_30_ & n57461;
  assign n58274 = ~n58272 & ~n58273;
  assign n58275 = ~n55477 & n57458;
  assign n58276 = n58274 & ~n58275;
  assign n58277 = ~n58265 & ~n58266;
  assign n58278 = ~n58267 & n58277;
  assign n58279 = ~n58271 & n58278;
  assign n58280 = n58276 & n58279;
  assign n58281 = n55477 & n58249;
  assign n58282 = ~n55477 & ~n58249;
  assign n58283 = ~n58281 & ~n58282;
  assign n58284 = n57464 & n58283;
  assign n9901 = ~n58280 | n58284;
  assign n58286 = P1_P1_REIP_REG_30_ & n58261;
  assign n58287 = ~P1_P1_REIP_REG_31_ & n58286;
  assign n58288 = P1_P1_REIP_REG_31_ & ~n58286;
  assign n58289 = ~n58287 & ~n58288;
  assign n58290 = n57455 & ~n58289;
  assign n58291 = P1_P1_EBX_REG_31_ & ~n57442;
  assign n58292 = n57444 & ~n58289;
  assign n58293 = P1_P1_EBX_REG_31_ & n58268;
  assign n58294 = ~P1_P1_EBX_REG_31_ & ~n58268;
  assign n58295 = ~n58293 & ~n58294;
  assign n58296 = n57446 & ~n58295;
  assign n58297 = P1_P1_REIP_REG_31_ & n57432;
  assign n58298 = P1_P1_PHYADDRPOINTER_REG_31_ & n57461;
  assign n58299 = ~n58297 & ~n58298;
  assign n58300 = ~n55500 & n57458;
  assign n58301 = n58299 & ~n58300;
  assign n58302 = ~n58296 & n58301;
  assign n58303 = ~n55500 & n58281;
  assign n58304 = n55500 & ~n58281;
  assign n58305 = ~n58303 & ~n58304;
  assign n58306 = n57464 & ~n58305;
  assign n58307 = ~n58290 & ~n58291;
  assign n58308 = ~n58292 & n58307;
  assign n58309 = n58302 & n58308;
  assign n9906 = n58306 | ~n58309;
  assign n58311 = ~P1_P1_DATAWIDTH_REG_1_ & ~P1_P1_REIP_REG_1_;
  assign n58312 = ~P1_P1_DATAWIDTH_REG_30_ & ~P1_P1_DATAWIDTH_REG_31_;
  assign n58313 = P1_P1_DATAWIDTH_REG_0_ & P1_P1_DATAWIDTH_REG_1_;
  assign n58314 = ~P1_P1_DATAWIDTH_REG_28_ & ~P1_P1_DATAWIDTH_REG_29_;
  assign n58315 = ~P1_P1_DATAWIDTH_REG_26_ & ~P1_P1_DATAWIDTH_REG_27_;
  assign n58316 = n58312 & ~n58313;
  assign n58317 = n58314 & n58316;
  assign n58318 = n58315 & n58317;
  assign n58319 = ~P1_P1_DATAWIDTH_REG_22_ & ~P1_P1_DATAWIDTH_REG_23_;
  assign n58320 = ~P1_P1_DATAWIDTH_REG_24_ & n58319;
  assign n58321 = ~P1_P1_DATAWIDTH_REG_25_ & n58320;
  assign n58322 = ~P1_P1_DATAWIDTH_REG_18_ & ~P1_P1_DATAWIDTH_REG_19_;
  assign n58323 = ~P1_P1_DATAWIDTH_REG_20_ & n58322;
  assign n58324 = ~P1_P1_DATAWIDTH_REG_21_ & n58323;
  assign n58325 = n58321 & n58324;
  assign n58326 = ~P1_P1_DATAWIDTH_REG_14_ & ~P1_P1_DATAWIDTH_REG_15_;
  assign n58327 = ~P1_P1_DATAWIDTH_REG_16_ & n58326;
  assign n58328 = ~P1_P1_DATAWIDTH_REG_17_ & n58327;
  assign n58329 = ~P1_P1_DATAWIDTH_REG_10_ & ~P1_P1_DATAWIDTH_REG_11_;
  assign n58330 = ~P1_P1_DATAWIDTH_REG_12_ & n58329;
  assign n58331 = ~P1_P1_DATAWIDTH_REG_13_ & n58330;
  assign n58332 = n58328 & n58331;
  assign n58333 = ~P1_P1_DATAWIDTH_REG_6_ & ~P1_P1_DATAWIDTH_REG_7_;
  assign n58334 = ~P1_P1_DATAWIDTH_REG_8_ & n58333;
  assign n58335 = ~P1_P1_DATAWIDTH_REG_9_ & n58334;
  assign n58336 = ~P1_P1_DATAWIDTH_REG_2_ & ~P1_P1_DATAWIDTH_REG_3_;
  assign n58337 = ~P1_P1_DATAWIDTH_REG_4_ & n58336;
  assign n58338 = ~P1_P1_DATAWIDTH_REG_5_ & n58337;
  assign n58339 = n58335 & n58338;
  assign n58340 = n58318 & n58325;
  assign n58341 = n58332 & n58340;
  assign n58342 = n58339 & n58341;
  assign n58343 = n58311 & n58342;
  assign n58344 = P1_P1_BYTEENABLE_REG_3_ & ~n58342;
  assign n58345 = ~P1_P1_DATAWIDTH_REG_0_ & ~P1_P1_REIP_REG_0_;
  assign n58346 = ~P1_P1_DATAWIDTH_REG_1_ & n58345;
  assign n58347 = n58342 & n58346;
  assign n58348 = ~n58343 & ~n58344;
  assign n9911 = n58347 | ~n58348;
  assign n58350 = P1_P1_REIP_REG_0_ & P1_P1_REIP_REG_1_;
  assign n58351 = P1_P1_DATAWIDTH_REG_0_ & ~P1_P1_REIP_REG_0_;
  assign n58352 = ~P1_P1_DATAWIDTH_REG_0_ & ~P1_P1_DATAWIDTH_REG_1_;
  assign n58353 = ~n58351 & ~n58352;
  assign n58354 = ~P1_P1_REIP_REG_1_ & ~n58353;
  assign n58355 = ~n58350 & ~n58354;
  assign n58356 = n58342 & ~n58355;
  assign n58357 = P1_P1_BYTEENABLE_REG_2_ & ~n58342;
  assign n9916 = n58356 | n58357;
  assign n58359 = P1_P1_REIP_REG_1_ & n58342;
  assign n58360 = P1_P1_BYTEENABLE_REG_1_ & ~n58342;
  assign n58361 = ~n58359 & ~n58360;
  assign n9921 = n58347 | ~n58361;
  assign n58363 = ~P1_P1_REIP_REG_0_ & ~P1_P1_REIP_REG_1_;
  assign n58364 = n58342 & ~n58363;
  assign n58365 = P1_P1_BYTEENABLE_REG_0_ & ~n58342;
  assign n9926 = n58364 | n58365;
  assign n58367 = P1_P1_W_R_N_REG & ~n43082;
  assign n58368 = ~P1_P1_READREQUEST_REG & n43082;
  assign n9931 = n58367 | n58368;
  assign n58370 = n43746 & n43979;
  assign n58371 = ~n43694 & n43979;
  assign n58372 = P1_P1_FLUSH_REG & ~n58371;
  assign n9936 = n58370 | n58372;
  assign n58374 = P1_P1_MORE_REG & ~n58371;
  assign n58375 = ~n43740 & n58371;
  assign n9941 = n58374 | n58375;
  assign n58377 = BS & ~n43299;
  assign n58378 = P1_P1_STATEBS16_REG & n43299;
  assign n58379 = ~P1_P1_STATE_REG_0_ & n43254;
  assign n58380 = ~n58377 & ~n58378;
  assign n9946 = n58379 | ~n58380;
  assign n58382 = ~n43624 & ~n43697;
  assign n58383 = ~n43342 & ~n58382;
  assign n58384 = ~P1_P1_STATEBS16_REG & n43624;
  assign n58385 = ~n43251 & ~n58384;
  assign n58386 = P1_P1_STATE2_REG_2_ & ~n58383;
  assign n58387 = n58385 & n58386;
  assign n58388 = P1_P1_STATE2_REG_0_ & ~n58387;
  assign n58389 = ~n43995 & ~n58388;
  assign n58390 = ~n43251 & n43336;
  assign n58391 = ~n43985 & ~n58390;
  assign n58392 = ~P1_P1_STATE2_REG_0_ & ~n58391;
  assign n58393 = ~n44057 & ~n58392;
  assign n58394 = ~n57431 & n58393;
  assign n58395 = ~n58389 & ~n58394;
  assign n58396 = P1_P1_REQUESTPENDING_REG & n58394;
  assign n9951 = n58395 | n58396;
  assign n58398 = P1_P1_D_C_N_REG & ~n43082;
  assign n58399 = ~P1_P1_CODEFETCH_REG & n43082;
  assign n58400 = ~n58398 & ~n58399;
  assign n9956 = n58379 | ~n58400;
  assign n58402 = P1_P1_MEMORYFETCH_REG & n43082;
  assign n58403 = P1_P1_M_IO_N_REG & ~n43082;
  assign n9961 = n58402 | n58403;
  assign n58405 = P1_P1_STATE2_REG_0_ & n51898;
  assign n58406 = n43693 & n43979;
  assign n58407 = P1_P1_CODEFETCH_REG & ~n58406;
  assign n9966 = n58405 | n58407;
  assign n58409 = P1_P1_STATE_REG_0_ & P1_P1_ADS_N_REG;
  assign n9971 = ~n43299 | n58409;
  assign n58411 = P1_P1_STATE2_REG_2_ & ~n43706;
  assign n58412 = ~n43701 & n58411;
  assign n58413 = ~n51898 & ~n57431;
  assign n58414 = ~n58412 & ~n58413;
  assign n58415 = P1_P1_READREQUEST_REG & n58413;
  assign n9976 = n58414 | n58415;
  assign n58417 = P1_P1_STATE2_REG_2_ & n43623;
  assign n58418 = ~n58413 & ~n58417;
  assign n58419 = P1_P1_MEMORYFETCH_REG & n58413;
  assign n9981 = n58418 | n58419;
  assign n58421 = P2_P3_STATE_REG_1_ & ~P2_P3_STATE_REG_0_;
  assign n58422 = P2_P3_BYTEENABLE_REG_3_ & n58421;
  assign n58423 = P2_P3_BE_N_REG_3_ & ~n58421;
  assign n9986 = n58422 | n58423;
  assign n58425 = P2_P3_BYTEENABLE_REG_2_ & n58421;
  assign n58426 = P2_P3_BE_N_REG_2_ & ~n58421;
  assign n9991 = n58425 | n58426;
  assign n58428 = P2_P3_BYTEENABLE_REG_1_ & n58421;
  assign n58429 = P2_P3_BE_N_REG_1_ & ~n58421;
  assign n9996 = n58428 | n58429;
  assign n58431 = P2_P3_BYTEENABLE_REG_0_ & n58421;
  assign n58432 = P2_P3_BE_N_REG_0_ & ~n58421;
  assign n10001 = n58431 | n58432;
  assign n58434 = P2_P3_STATE_REG_2_ & n58421;
  assign n58435 = P2_P3_REIP_REG_30_ & n58434;
  assign n58436 = ~P2_P3_STATE_REG_2_ & n58421;
  assign n58437 = P2_P3_REIP_REG_31_ & n58436;
  assign n58438 = P2_P3_ADDRESS_REG_29_ & ~n58421;
  assign n58439 = ~n58435 & ~n58437;
  assign n10006 = n58438 | ~n58439;
  assign n58441 = P2_P3_REIP_REG_29_ & n58434;
  assign n58442 = P2_P3_REIP_REG_30_ & n58436;
  assign n58443 = P2_P3_ADDRESS_REG_28_ & ~n58421;
  assign n58444 = ~n58441 & ~n58442;
  assign n10011 = n58443 | ~n58444;
  assign n58446 = P2_P3_REIP_REG_28_ & n58434;
  assign n58447 = P2_P3_REIP_REG_29_ & n58436;
  assign n58448 = P2_P3_ADDRESS_REG_27_ & ~n58421;
  assign n58449 = ~n58446 & ~n58447;
  assign n10016 = n58448 | ~n58449;
  assign n58451 = P2_P3_REIP_REG_27_ & n58434;
  assign n58452 = P2_P3_REIP_REG_28_ & n58436;
  assign n58453 = P2_P3_ADDRESS_REG_26_ & ~n58421;
  assign n58454 = ~n58451 & ~n58452;
  assign n10021 = n58453 | ~n58454;
  assign n58456 = P2_P3_REIP_REG_26_ & n58434;
  assign n58457 = P2_P3_REIP_REG_27_ & n58436;
  assign n58458 = P2_P3_ADDRESS_REG_25_ & ~n58421;
  assign n58459 = ~n58456 & ~n58457;
  assign n10026 = n58458 | ~n58459;
  assign n58461 = P2_P3_REIP_REG_25_ & n58434;
  assign n58462 = P2_P3_REIP_REG_26_ & n58436;
  assign n58463 = P2_P3_ADDRESS_REG_24_ & ~n58421;
  assign n58464 = ~n58461 & ~n58462;
  assign n10031 = n58463 | ~n58464;
  assign n58466 = P2_P3_REIP_REG_24_ & n58434;
  assign n58467 = P2_P3_REIP_REG_25_ & n58436;
  assign n58468 = P2_P3_ADDRESS_REG_23_ & ~n58421;
  assign n58469 = ~n58466 & ~n58467;
  assign n10036 = n58468 | ~n58469;
  assign n58471 = P2_P3_REIP_REG_23_ & n58434;
  assign n58472 = P2_P3_REIP_REG_24_ & n58436;
  assign n58473 = P2_P3_ADDRESS_REG_22_ & ~n58421;
  assign n58474 = ~n58471 & ~n58472;
  assign n10041 = n58473 | ~n58474;
  assign n58476 = P2_P3_REIP_REG_22_ & n58434;
  assign n58477 = P2_P3_REIP_REG_23_ & n58436;
  assign n58478 = P2_P3_ADDRESS_REG_21_ & ~n58421;
  assign n58479 = ~n58476 & ~n58477;
  assign n10046 = n58478 | ~n58479;
  assign n58481 = P2_P3_REIP_REG_21_ & n58434;
  assign n58482 = P2_P3_REIP_REG_22_ & n58436;
  assign n58483 = P2_P3_ADDRESS_REG_20_ & ~n58421;
  assign n58484 = ~n58481 & ~n58482;
  assign n10051 = n58483 | ~n58484;
  assign n58486 = P2_P3_REIP_REG_20_ & n58434;
  assign n58487 = P2_P3_REIP_REG_21_ & n58436;
  assign n58488 = P2_P3_ADDRESS_REG_19_ & ~n58421;
  assign n58489 = ~n58486 & ~n58487;
  assign n10056 = n58488 | ~n58489;
  assign n58491 = P2_P3_REIP_REG_19_ & n58434;
  assign n58492 = P2_P3_REIP_REG_20_ & n58436;
  assign n58493 = P2_P3_ADDRESS_REG_18_ & ~n58421;
  assign n58494 = ~n58491 & ~n58492;
  assign n10061 = n58493 | ~n58494;
  assign n58496 = P2_P3_REIP_REG_18_ & n58434;
  assign n58497 = P2_P3_REIP_REG_19_ & n58436;
  assign n58498 = P2_P3_ADDRESS_REG_17_ & ~n58421;
  assign n58499 = ~n58496 & ~n58497;
  assign n10066 = n58498 | ~n58499;
  assign n58501 = P2_P3_REIP_REG_17_ & n58434;
  assign n58502 = P2_P3_REIP_REG_18_ & n58436;
  assign n58503 = P2_P3_ADDRESS_REG_16_ & ~n58421;
  assign n58504 = ~n58501 & ~n58502;
  assign n10071 = n58503 | ~n58504;
  assign n58506 = P2_P3_REIP_REG_16_ & n58434;
  assign n58507 = P2_P3_REIP_REG_17_ & n58436;
  assign n58508 = P2_P3_ADDRESS_REG_15_ & ~n58421;
  assign n58509 = ~n58506 & ~n58507;
  assign n10076 = n58508 | ~n58509;
  assign n58511 = P2_P3_REIP_REG_15_ & n58434;
  assign n58512 = P2_P3_REIP_REG_16_ & n58436;
  assign n58513 = P2_P3_ADDRESS_REG_14_ & ~n58421;
  assign n58514 = ~n58511 & ~n58512;
  assign n10081 = n58513 | ~n58514;
  assign n58516 = P2_P3_REIP_REG_14_ & n58434;
  assign n58517 = P2_P3_REIP_REG_15_ & n58436;
  assign n58518 = P2_P3_ADDRESS_REG_13_ & ~n58421;
  assign n58519 = ~n58516 & ~n58517;
  assign n10086 = n58518 | ~n58519;
  assign n58521 = P2_P3_REIP_REG_13_ & n58434;
  assign n58522 = P2_P3_REIP_REG_14_ & n58436;
  assign n58523 = P2_P3_ADDRESS_REG_12_ & ~n58421;
  assign n58524 = ~n58521 & ~n58522;
  assign n10091 = n58523 | ~n58524;
  assign n58526 = P2_P3_REIP_REG_12_ & n58434;
  assign n58527 = P2_P3_REIP_REG_13_ & n58436;
  assign n58528 = P2_P3_ADDRESS_REG_11_ & ~n58421;
  assign n58529 = ~n58526 & ~n58527;
  assign n10096 = n58528 | ~n58529;
  assign n58531 = P2_P3_REIP_REG_11_ & n58434;
  assign n58532 = P2_P3_REIP_REG_12_ & n58436;
  assign n58533 = P2_P3_ADDRESS_REG_10_ & ~n58421;
  assign n58534 = ~n58531 & ~n58532;
  assign n10101 = n58533 | ~n58534;
  assign n58536 = P2_P3_REIP_REG_10_ & n58434;
  assign n58537 = P2_P3_REIP_REG_11_ & n58436;
  assign n58538 = P2_P3_ADDRESS_REG_9_ & ~n58421;
  assign n58539 = ~n58536 & ~n58537;
  assign n10106 = n58538 | ~n58539;
  assign n58541 = P2_P3_REIP_REG_9_ & n58434;
  assign n58542 = P2_P3_REIP_REG_10_ & n58436;
  assign n58543 = P2_P3_ADDRESS_REG_8_ & ~n58421;
  assign n58544 = ~n58541 & ~n58542;
  assign n10111 = n58543 | ~n58544;
  assign n58546 = P2_P3_REIP_REG_8_ & n58434;
  assign n58547 = P2_P3_REIP_REG_9_ & n58436;
  assign n58548 = P2_P3_ADDRESS_REG_7_ & ~n58421;
  assign n58549 = ~n58546 & ~n58547;
  assign n10116 = n58548 | ~n58549;
  assign n58551 = P2_P3_REIP_REG_7_ & n58434;
  assign n58552 = P2_P3_REIP_REG_8_ & n58436;
  assign n58553 = P2_P3_ADDRESS_REG_6_ & ~n58421;
  assign n58554 = ~n58551 & ~n58552;
  assign n10121 = n58553 | ~n58554;
  assign n58556 = P2_P3_REIP_REG_6_ & n58434;
  assign n58557 = P2_P3_REIP_REG_7_ & n58436;
  assign n58558 = P2_P3_ADDRESS_REG_5_ & ~n58421;
  assign n58559 = ~n58556 & ~n58557;
  assign n10126 = n58558 | ~n58559;
  assign n58561 = P2_P3_REIP_REG_5_ & n58434;
  assign n58562 = P2_P3_REIP_REG_6_ & n58436;
  assign n58563 = P2_P3_ADDRESS_REG_4_ & ~n58421;
  assign n58564 = ~n58561 & ~n58562;
  assign n10131 = n58563 | ~n58564;
  assign n58566 = P2_P3_REIP_REG_4_ & n58434;
  assign n58567 = P2_P3_REIP_REG_5_ & n58436;
  assign n58568 = P2_P3_ADDRESS_REG_3_ & ~n58421;
  assign n58569 = ~n58566 & ~n58567;
  assign n10136 = n58568 | ~n58569;
  assign n58571 = P2_P3_REIP_REG_3_ & n58434;
  assign n58572 = P2_P3_REIP_REG_4_ & n58436;
  assign n58573 = P2_P3_ADDRESS_REG_2_ & ~n58421;
  assign n58574 = ~n58571 & ~n58572;
  assign n10141 = n58573 | ~n58574;
  assign n58576 = P2_P3_REIP_REG_2_ & n58434;
  assign n58577 = P2_P3_REIP_REG_3_ & n58436;
  assign n58578 = P2_P3_ADDRESS_REG_1_ & ~n58421;
  assign n58579 = ~n58576 & ~n58577;
  assign n10146 = n58578 | ~n58579;
  assign n58581 = P2_P3_REIP_REG_1_ & n58434;
  assign n58582 = P2_P3_REIP_REG_2_ & n58436;
  assign n58583 = P2_P3_ADDRESS_REG_0_ & ~n58421;
  assign n58584 = ~n58581 & ~n58582;
  assign n10151 = n58583 | ~n58584;
  assign n58586 = ~P2_P3_STATE_REG_2_ & P2_P3_STATE_REG_1_;
  assign n58587 = NA & n58586;
  assign n58588 = P2_P3_STATE_REG_0_ & ~n58587;
  assign n58589 = ~HOLD & ~P2_P3_REQUESTPENDING_REG;
  assign n58590 = P2_P3_D_C_N_REG & ~P2_P3_ADS_N_REG;
  assign n58591 = P2_P3_M_IO_N_REG & n58590;
  assign n58592 = P2_P3_W_R_N_REG & n58591;
  assign n58593 = P4_RD_REG & n58592;
  assign n58594 = P2_READY22_REG & ~n58593;
  assign n58595 = n58586 & ~n58589;
  assign n58596 = n58594 & n58595;
  assign n58597 = ~P2_P3_STATE_REG_2_ & ~P2_P3_STATE_REG_1_;
  assign n58598 = HOLD & ~P2_P3_REQUESTPENDING_REG;
  assign n58599 = n58597 & n58598;
  assign n58600 = ~n58596 & ~n58599;
  assign n58601 = n58588 & ~n58600;
  assign n58602 = ~n58434 & ~n58601;
  assign n58603 = ~HOLD & P2_P3_REQUESTPENDING_REG;
  assign n58604 = P2_P3_STATE_REG_0_ & ~n58603;
  assign n58605 = ~n58589 & n58604;
  assign n58606 = ~NA & ~P2_P3_STATE_REG_0_;
  assign n58607 = n58589 & ~n58594;
  assign n58608 = ~n58594 & n58603;
  assign n58609 = ~n58607 & ~n58608;
  assign n58610 = P2_P3_STATE_REG_1_ & n58609;
  assign n58611 = ~n58605 & ~n58606;
  assign n58612 = ~n58610 & n58611;
  assign n58613 = P2_P3_STATE_REG_2_ & ~n58612;
  assign n10156 = ~n58602 | n58613;
  assign n58615 = P2_P3_STATE_REG_2_ & ~n58604;
  assign n58616 = P2_P3_STATE_REG_0_ & P2_P3_REQUESTPENDING_REG;
  assign n58617 = ~P2_P3_STATE_REG_2_ & n58616;
  assign n58618 = ~n58615 & ~n58617;
  assign n58619 = ~P2_P3_STATE_REG_1_ & ~n58618;
  assign n58620 = HOLD & ~n58594;
  assign n58621 = P2_P3_STATE_REG_0_ & ~n58620;
  assign n58622 = P2_P3_STATE_REG_2_ & ~n58621;
  assign n58623 = ~n58607 & ~n58622;
  assign n58624 = P2_P3_STATE_REG_1_ & n58623;
  assign n58625 = n58421 & n58594;
  assign n58626 = ~n58436 & ~n58625;
  assign n58627 = ~n58619 & ~n58624;
  assign n10161 = ~n58626 | ~n58627;
  assign n58629 = P2_P3_STATE_REG_1_ & ~n58608;
  assign n58630 = n58616 & ~n58629;
  assign n58631 = ~P2_P3_STATE_REG_2_ & ~n58630;
  assign n58632 = P2_P3_STATE_REG_2_ & n58604;
  assign n58633 = NA & ~P2_P3_STATE_REG_0_;
  assign n58634 = P2_P3_STATE_REG_2_ & ~n58603;
  assign n58635 = ~n58633 & ~n58634;
  assign n58636 = ~P2_P3_STATE_REG_1_ & ~n58635;
  assign n58637 = ~n58631 & ~n58632;
  assign n10166 = n58636 | ~n58637;
  assign n58639 = ~BS & ~n58597;
  assign n58640 = P2_P3_STATE_REG_0_ & n58586;
  assign n58641 = ~P2_P3_STATE_REG_1_ & ~P2_P3_STATE_REG_0_;
  assign n58642 = ~n58640 & ~n58641;
  assign n58643 = n58639 & ~n58642;
  assign n58644 = P2_P3_DATAWIDTH_REG_0_ & n58642;
  assign n10171 = n58643 | n58644;
  assign n58646 = P2_P3_DATAWIDTH_REG_1_ & n58642;
  assign n58647 = ~n58639 & ~n58642;
  assign n10176 = n58646 | n58647;
  assign n10181 = P2_P3_DATAWIDTH_REG_2_ & n58642;
  assign n10186 = P2_P3_DATAWIDTH_REG_3_ & n58642;
  assign n10191 = P2_P3_DATAWIDTH_REG_4_ & n58642;
  assign n10196 = P2_P3_DATAWIDTH_REG_5_ & n58642;
  assign n10201 = P2_P3_DATAWIDTH_REG_6_ & n58642;
  assign n10206 = P2_P3_DATAWIDTH_REG_7_ & n58642;
  assign n10211 = P2_P3_DATAWIDTH_REG_8_ & n58642;
  assign n10216 = P2_P3_DATAWIDTH_REG_9_ & n58642;
  assign n10221 = P2_P3_DATAWIDTH_REG_10_ & n58642;
  assign n10226 = P2_P3_DATAWIDTH_REG_11_ & n58642;
  assign n10231 = P2_P3_DATAWIDTH_REG_12_ & n58642;
  assign n10236 = P2_P3_DATAWIDTH_REG_13_ & n58642;
  assign n10241 = P2_P3_DATAWIDTH_REG_14_ & n58642;
  assign n10246 = P2_P3_DATAWIDTH_REG_15_ & n58642;
  assign n10251 = P2_P3_DATAWIDTH_REG_16_ & n58642;
  assign n10256 = P2_P3_DATAWIDTH_REG_17_ & n58642;
  assign n10261 = P2_P3_DATAWIDTH_REG_18_ & n58642;
  assign n10266 = P2_P3_DATAWIDTH_REG_19_ & n58642;
  assign n10271 = P2_P3_DATAWIDTH_REG_20_ & n58642;
  assign n10276 = P2_P3_DATAWIDTH_REG_21_ & n58642;
  assign n10281 = P2_P3_DATAWIDTH_REG_22_ & n58642;
  assign n10286 = P2_P3_DATAWIDTH_REG_23_ & n58642;
  assign n10291 = P2_P3_DATAWIDTH_REG_24_ & n58642;
  assign n10296 = P2_P3_DATAWIDTH_REG_25_ & n58642;
  assign n10301 = P2_P3_DATAWIDTH_REG_26_ & n58642;
  assign n10306 = P2_P3_DATAWIDTH_REG_27_ & n58642;
  assign n10311 = P2_P3_DATAWIDTH_REG_28_ & n58642;
  assign n10316 = P2_P3_DATAWIDTH_REG_29_ & n58642;
  assign n10321 = P2_P3_DATAWIDTH_REG_30_ & n58642;
  assign n10326 = P2_P3_DATAWIDTH_REG_31_ & n58642;
  assign n58679 = P2_P3_STATE2_REG_2_ & P2_P3_STATE2_REG_1_;
  assign n58680 = P2_P3_STATE2_REG_1_ & n58594;
  assign n58681 = ~P2_P3_STATE2_REG_0_ & ~n58680;
  assign n58682 = ~P2_P3_STATEBS16_REG & ~n58594;
  assign n58683 = P2_P3_STATE_REG_2_ & ~P2_P3_STATE_REG_1_;
  assign n58684 = ~n58586 & ~n58683;
  assign n58685 = ~P2_P3_STATE_REG_0_ & ~n58684;
  assign n58686 = n58682 & n58685;
  assign n58687 = P2_P3_INSTQUEUERD_ADDR_REG_1_ & P2_P3_INSTQUEUERD_ADDR_REG_0_;
  assign n58688 = ~P2_P3_INSTQUEUERD_ADDR_REG_2_ & n58687;
  assign n58689 = P2_P3_INSTQUEUERD_ADDR_REG_3_ & n58688;
  assign n58690 = P2_P3_INSTQUEUE_REG_11__5_ & n58689;
  assign n58691 = P2_P3_INSTQUEUERD_ADDR_REG_1_ & ~P2_P3_INSTQUEUERD_ADDR_REG_0_;
  assign n58692 = ~P2_P3_INSTQUEUERD_ADDR_REG_2_ & n58691;
  assign n58693 = P2_P3_INSTQUEUERD_ADDR_REG_3_ & n58692;
  assign n58694 = P2_P3_INSTQUEUE_REG_10__5_ & n58693;
  assign n58695 = ~n58690 & ~n58694;
  assign n58696 = ~P2_P3_INSTQUEUERD_ADDR_REG_1_ & P2_P3_INSTQUEUERD_ADDR_REG_0_;
  assign n58697 = ~P2_P3_INSTQUEUERD_ADDR_REG_2_ & n58696;
  assign n58698 = P2_P3_INSTQUEUERD_ADDR_REG_3_ & n58697;
  assign n58699 = P2_P3_INSTQUEUE_REG_9__5_ & n58698;
  assign n58700 = ~P2_P3_INSTQUEUERD_ADDR_REG_1_ & ~P2_P3_INSTQUEUERD_ADDR_REG_0_;
  assign n58701 = ~P2_P3_INSTQUEUERD_ADDR_REG_2_ & n58700;
  assign n58702 = P2_P3_INSTQUEUERD_ADDR_REG_3_ & n58701;
  assign n58703 = P2_P3_INSTQUEUE_REG_8__5_ & n58702;
  assign n58704 = ~n58699 & ~n58703;
  assign n58705 = P2_P3_INSTQUEUERD_ADDR_REG_3_ & P2_P3_INSTQUEUERD_ADDR_REG_2_;
  assign n58706 = n58687 & n58705;
  assign n58707 = P2_P3_INSTQUEUE_REG_15__5_ & n58706;
  assign n58708 = n58691 & n58705;
  assign n58709 = P2_P3_INSTQUEUE_REG_14__5_ & n58708;
  assign n58710 = n58696 & n58705;
  assign n58711 = P2_P3_INSTQUEUE_REG_13__5_ & n58710;
  assign n58712 = n58700 & n58705;
  assign n58713 = P2_P3_INSTQUEUE_REG_12__5_ & n58712;
  assign n58714 = ~n58707 & ~n58709;
  assign n58715 = ~n58711 & n58714;
  assign n58716 = ~n58713 & n58715;
  assign n58717 = ~P2_P3_INSTQUEUERD_ADDR_REG_3_ & P2_P3_INSTQUEUERD_ADDR_REG_2_;
  assign n58718 = n58687 & n58717;
  assign n58719 = P2_P3_INSTQUEUE_REG_7__5_ & n58718;
  assign n58720 = n58691 & n58717;
  assign n58721 = P2_P3_INSTQUEUE_REG_6__5_ & n58720;
  assign n58722 = n58696 & n58717;
  assign n58723 = P2_P3_INSTQUEUE_REG_5__5_ & n58722;
  assign n58724 = n58700 & n58717;
  assign n58725 = P2_P3_INSTQUEUE_REG_4__5_ & n58724;
  assign n58726 = ~n58719 & ~n58721;
  assign n58727 = ~n58723 & n58726;
  assign n58728 = ~n58725 & n58727;
  assign n58729 = ~P2_P3_INSTQUEUERD_ADDR_REG_3_ & n58688;
  assign n58730 = P2_P3_INSTQUEUE_REG_3__5_ & n58729;
  assign n58731 = ~P2_P3_INSTQUEUERD_ADDR_REG_3_ & ~P2_P3_INSTQUEUERD_ADDR_REG_2_;
  assign n58732 = n58691 & n58731;
  assign n58733 = P2_P3_INSTQUEUE_REG_2__5_ & n58732;
  assign n58734 = n58696 & n58731;
  assign n58735 = P2_P3_INSTQUEUE_REG_1__5_ & n58734;
  assign n58736 = ~P2_P3_INSTQUEUERD_ADDR_REG_3_ & n58701;
  assign n58737 = P2_P3_INSTQUEUE_REG_0__5_ & n58736;
  assign n58738 = ~n58730 & ~n58733;
  assign n58739 = ~n58735 & n58738;
  assign n58740 = ~n58737 & n58739;
  assign n58741 = n58695 & n58704;
  assign n58742 = n58716 & n58741;
  assign n58743 = n58728 & n58742;
  assign n58744 = n58740 & n58743;
  assign n58745 = P2_P3_INSTQUEUE_REG_11__6_ & n58689;
  assign n58746 = P2_P3_INSTQUEUE_REG_10__6_ & n58693;
  assign n58747 = ~n58745 & ~n58746;
  assign n58748 = P2_P3_INSTQUEUE_REG_9__6_ & n58698;
  assign n58749 = P2_P3_INSTQUEUE_REG_8__6_ & n58702;
  assign n58750 = ~n58748 & ~n58749;
  assign n58751 = P2_P3_INSTQUEUE_REG_15__6_ & n58706;
  assign n58752 = P2_P3_INSTQUEUE_REG_14__6_ & n58708;
  assign n58753 = P2_P3_INSTQUEUE_REG_13__6_ & n58710;
  assign n58754 = P2_P3_INSTQUEUE_REG_12__6_ & n58712;
  assign n58755 = ~n58751 & ~n58752;
  assign n58756 = ~n58753 & n58755;
  assign n58757 = ~n58754 & n58756;
  assign n58758 = P2_P3_INSTQUEUE_REG_7__6_ & n58718;
  assign n58759 = P2_P3_INSTQUEUE_REG_6__6_ & n58720;
  assign n58760 = P2_P3_INSTQUEUE_REG_5__6_ & n58722;
  assign n58761 = P2_P3_INSTQUEUE_REG_4__6_ & n58724;
  assign n58762 = ~n58758 & ~n58759;
  assign n58763 = ~n58760 & n58762;
  assign n58764 = ~n58761 & n58763;
  assign n58765 = P2_P3_INSTQUEUE_REG_3__6_ & n58729;
  assign n58766 = P2_P3_INSTQUEUE_REG_2__6_ & n58732;
  assign n58767 = P2_P3_INSTQUEUE_REG_1__6_ & n58734;
  assign n58768 = P2_P3_INSTQUEUE_REG_0__6_ & n58736;
  assign n58769 = ~n58765 & ~n58766;
  assign n58770 = ~n58767 & n58769;
  assign n58771 = ~n58768 & n58770;
  assign n58772 = n58747 & n58750;
  assign n58773 = n58757 & n58772;
  assign n58774 = n58764 & n58773;
  assign n58775 = n58771 & n58774;
  assign n58776 = n58744 & n58775;
  assign n58777 = P2_P3_INSTQUEUE_REG_11__4_ & n58689;
  assign n58778 = P2_P3_INSTQUEUE_REG_10__4_ & n58693;
  assign n58779 = ~n58777 & ~n58778;
  assign n58780 = P2_P3_INSTQUEUE_REG_9__4_ & n58698;
  assign n58781 = P2_P3_INSTQUEUE_REG_8__4_ & n58702;
  assign n58782 = ~n58780 & ~n58781;
  assign n58783 = P2_P3_INSTQUEUE_REG_15__4_ & n58706;
  assign n58784 = P2_P3_INSTQUEUE_REG_14__4_ & n58708;
  assign n58785 = P2_P3_INSTQUEUE_REG_13__4_ & n58710;
  assign n58786 = P2_P3_INSTQUEUE_REG_12__4_ & n58712;
  assign n58787 = ~n58783 & ~n58784;
  assign n58788 = ~n58785 & n58787;
  assign n58789 = ~n58786 & n58788;
  assign n58790 = P2_P3_INSTQUEUE_REG_7__4_ & n58718;
  assign n58791 = P2_P3_INSTQUEUE_REG_6__4_ & n58720;
  assign n58792 = P2_P3_INSTQUEUE_REG_5__4_ & n58722;
  assign n58793 = P2_P3_INSTQUEUE_REG_4__4_ & n58724;
  assign n58794 = ~n58790 & ~n58791;
  assign n58795 = ~n58792 & n58794;
  assign n58796 = ~n58793 & n58795;
  assign n58797 = P2_P3_INSTQUEUE_REG_3__4_ & n58729;
  assign n58798 = P2_P3_INSTQUEUE_REG_2__4_ & n58732;
  assign n58799 = P2_P3_INSTQUEUE_REG_1__4_ & n58734;
  assign n58800 = P2_P3_INSTQUEUE_REG_0__4_ & n58736;
  assign n58801 = ~n58797 & ~n58798;
  assign n58802 = ~n58799 & n58801;
  assign n58803 = ~n58800 & n58802;
  assign n58804 = n58779 & n58782;
  assign n58805 = n58789 & n58804;
  assign n58806 = n58796 & n58805;
  assign n58807 = n58803 & n58806;
  assign n58808 = P2_P3_INSTQUEUE_REG_11__7_ & n58689;
  assign n58809 = P2_P3_INSTQUEUE_REG_10__7_ & n58693;
  assign n58810 = ~n58808 & ~n58809;
  assign n58811 = P2_P3_INSTQUEUE_REG_9__7_ & n58698;
  assign n58812 = P2_P3_INSTQUEUE_REG_8__7_ & n58702;
  assign n58813 = ~n58811 & ~n58812;
  assign n58814 = P2_P3_INSTQUEUE_REG_15__7_ & n58706;
  assign n58815 = P2_P3_INSTQUEUE_REG_14__7_ & n58708;
  assign n58816 = P2_P3_INSTQUEUE_REG_13__7_ & n58710;
  assign n58817 = P2_P3_INSTQUEUE_REG_12__7_ & n58712;
  assign n58818 = ~n58814 & ~n58815;
  assign n58819 = ~n58816 & n58818;
  assign n58820 = ~n58817 & n58819;
  assign n58821 = P2_P3_INSTQUEUE_REG_7__7_ & n58718;
  assign n58822 = P2_P3_INSTQUEUE_REG_6__7_ & n58720;
  assign n58823 = P2_P3_INSTQUEUE_REG_5__7_ & n58722;
  assign n58824 = P2_P3_INSTQUEUE_REG_4__7_ & n58724;
  assign n58825 = ~n58821 & ~n58822;
  assign n58826 = ~n58823 & n58825;
  assign n58827 = ~n58824 & n58826;
  assign n58828 = P2_P3_INSTQUEUE_REG_3__7_ & n58729;
  assign n58829 = P2_P3_INSTQUEUE_REG_2__7_ & n58732;
  assign n58830 = P2_P3_INSTQUEUE_REG_1__7_ & n58734;
  assign n58831 = P2_P3_INSTQUEUE_REG_0__7_ & n58736;
  assign n58832 = ~n58828 & ~n58829;
  assign n58833 = ~n58830 & n58832;
  assign n58834 = ~n58831 & n58833;
  assign n58835 = n58810 & n58813;
  assign n58836 = n58820 & n58835;
  assign n58837 = n58827 & n58836;
  assign n58838 = n58834 & n58837;
  assign n58839 = P2_P3_INSTQUEUE_REG_11__3_ & n58689;
  assign n58840 = P2_P3_INSTQUEUE_REG_10__3_ & n58693;
  assign n58841 = ~n58839 & ~n58840;
  assign n58842 = P2_P3_INSTQUEUE_REG_9__3_ & n58698;
  assign n58843 = P2_P3_INSTQUEUE_REG_8__3_ & n58702;
  assign n58844 = ~n58842 & ~n58843;
  assign n58845 = P2_P3_INSTQUEUE_REG_15__3_ & n58706;
  assign n58846 = P2_P3_INSTQUEUE_REG_14__3_ & n58708;
  assign n58847 = P2_P3_INSTQUEUE_REG_13__3_ & n58710;
  assign n58848 = P2_P3_INSTQUEUE_REG_12__3_ & n58712;
  assign n58849 = ~n58845 & ~n58846;
  assign n58850 = ~n58847 & n58849;
  assign n58851 = ~n58848 & n58850;
  assign n58852 = P2_P3_INSTQUEUE_REG_7__3_ & n58718;
  assign n58853 = P2_P3_INSTQUEUE_REG_6__3_ & n58720;
  assign n58854 = P2_P3_INSTQUEUE_REG_5__3_ & n58722;
  assign n58855 = P2_P3_INSTQUEUE_REG_4__3_ & n58724;
  assign n58856 = ~n58852 & ~n58853;
  assign n58857 = ~n58854 & n58856;
  assign n58858 = ~n58855 & n58857;
  assign n58859 = P2_P3_INSTQUEUE_REG_3__3_ & n58729;
  assign n58860 = P2_P3_INSTQUEUE_REG_2__3_ & n58732;
  assign n58861 = P2_P3_INSTQUEUE_REG_1__3_ & n58734;
  assign n58862 = P2_P3_INSTQUEUE_REG_0__3_ & n58736;
  assign n58863 = ~n58859 & ~n58860;
  assign n58864 = ~n58861 & n58863;
  assign n58865 = ~n58862 & n58864;
  assign n58866 = n58841 & n58844;
  assign n58867 = n58851 & n58866;
  assign n58868 = n58858 & n58867;
  assign n58869 = n58865 & n58868;
  assign n58870 = P2_P3_INSTQUEUE_REG_11__2_ & n58689;
  assign n58871 = P2_P3_INSTQUEUE_REG_10__2_ & n58693;
  assign n58872 = ~n58870 & ~n58871;
  assign n58873 = P2_P3_INSTQUEUE_REG_9__2_ & n58698;
  assign n58874 = P2_P3_INSTQUEUE_REG_8__2_ & n58702;
  assign n58875 = ~n58873 & ~n58874;
  assign n58876 = P2_P3_INSTQUEUE_REG_15__2_ & n58706;
  assign n58877 = P2_P3_INSTQUEUE_REG_14__2_ & n58708;
  assign n58878 = P2_P3_INSTQUEUE_REG_13__2_ & n58710;
  assign n58879 = P2_P3_INSTQUEUE_REG_12__2_ & n58712;
  assign n58880 = ~n58876 & ~n58877;
  assign n58881 = ~n58878 & n58880;
  assign n58882 = ~n58879 & n58881;
  assign n58883 = P2_P3_INSTQUEUE_REG_7__2_ & n58718;
  assign n58884 = P2_P3_INSTQUEUE_REG_6__2_ & n58720;
  assign n58885 = P2_P3_INSTQUEUE_REG_5__2_ & n58722;
  assign n58886 = P2_P3_INSTQUEUE_REG_4__2_ & n58724;
  assign n58887 = ~n58883 & ~n58884;
  assign n58888 = ~n58885 & n58887;
  assign n58889 = ~n58886 & n58888;
  assign n58890 = P2_P3_INSTQUEUE_REG_3__2_ & n58729;
  assign n58891 = P2_P3_INSTQUEUE_REG_2__2_ & n58732;
  assign n58892 = P2_P3_INSTQUEUE_REG_1__2_ & n58734;
  assign n58893 = P2_P3_INSTQUEUE_REG_0__2_ & n58736;
  assign n58894 = ~n58890 & ~n58891;
  assign n58895 = ~n58892 & n58894;
  assign n58896 = ~n58893 & n58895;
  assign n58897 = n58872 & n58875;
  assign n58898 = n58882 & n58897;
  assign n58899 = n58889 & n58898;
  assign n58900 = n58896 & n58899;
  assign n58901 = ~n58838 & ~n58869;
  assign n58902 = n58900 & n58901;
  assign n58903 = n58776 & n58807;
  assign n58904 = n58902 & n58903;
  assign n58905 = P2_P3_INSTQUEUE_REG_11__1_ & n58689;
  assign n58906 = P2_P3_INSTQUEUE_REG_10__1_ & n58693;
  assign n58907 = ~n58905 & ~n58906;
  assign n58908 = P2_P3_INSTQUEUE_REG_9__1_ & n58698;
  assign n58909 = P2_P3_INSTQUEUE_REG_8__1_ & n58702;
  assign n58910 = ~n58908 & ~n58909;
  assign n58911 = P2_P3_INSTQUEUE_REG_15__1_ & n58706;
  assign n58912 = P2_P3_INSTQUEUE_REG_14__1_ & n58708;
  assign n58913 = P2_P3_INSTQUEUE_REG_13__1_ & n58710;
  assign n58914 = P2_P3_INSTQUEUE_REG_12__1_ & n58712;
  assign n58915 = ~n58911 & ~n58912;
  assign n58916 = ~n58913 & n58915;
  assign n58917 = ~n58914 & n58916;
  assign n58918 = P2_P3_INSTQUEUE_REG_7__1_ & n58718;
  assign n58919 = P2_P3_INSTQUEUE_REG_6__1_ & n58720;
  assign n58920 = P2_P3_INSTQUEUE_REG_5__1_ & n58722;
  assign n58921 = P2_P3_INSTQUEUE_REG_4__1_ & n58724;
  assign n58922 = ~n58918 & ~n58919;
  assign n58923 = ~n58920 & n58922;
  assign n58924 = ~n58921 & n58923;
  assign n58925 = P2_P3_INSTQUEUE_REG_3__1_ & n58729;
  assign n58926 = P2_P3_INSTQUEUE_REG_2__1_ & n58732;
  assign n58927 = P2_P3_INSTQUEUE_REG_1__1_ & n58734;
  assign n58928 = P2_P3_INSTQUEUE_REG_0__1_ & n58736;
  assign n58929 = ~n58925 & ~n58926;
  assign n58930 = ~n58927 & n58929;
  assign n58931 = ~n58928 & n58930;
  assign n58932 = n58907 & n58910;
  assign n58933 = n58917 & n58932;
  assign n58934 = n58924 & n58933;
  assign n58935 = n58931 & n58934;
  assign n58936 = P2_P3_INSTQUEUE_REG_11__0_ & n58689;
  assign n58937 = P2_P3_INSTQUEUE_REG_10__0_ & n58693;
  assign n58938 = ~n58936 & ~n58937;
  assign n58939 = P2_P3_INSTQUEUE_REG_9__0_ & n58698;
  assign n58940 = P2_P3_INSTQUEUE_REG_8__0_ & n58702;
  assign n58941 = ~n58939 & ~n58940;
  assign n58942 = P2_P3_INSTQUEUE_REG_15__0_ & n58706;
  assign n58943 = P2_P3_INSTQUEUE_REG_14__0_ & n58708;
  assign n58944 = P2_P3_INSTQUEUE_REG_13__0_ & n58710;
  assign n58945 = P2_P3_INSTQUEUE_REG_12__0_ & n58712;
  assign n58946 = ~n58942 & ~n58943;
  assign n58947 = ~n58944 & n58946;
  assign n58948 = ~n58945 & n58947;
  assign n58949 = P2_P3_INSTQUEUE_REG_7__0_ & n58718;
  assign n58950 = P2_P3_INSTQUEUE_REG_6__0_ & n58720;
  assign n58951 = P2_P3_INSTQUEUE_REG_5__0_ & n58722;
  assign n58952 = P2_P3_INSTQUEUE_REG_4__0_ & n58724;
  assign n58953 = ~n58949 & ~n58950;
  assign n58954 = ~n58951 & n58953;
  assign n58955 = ~n58952 & n58954;
  assign n58956 = P2_P3_INSTQUEUE_REG_3__0_ & n58729;
  assign n58957 = P2_P3_INSTQUEUE_REG_2__0_ & n58732;
  assign n58958 = P2_P3_INSTQUEUE_REG_1__0_ & n58734;
  assign n58959 = P2_P3_INSTQUEUE_REG_0__0_ & n58736;
  assign n58960 = ~n58956 & ~n58957;
  assign n58961 = ~n58958 & n58960;
  assign n58962 = ~n58959 & n58961;
  assign n58963 = n58938 & n58941;
  assign n58964 = n58948 & n58963;
  assign n58965 = n58955 & n58964;
  assign n58966 = n58962 & n58965;
  assign n58967 = n58935 & ~n58966;
  assign n58968 = n58904 & n58967;
  assign n58969 = n58686 & n58968;
  assign n58970 = ~P2_P3_STATE2_REG_1_ & ~n58969;
  assign n58971 = ~n58594 & n58685;
  assign n58972 = ~n58900 & ~n58935;
  assign n58973 = n58971 & n58972;
  assign n58974 = ~n58594 & ~n58900;
  assign n58975 = n58935 & n58974;
  assign n58976 = ~n58594 & n58900;
  assign n58977 = n58935 & ~n58971;
  assign n58978 = n58976 & ~n58977;
  assign n58979 = ~n58973 & ~n58975;
  assign n58980 = ~n58978 & n58979;
  assign n58981 = P2_P3_INSTQUEUERD_ADDR_REG_4_ & ~P2_P3_INSTQUEUEWR_ADDR_REG_4_;
  assign n58982 = ~P2_P3_INSTQUEUERD_ADDR_REG_3_ & P2_P3_INSTQUEUEWR_ADDR_REG_3_;
  assign n58983 = P2_P3_INSTQUEUERD_ADDR_REG_3_ & ~P2_P3_INSTQUEUEWR_ADDR_REG_3_;
  assign n58984 = ~P2_P3_INSTQUEUERD_ADDR_REG_2_ & P2_P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n58985 = P2_P3_INSTQUEUERD_ADDR_REG_2_ & ~P2_P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n58986 = P2_P3_INSTQUEUERD_ADDR_REG_0_ & ~P2_P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n58987 = P2_P3_INSTQUEUEWR_ADDR_REG_1_ & ~n58986;
  assign n58988 = ~P2_P3_INSTQUEUEWR_ADDR_REG_1_ & n58986;
  assign n58989 = ~P2_P3_INSTQUEUERD_ADDR_REG_1_ & ~n58988;
  assign n58990 = ~n58987 & ~n58989;
  assign n58991 = ~n58985 & ~n58990;
  assign n58992 = ~n58984 & ~n58991;
  assign n58993 = ~n58983 & ~n58992;
  assign n58994 = ~n58982 & ~n58993;
  assign n58995 = ~P2_P3_INSTQUEUERD_ADDR_REG_4_ & P2_P3_INSTQUEUEWR_ADDR_REG_4_;
  assign n58996 = n58994 & ~n58995;
  assign n58997 = ~n58981 & ~n58996;
  assign n58998 = ~n58981 & ~n58995;
  assign n58999 = ~n58994 & ~n58998;
  assign n59000 = n58994 & n58998;
  assign n59001 = ~n58999 & ~n59000;
  assign n59002 = ~n58982 & ~n58983;
  assign n59003 = ~n58992 & ~n59002;
  assign n59004 = n58992 & n59002;
  assign n59005 = ~n59003 & ~n59004;
  assign n59006 = ~P2_P3_INSTQUEUERD_ADDR_REG_1_ & P2_P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n59007 = P2_P3_INSTQUEUERD_ADDR_REG_1_ & ~P2_P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n59008 = ~n59006 & ~n59007;
  assign n59009 = ~n58986 & ~n59008;
  assign n59010 = n58986 & n59008;
  assign n59011 = ~n59009 & ~n59010;
  assign n59012 = ~n58984 & ~n58985;
  assign n59013 = ~n58990 & ~n59012;
  assign n59014 = n58990 & n59012;
  assign n59015 = ~n59013 & ~n59014;
  assign n59016 = n59001 & n59005;
  assign n59017 = n59011 & n59016;
  assign n59018 = n59015 & n59017;
  assign n59019 = n58997 & ~n59018;
  assign n59020 = ~n58935 & ~n59019;
  assign n59021 = n58935 & ~n59019;
  assign n59022 = ~n59020 & ~n59021;
  assign n59023 = ~n58838 & n58869;
  assign n59024 = ~n58744 & ~n58775;
  assign n59025 = n58807 & n59024;
  assign n59026 = n59023 & n59025;
  assign n59027 = n58966 & n59026;
  assign n59028 = n59022 & n59027;
  assign n59029 = ~n58900 & ~n59028;
  assign n59030 = ~n58869 & ~n58966;
  assign n59031 = ~n58838 & n59030;
  assign n59032 = n58903 & n59031;
  assign n59033 = ~n59020 & n59032;
  assign n59034 = ~n59021 & n59033;
  assign n59035 = n58900 & ~n59034;
  assign n59036 = ~n59029 & ~n59035;
  assign n59037 = n58980 & n59036;
  assign n59038 = ~P2_P3_FLUSH_REG & ~P2_P3_MORE_REG;
  assign n59039 = n59037 & ~n59038;
  assign n59040 = ~n58935 & n58966;
  assign n59041 = ~n58900 & n59040;
  assign n59042 = n59026 & n59041;
  assign n59043 = ~n59019 & n59042;
  assign n59044 = n58935 & n58966;
  assign n59045 = ~n58900 & n59044;
  assign n59046 = n59026 & n59045;
  assign n59047 = ~n59019 & n59046;
  assign n59048 = n58968 & ~n59019;
  assign n59049 = ~n58935 & ~n58966;
  assign n59050 = n58904 & n59049;
  assign n59051 = ~n59019 & n59050;
  assign n59052 = ~n59043 & ~n59047;
  assign n59053 = ~n59048 & n59052;
  assign n59054 = ~n59051 & n59053;
  assign n59055 = ~n58744 & n58775;
  assign n59056 = ~n58807 & n59055;
  assign n59057 = n58902 & n59056;
  assign n59058 = n59049 & n59057;
  assign n59059 = ~P2_P3_INSTQUEUERD_ADDR_REG_0_ & P2_P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n59060 = ~n58986 & ~n59059;
  assign n59061 = n59011 & n59060;
  assign n59062 = ~n59015 & ~n59061;
  assign n59063 = n59016 & ~n59062;
  assign n59064 = n58997 & ~n59063;
  assign n59065 = n59058 & ~n59064;
  assign n59066 = n59044 & n59057;
  assign n59067 = ~n59064 & n59066;
  assign n59068 = n58902 & n59025;
  assign n59069 = n58967 & n59068;
  assign n59070 = n59001 & ~n59062;
  assign n59071 = n59005 & n59070;
  assign n59072 = n58997 & ~n59071;
  assign n59073 = n59069 & ~n59072;
  assign n59074 = n59049 & n59068;
  assign n59075 = ~n59011 & ~n59060;
  assign n59076 = n59016 & ~n59075;
  assign n59077 = n59015 & n59076;
  assign n59078 = n58997 & ~n59077;
  assign n59079 = n59074 & ~n59078;
  assign n59080 = ~n59065 & ~n59067;
  assign n59081 = ~n59073 & n59080;
  assign n59082 = ~n59079 & n59081;
  assign n59083 = n59054 & n59082;
  assign n59084 = ~n59037 & ~n59083;
  assign n59085 = ~n58935 & ~n59078;
  assign n59086 = n58935 & ~n59072;
  assign n59087 = ~n59085 & ~n59086;
  assign n59088 = ~n58966 & n59068;
  assign n59089 = n59087 & n59088;
  assign n59090 = n58869 & n58900;
  assign n59091 = n58744 & ~n58775;
  assign n59092 = n59090 & n59091;
  assign n59093 = n59044 & n59092;
  assign n59094 = ~n58838 & n59093;
  assign n59095 = n58904 & ~n58966;
  assign n59096 = ~n59042 & ~n59094;
  assign n59097 = ~n59095 & n59096;
  assign n59098 = n58775 & n58869;
  assign n59099 = ~n58807 & n58900;
  assign n59100 = ~n58838 & n59044;
  assign n59101 = n59099 & n59100;
  assign n59102 = n58744 & ~n58900;
  assign n59103 = n58807 & n58838;
  assign n59104 = n59102 & n59103;
  assign n59105 = ~n59101 & ~n59104;
  assign n59106 = n59098 & ~n59105;
  assign n59107 = n59049 & n59103;
  assign n59108 = n59092 & n59107;
  assign n59109 = n58869 & ~n58900;
  assign n59110 = n58838 & n59040;
  assign n59111 = n59025 & n59109;
  assign n59112 = n59110 & n59111;
  assign n59113 = ~n58935 & n59068;
  assign n59114 = ~n59112 & ~n59113;
  assign n59115 = ~n59106 & ~n59108;
  assign n59116 = n59114 & n59115;
  assign n59117 = n58775 & ~n58838;
  assign n59118 = ~n59091 & ~n59117;
  assign n59119 = n58869 & n59118;
  assign n59120 = ~n58900 & ~n59119;
  assign n59121 = ~n58838 & ~n59091;
  assign n59122 = ~n59055 & n59121;
  assign n59123 = ~n58869 & n59122;
  assign n59124 = n58967 & ~n59123;
  assign n59125 = n59024 & n59044;
  assign n59126 = n58744 & n58838;
  assign n59127 = ~n58901 & ~n59126;
  assign n59128 = ~n58935 & n59127;
  assign n59129 = n58775 & n58807;
  assign n59130 = n58966 & n59129;
  assign n59131 = ~n59125 & ~n59128;
  assign n59132 = ~n59130 & n59131;
  assign n59133 = ~n59124 & n59132;
  assign n59134 = n58900 & ~n59133;
  assign n59135 = ~n58869 & ~n59129;
  assign n59136 = n58744 & n59135;
  assign n59137 = n58838 & n58935;
  assign n59138 = n58966 & ~n59137;
  assign n59139 = n58869 & ~n59138;
  assign n59140 = ~n58744 & n59139;
  assign n59141 = ~n58838 & ~n59024;
  assign n59142 = ~n58967 & n59141;
  assign n59143 = ~n58807 & ~n59142;
  assign n59144 = n58775 & ~n58935;
  assign n59145 = n58838 & n59144;
  assign n59146 = n58807 & ~n58935;
  assign n59147 = n59055 & n59146;
  assign n59148 = ~n59024 & n59040;
  assign n59149 = ~n59145 & ~n59147;
  assign n59150 = ~n59148 & n59149;
  assign n59151 = ~n59136 & ~n59140;
  assign n59152 = ~n59143 & n59151;
  assign n59153 = n59150 & n59152;
  assign n59154 = ~n59120 & ~n59134;
  assign n59155 = n59153 & n59154;
  assign n59156 = n59116 & n59155;
  assign n59157 = ~n59093 & n59156;
  assign n59158 = P2_P3_INSTQUEUERD_ADDR_REG_0_ & ~n59157;
  assign n59159 = n59097 & ~n59158;
  assign n59160 = ~P2_P3_INSTQUEUERD_ADDR_REG_2_ & ~n59159;
  assign n59161 = P2_P3_INSTQUEUERD_ADDR_REG_1_ & n59160;
  assign n59162 = P2_P3_INSTQUEUERD_ADDR_REG_2_ & ~n59097;
  assign n59163 = ~P2_P3_INSTQUEUERD_ADDR_REG_1_ & n59162;
  assign n59164 = ~P2_P3_INSTQUEUERD_ADDR_REG_2_ & P2_P3_INSTQUEUERD_ADDR_REG_1_;
  assign n59165 = P2_P3_INSTQUEUERD_ADDR_REG_2_ & ~P2_P3_INSTQUEUERD_ADDR_REG_1_;
  assign n59166 = ~n59164 & ~n59165;
  assign n59167 = n59046 & ~n59166;
  assign n59168 = P2_P3_INSTQUEUERD_ADDR_REG_2_ & ~n58687;
  assign n59169 = ~n58688 & ~n59168;
  assign n59170 = ~n59044 & ~n59049;
  assign n59171 = n59169 & ~n59170;
  assign n59172 = n59057 & n59171;
  assign n59173 = ~n59167 & ~n59172;
  assign n59174 = n58935 & n59098;
  assign n59175 = ~n59099 & ~n59104;
  assign n59176 = n59174 & ~n59175;
  assign n59177 = n59103 & ~n59170;
  assign n59178 = n59092 & n59177;
  assign n59179 = ~n59176 & ~n59178;
  assign n59180 = n59114 & n59179;
  assign n59181 = n59155 & n59180;
  assign n59182 = n59168 & ~n59181;
  assign n59183 = n59173 & ~n59182;
  assign n59184 = ~n59161 & ~n59163;
  assign n59185 = n59183 & n59184;
  assign n59186 = n58807 & n58966;
  assign n59187 = ~n58869 & ~n59040;
  assign n59188 = n59121 & ~n59186;
  assign n59189 = n59187 & n59188;
  assign n59190 = ~n59147 & n59189;
  assign n59191 = n58900 & ~n59190;
  assign n59192 = ~n58900 & ~n59027;
  assign n59193 = n58967 & ~n59122;
  assign n59194 = ~n59191 & ~n59192;
  assign n59195 = ~n59193 & n59194;
  assign n59196 = n59064 & n59066;
  assign n59197 = n59019 & n59046;
  assign n59198 = n59019 & n59050;
  assign n59199 = ~n59197 & ~n59198;
  assign n59200 = ~n58594 & ~n59199;
  assign n59201 = ~n59196 & ~n59200;
  assign n59202 = n59058 & n59064;
  assign n59203 = ~n59055 & n59099;
  assign n59204 = ~n59202 & ~n59203;
  assign n59205 = n59019 & n59042;
  assign n59206 = n58968 & n59019;
  assign n59207 = ~n59205 & ~n59206;
  assign n59208 = n58971 & ~n59207;
  assign n59209 = n59204 & ~n59208;
  assign n59210 = n59195 & n59201;
  assign n59211 = n59209 & n59210;
  assign n59212 = ~n59185 & ~n59211;
  assign n59213 = P2_P3_INSTQUEUERD_ADDR_REG_2_ & n59211;
  assign n59214 = ~n59212 & ~n59213;
  assign n59215 = P2_P3_INSTQUEUERD_ADDR_REG_1_ & n58717;
  assign n59216 = ~n59159 & n59215;
  assign n59217 = P2_P3_INSTQUEUERD_ADDR_REG_2_ & n58687;
  assign n59218 = P2_P3_INSTQUEUERD_ADDR_REG_3_ & ~n59217;
  assign n59219 = ~n59180 & n59218;
  assign n59220 = P2_P3_INSTQUEUERD_ADDR_REG_2_ & P2_P3_INSTQUEUERD_ADDR_REG_1_;
  assign n59221 = ~P2_P3_INSTQUEUERD_ADDR_REG_3_ & n59220;
  assign n59222 = P2_P3_INSTQUEUERD_ADDR_REG_3_ & ~n59220;
  assign n59223 = ~n59221 & ~n59222;
  assign n59224 = n59046 & ~n59223;
  assign n59225 = ~n59219 & ~n59224;
  assign n59226 = ~n58807 & n59094;
  assign n59227 = n58807 & n59094;
  assign n59228 = ~n58968 & ~n59050;
  assign n59229 = ~n59042 & n59228;
  assign n59230 = ~n59226 & ~n59227;
  assign n59231 = n59229 & n59230;
  assign n59232 = n59155 & n59231;
  assign n59233 = n59222 & ~n59232;
  assign n59234 = P2_P3_INSTQUEUERD_ADDR_REG_3_ & ~P2_P3_INSTQUEUERD_ADDR_REG_0_;
  assign n59235 = ~n59155 & n59234;
  assign n59236 = ~n58687 & n58731;
  assign n59237 = ~P2_P3_INSTQUEUERD_ADDR_REG_2_ & ~n58687;
  assign n59238 = P2_P3_INSTQUEUERD_ADDR_REG_3_ & ~n59237;
  assign n59239 = ~n59236 & ~n59238;
  assign n59240 = ~n59170 & n59239;
  assign n59241 = n59057 & n59240;
  assign n59242 = ~n59235 & ~n59241;
  assign n59243 = n59225 & ~n59233;
  assign n59244 = n59242 & n59243;
  assign n59245 = ~n59216 & n59244;
  assign n59246 = ~n59211 & ~n59245;
  assign n59247 = P2_P3_INSTQUEUERD_ADDR_REG_3_ & n59211;
  assign n59248 = ~n59246 & ~n59247;
  assign n59249 = ~n59214 & ~n59248;
  assign n59250 = P2_P3_INSTQUEUERD_ADDR_REG_4_ & n59211;
  assign n59251 = P2_P3_INSTQUEUERD_ADDR_REG_3_ & n59220;
  assign n59252 = ~P2_P3_INSTQUEUERD_ADDR_REG_4_ & n59251;
  assign n59253 = P2_P3_INSTQUEUERD_ADDR_REG_4_ & ~n59251;
  assign n59254 = ~n59252 & ~n59253;
  assign n59255 = n59046 & ~n59254;
  assign n59256 = ~n59211 & n59255;
  assign n59257 = ~n59250 & ~n59256;
  assign n59258 = ~n59249 & n59257;
  assign n59259 = ~P2_P3_INSTQUEUEWR_ADDR_REG_3_ & ~n59248;
  assign n59260 = ~P2_P3_INSTQUEUEWR_ADDR_REG_4_ & ~n59257;
  assign n59261 = P2_P3_INSTQUEUEWR_ADDR_REG_2_ & n59214;
  assign n59262 = P2_P3_INSTQUEUEWR_ADDR_REG_3_ & n59248;
  assign n59263 = n59055 & n59101;
  assign n59264 = ~n59058 & ~n59263;
  assign n59265 = n59093 & n59103;
  assign n59266 = n59156 & ~n59265;
  assign n59267 = n59264 & n59266;
  assign n59268 = ~P2_P3_INSTQUEUERD_ADDR_REG_0_ & ~n59267;
  assign n59269 = P2_P3_INSTQUEUERD_ADDR_REG_0_ & ~n59097;
  assign n59270 = P2_P3_INSTQUEUERD_ADDR_REG_0_ & n59046;
  assign n59271 = ~n59268 & ~n59269;
  assign n59272 = ~n59270 & n59271;
  assign n59273 = ~n59211 & ~n59272;
  assign n59274 = P2_P3_INSTQUEUERD_ADDR_REG_0_ & n59211;
  assign n59275 = ~n59273 & ~n59274;
  assign n59276 = P2_P3_INSTQUEUEWR_ADDR_REG_0_ & n59275;
  assign n59277 = ~P2_P3_INSTQUEUEWR_ADDR_REG_1_ & ~n59276;
  assign n59278 = ~P2_P3_INSTQUEUEWR_ADDR_REG_2_ & ~n59214;
  assign n59279 = ~P2_P3_INSTQUEUERD_ADDR_REG_1_ & ~n59159;
  assign n59280 = ~P2_P3_INSTQUEUERD_ADDR_REG_1_ & n59046;
  assign n59281 = ~n58687 & ~n58700;
  assign n59282 = ~n59264 & n59281;
  assign n59283 = ~n59280 & ~n59282;
  assign n59284 = n58691 & ~n59266;
  assign n59285 = n59283 & ~n59284;
  assign n59286 = ~n59279 & n59285;
  assign n59287 = ~n59211 & ~n59286;
  assign n59288 = P2_P3_INSTQUEUERD_ADDR_REG_1_ & n59211;
  assign n59289 = ~n59287 & ~n59288;
  assign n59290 = P2_P3_INSTQUEUEWR_ADDR_REG_1_ & n59276;
  assign n59291 = ~n59289 & ~n59290;
  assign n59292 = ~n59277 & ~n59278;
  assign n59293 = ~n59291 & n59292;
  assign n59294 = ~n59261 & ~n59262;
  assign n59295 = ~n59293 & n59294;
  assign n59296 = ~n59259 & ~n59260;
  assign n59297 = ~n59295 & n59296;
  assign n59298 = P2_P3_INSTQUEUEWR_ADDR_REG_4_ & n59257;
  assign n59299 = ~n59297 & ~n59298;
  assign n59300 = ~n59039 & ~n59084;
  assign n59301 = ~n59089 & n59300;
  assign n59302 = n59258 & n59301;
  assign n59303 = ~n59299 & n59302;
  assign n59304 = n58970 & n59303;
  assign n59305 = P2_P3_STATE2_REG_0_ & ~n59304;
  assign n59306 = ~n58681 & ~n59305;
  assign n59307 = P2_P3_STATE2_REG_2_ & n59306;
  assign n59308 = P2_P3_STATE2_REG_0_ & ~n59307;
  assign n59309 = n58679 & n59308;
  assign n59310 = P2_P3_STATE2_REG_3_ & ~n59308;
  assign n10331 = n59309 | n59310;
  assign n59312 = ~P2_P3_STATE2_REG_2_ & ~n58594;
  assign n59313 = P2_P3_STATE2_REG_0_ & ~n59312;
  assign n59314 = ~P2_P3_STATE2_REG_0_ & ~P2_P3_STATEBS16_REG;
  assign n59315 = ~n59313 & ~n59314;
  assign n59316 = P2_P3_STATE2_REG_1_ & n59315;
  assign n59317 = P2_P3_STATE2_REG_2_ & ~P2_P3_STATE2_REG_1_;
  assign n59318 = ~n59316 & ~n59317;
  assign n59319 = P2_P3_STATE2_REG_2_ & ~n59308;
  assign n10336 = ~n59318 | n59319;
  assign n59321 = P2_P3_STATE2_REG_0_ & n59317;
  assign n59322 = ~n59307 & n59321;
  assign n59323 = ~P2_P3_STATE2_REG_2_ & P2_P3_STATE2_REG_0_;
  assign n59324 = n58594 & n59323;
  assign n59325 = ~n59307 & ~n59324;
  assign n59326 = P2_P3_STATE2_REG_1_ & ~n59325;
  assign n59327 = ~P2_P3_STATE2_REG_3_ & ~P2_P3_STATE2_REG_1_;
  assign n59328 = ~n58594 & n59327;
  assign n59329 = n59308 & n59328;
  assign n59330 = P2_P3_STATE2_REG_1_ & ~P2_P3_STATE2_REG_0_;
  assign n59331 = ~P2_P3_STATE2_REG_2_ & n59330;
  assign n59332 = ~P2_P3_STATEBS16_REG & n59331;
  assign n59333 = ~n59322 & ~n59326;
  assign n59334 = ~n59329 & n59333;
  assign n10341 = n59332 | ~n59334;
  assign n59336 = P2_P3_STATE2_REG_3_ & ~P2_P3_INSTQUEUERD_ADDR_REG_4_;
  assign n59337 = ~P2_P3_STATE2_REG_2_ & ~P2_P3_STATE2_REG_1_;
  assign n59338 = n59336 & n59337;
  assign n59339 = ~n59307 & ~n59338;
  assign n59340 = ~P2_P3_STATE2_REG_0_ & n59339;
  assign n59341 = P2_P3_INSTADDRPOINTER_REG_0_ & P2_P3_INSTADDRPOINTER_REG_31_;
  assign n59342 = P2_P3_INSTADDRPOINTER_REG_0_ & ~P2_P3_INSTADDRPOINTER_REG_31_;
  assign n59343 = ~n59341 & ~n59342;
  assign n59344 = P2_P3_FLUSH_REG & n59343;
  assign n59345 = P2_P3_INSTQUEUERD_ADDR_REG_0_ & ~P2_P3_FLUSH_REG;
  assign n59346 = ~n59344 & ~n59345;
  assign n59347 = P2_P3_INSTADDRPOINTER_REG_0_ & ~P2_P3_INSTADDRPOINTER_REG_1_;
  assign n59348 = ~P2_P3_INSTADDRPOINTER_REG_0_ & P2_P3_INSTADDRPOINTER_REG_1_;
  assign n59349 = ~n59347 & ~n59348;
  assign n59350 = P2_P3_INSTADDRPOINTER_REG_31_ & ~n59349;
  assign n59351 = P2_P3_INSTADDRPOINTER_REG_1_ & ~P2_P3_INSTADDRPOINTER_REG_31_;
  assign n59352 = ~n59350 & ~n59351;
  assign n59353 = ~n59343 & n59352;
  assign n59354 = P2_P3_FLUSH_REG & n59353;
  assign n59355 = P2_P3_INSTQUEUERD_ADDR_REG_1_ & ~P2_P3_FLUSH_REG;
  assign n59356 = ~n59354 & ~n59355;
  assign n59357 = n59346 & n59356;
  assign n59358 = P2_P3_INSTQUEUERD_ADDR_REG_3_ & ~P2_P3_FLUSH_REG;
  assign n59359 = ~n59343 & ~n59352;
  assign n59360 = P2_P3_FLUSH_REG & n59359;
  assign n59361 = P2_P3_INSTQUEUERD_ADDR_REG_2_ & ~P2_P3_FLUSH_REG;
  assign n59362 = ~n59360 & ~n59361;
  assign n59363 = ~n59357 & n59358;
  assign n59364 = ~n59362 & n59363;
  assign n59365 = P2_P3_INSTQUEUERD_ADDR_REG_4_ & ~P2_P3_FLUSH_REG;
  assign n59366 = ~n59364 & ~n59365;
  assign n59367 = n58679 & n59366;
  assign n59368 = ~n59307 & ~n59367;
  assign n59369 = P2_P3_STATE2_REG_0_ & ~n59368;
  assign n59370 = P2_P3_STATE2_REG_3_ & P2_P3_STATE2_REG_0_;
  assign n59371 = n59337 & n59370;
  assign n59372 = ~n59324 & ~n59371;
  assign n59373 = ~n59303 & n59321;
  assign n59374 = n59372 & ~n59373;
  assign n59375 = ~n59340 & ~n59369;
  assign n10346 = ~n59374 | ~n59375;
  assign n59377 = P2_P3_INSTQUEUEWR_ADDR_REG_1_ & P2_P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n59378 = P2_P3_INSTQUEUEWR_ADDR_REG_2_ & n59377;
  assign n59379 = P2_P3_INSTQUEUEWR_ADDR_REG_3_ & n59378;
  assign n59380 = P2_P3_STATE2_REG_3_ & ~n59379;
  assign n59381 = ~P2_P3_STATE2_REG_2_ & P2_P3_STATE2_REG_1_;
  assign n59382 = ~n59317 & ~n59381;
  assign n59383 = ~n59336 & n59382;
  assign n59384 = ~P2_P3_STATE2_REG_0_ & ~n59383;
  assign n59385 = ~n59380 & n59384;
  assign n59386 = ~P2_P3_INSTQUEUEWR_ADDR_REG_2_ & n59377;
  assign n59387 = P2_P3_INSTQUEUEWR_ADDR_REG_2_ & ~n59377;
  assign n59388 = ~n59386 & ~n59387;
  assign n59389 = ~P2_P3_INSTQUEUEWR_ADDR_REG_3_ & n59378;
  assign n59390 = P2_P3_INSTQUEUEWR_ADDR_REG_3_ & ~n59378;
  assign n59391 = ~n59389 & ~n59390;
  assign n59392 = ~n59388 & ~n59391;
  assign n59393 = ~P2_P3_INSTQUEUEWR_ADDR_REG_1_ & P2_P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n59394 = P2_P3_INSTQUEUEWR_ADDR_REG_1_ & ~P2_P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n59395 = ~n59393 & ~n59394;
  assign n59396 = ~P2_P3_INSTQUEUEWR_ADDR_REG_0_ & ~n59395;
  assign n59397 = n59392 & n59396;
  assign n59398 = ~n59379 & ~n59397;
  assign n59399 = ~P2_P3_STATE2_REG_3_ & ~P2_P3_STATE2_REG_2_;
  assign n59400 = ~P2_P3_STATEBS16_REG & n59399;
  assign n59401 = ~P2_P3_STATE2_REG_2_ & ~n59400;
  assign n59402 = P2_P3_INSTQUEUEWR_ADDR_REG_0_ & ~n59395;
  assign n59403 = ~P2_P3_INSTQUEUEWR_ADDR_REG_0_ & n59395;
  assign n59404 = ~n59402 & ~n59403;
  assign n59405 = ~P2_P3_INSTQUEUEWR_ADDR_REG_0_ & ~n59404;
  assign n59406 = P2_P3_INSTQUEUEWR_ADDR_REG_0_ & n59404;
  assign n59407 = ~n59405 & ~n59406;
  assign n59408 = ~P2_P3_INSTQUEUEWR_ADDR_REG_0_ & ~n59407;
  assign n59409 = ~n59388 & ~n59396;
  assign n59410 = n59388 & n59396;
  assign n59411 = ~n59409 & ~n59410;
  assign n59412 = P2_P3_INSTQUEUEWR_ADDR_REG_0_ & ~n59404;
  assign n59413 = ~n59411 & ~n59412;
  assign n59414 = n59411 & n59412;
  assign n59415 = ~n59413 & ~n59414;
  assign n59416 = ~n59388 & n59391;
  assign n59417 = n59396 & n59416;
  assign n59418 = ~n59388 & n59396;
  assign n59419 = ~n59391 & ~n59418;
  assign n59420 = ~n59417 & ~n59419;
  assign n59421 = n59411 & ~n59420;
  assign n59422 = ~n59412 & ~n59420;
  assign n59423 = ~n59421 & ~n59422;
  assign n59424 = ~n59411 & n59420;
  assign n59425 = n59412 & n59424;
  assign n59426 = n59423 & ~n59425;
  assign n59427 = ~n59415 & ~n59426;
  assign n59428 = n59408 & n59427;
  assign n59429 = ~n59411 & ~n59420;
  assign n59430 = n59412 & n59429;
  assign n59431 = ~n59428 & ~n59430;
  assign n59432 = n59401 & ~n59431;
  assign n59433 = n59398 & ~n59432;
  assign n59434 = n59385 & ~n59433;
  assign n59435 = P2_P3_INSTQUEUE_REG_15__7_ & ~n59434;
  assign n59436 = P2_P3_STATEBS16_REG & n59399;
  assign n59437 = n59384 & n59436;
  assign n59438 = P2_BUF2_REG_23_ & n59437;
  assign n59439 = n59430 & n59438;
  assign n59440 = P2_P3_STATE2_REG_3_ & n59384;
  assign n59441 = ~n58838 & n59440;
  assign n59442 = n59379 & n59441;
  assign n59443 = ~n59439 & ~n59442;
  assign n59444 = P2_BUF2_REG_31_ & n59437;
  assign n59445 = n59428 & n59444;
  assign n59446 = n59443 & ~n59445;
  assign n59447 = n59431 & n59436;
  assign n59448 = n59401 & ~n59447;
  assign n59449 = ~n59398 & ~n59448;
  assign n59450 = P2_BUF2_REG_7_ & n59384;
  assign n59451 = n59449 & n59450;
  assign n59452 = ~n59435 & n59446;
  assign n10351 = n59451 | ~n59452;
  assign n59454 = P2_P3_INSTQUEUE_REG_15__6_ & ~n59434;
  assign n59455 = P2_BUF2_REG_22_ & n59437;
  assign n59456 = n59430 & n59455;
  assign n59457 = ~n58775 & n59440;
  assign n59458 = n59379 & n59457;
  assign n59459 = ~n59456 & ~n59458;
  assign n59460 = P2_BUF2_REG_30_ & n59437;
  assign n59461 = n59428 & n59460;
  assign n59462 = n59459 & ~n59461;
  assign n59463 = P2_BUF2_REG_6_ & n59384;
  assign n59464 = n59449 & n59463;
  assign n59465 = ~n59454 & n59462;
  assign n10356 = n59464 | ~n59465;
  assign n59467 = P2_P3_INSTQUEUE_REG_15__5_ & ~n59434;
  assign n59468 = P2_BUF2_REG_21_ & n59437;
  assign n59469 = n59430 & n59468;
  assign n59470 = ~n58744 & n59440;
  assign n59471 = n59379 & n59470;
  assign n59472 = ~n59469 & ~n59471;
  assign n59473 = P2_BUF2_REG_29_ & n59437;
  assign n59474 = n59428 & n59473;
  assign n59475 = n59472 & ~n59474;
  assign n59476 = P2_BUF2_REG_5_ & n59384;
  assign n59477 = n59449 & n59476;
  assign n59478 = ~n59467 & n59475;
  assign n10361 = n59477 | ~n59478;
  assign n59480 = P2_P3_INSTQUEUE_REG_15__4_ & ~n59434;
  assign n59481 = P2_BUF2_REG_20_ & n59437;
  assign n59482 = n59430 & n59481;
  assign n59483 = ~n58807 & n59440;
  assign n59484 = n59379 & n59483;
  assign n59485 = ~n59482 & ~n59484;
  assign n59486 = P2_BUF2_REG_28_ & n59437;
  assign n59487 = n59428 & n59486;
  assign n59488 = n59485 & ~n59487;
  assign n59489 = P2_BUF2_REG_4_ & n59384;
  assign n59490 = n59449 & n59489;
  assign n59491 = ~n59480 & n59488;
  assign n10366 = n59490 | ~n59491;
  assign n59493 = P2_P3_INSTQUEUE_REG_15__3_ & ~n59434;
  assign n59494 = P2_BUF2_REG_19_ & n59437;
  assign n59495 = n59430 & n59494;
  assign n59496 = ~n58869 & n59440;
  assign n59497 = n59379 & n59496;
  assign n59498 = ~n59495 & ~n59497;
  assign n59499 = P2_BUF2_REG_27_ & n59437;
  assign n59500 = n59428 & n59499;
  assign n59501 = n59498 & ~n59500;
  assign n59502 = P2_BUF2_REG_3_ & n59384;
  assign n59503 = n59449 & n59502;
  assign n59504 = ~n59493 & n59501;
  assign n10371 = n59503 | ~n59504;
  assign n59506 = P2_P3_INSTQUEUE_REG_15__2_ & ~n59434;
  assign n59507 = P2_BUF2_REG_18_ & n59437;
  assign n59508 = n59430 & n59507;
  assign n59509 = ~n58900 & n59440;
  assign n59510 = n59379 & n59509;
  assign n59511 = ~n59508 & ~n59510;
  assign n59512 = P2_BUF2_REG_26_ & n59437;
  assign n59513 = n59428 & n59512;
  assign n59514 = n59511 & ~n59513;
  assign n59515 = P2_BUF2_REG_2_ & n59384;
  assign n59516 = n59449 & n59515;
  assign n59517 = ~n59506 & n59514;
  assign n10376 = n59516 | ~n59517;
  assign n59519 = P2_P3_INSTQUEUE_REG_15__1_ & ~n59434;
  assign n59520 = P2_BUF2_REG_17_ & n59437;
  assign n59521 = n59430 & n59520;
  assign n59522 = ~n58935 & n59440;
  assign n59523 = n59379 & n59522;
  assign n59524 = ~n59521 & ~n59523;
  assign n59525 = P2_BUF2_REG_25_ & n59437;
  assign n59526 = n59428 & n59525;
  assign n59527 = n59524 & ~n59526;
  assign n59528 = P2_BUF2_REG_1_ & n59384;
  assign n59529 = n59449 & n59528;
  assign n59530 = ~n59519 & n59527;
  assign n10381 = n59529 | ~n59530;
  assign n59532 = P2_P3_INSTQUEUE_REG_15__0_ & ~n59434;
  assign n59533 = P2_BUF2_REG_16_ & n59437;
  assign n59534 = n59430 & n59533;
  assign n59535 = ~n58966 & n59440;
  assign n59536 = n59379 & n59535;
  assign n59537 = ~n59534 & ~n59536;
  assign n59538 = P2_BUF2_REG_24_ & n59437;
  assign n59539 = n59428 & n59538;
  assign n59540 = n59537 & ~n59539;
  assign n59541 = P2_BUF2_REG_0_ & n59384;
  assign n59542 = n59449 & n59541;
  assign n59543 = ~n59532 & n59540;
  assign n10386 = n59542 | ~n59543;
  assign n59545 = P2_P3_INSTQUEUEWR_ADDR_REG_3_ & P2_P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n59546 = P2_P3_INSTQUEUEWR_ADDR_REG_2_ & ~P2_P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n59547 = n59545 & n59546;
  assign n59548 = P2_P3_STATE2_REG_3_ & ~n59547;
  assign n59549 = n59384 & ~n59548;
  assign n59550 = n59392 & n59402;
  assign n59551 = ~n59547 & ~n59550;
  assign n59552 = P2_P3_INSTQUEUEWR_ADDR_REG_0_ & ~n59407;
  assign n59553 = n59427 & n59552;
  assign n59554 = n59405 & n59429;
  assign n59555 = ~n59553 & ~n59554;
  assign n59556 = n59401 & ~n59555;
  assign n59557 = n59551 & ~n59556;
  assign n59558 = n59549 & ~n59557;
  assign n59559 = P2_P3_INSTQUEUE_REG_14__7_ & ~n59558;
  assign n59560 = n59438 & n59554;
  assign n59561 = n59441 & n59547;
  assign n59562 = ~n59560 & ~n59561;
  assign n59563 = n59444 & n59553;
  assign n59564 = n59562 & ~n59563;
  assign n59565 = n59436 & n59555;
  assign n59566 = n59401 & ~n59565;
  assign n59567 = ~n59551 & ~n59566;
  assign n59568 = n59450 & n59567;
  assign n59569 = ~n59559 & n59564;
  assign n10391 = n59568 | ~n59569;
  assign n59571 = P2_P3_INSTQUEUE_REG_14__6_ & ~n59558;
  assign n59572 = n59455 & n59554;
  assign n59573 = n59457 & n59547;
  assign n59574 = ~n59572 & ~n59573;
  assign n59575 = n59460 & n59553;
  assign n59576 = n59574 & ~n59575;
  assign n59577 = n59463 & n59567;
  assign n59578 = ~n59571 & n59576;
  assign n10396 = n59577 | ~n59578;
  assign n59580 = P2_P3_INSTQUEUE_REG_14__5_ & ~n59558;
  assign n59581 = n59468 & n59554;
  assign n59582 = n59470 & n59547;
  assign n59583 = ~n59581 & ~n59582;
  assign n59584 = n59473 & n59553;
  assign n59585 = n59583 & ~n59584;
  assign n59586 = n59476 & n59567;
  assign n59587 = ~n59580 & n59585;
  assign n10401 = n59586 | ~n59587;
  assign n59589 = P2_P3_INSTQUEUE_REG_14__4_ & ~n59558;
  assign n59590 = n59481 & n59554;
  assign n59591 = n59483 & n59547;
  assign n59592 = ~n59590 & ~n59591;
  assign n59593 = n59486 & n59553;
  assign n59594 = n59592 & ~n59593;
  assign n59595 = n59489 & n59567;
  assign n59596 = ~n59589 & n59594;
  assign n10406 = n59595 | ~n59596;
  assign n59598 = P2_P3_INSTQUEUE_REG_14__3_ & ~n59558;
  assign n59599 = n59494 & n59554;
  assign n59600 = n59496 & n59547;
  assign n59601 = ~n59599 & ~n59600;
  assign n59602 = n59499 & n59553;
  assign n59603 = n59601 & ~n59602;
  assign n59604 = n59502 & n59567;
  assign n59605 = ~n59598 & n59603;
  assign n10411 = n59604 | ~n59605;
  assign n59607 = P2_P3_INSTQUEUE_REG_14__2_ & ~n59558;
  assign n59608 = n59507 & n59554;
  assign n59609 = n59509 & n59547;
  assign n59610 = ~n59608 & ~n59609;
  assign n59611 = n59512 & n59553;
  assign n59612 = n59610 & ~n59611;
  assign n59613 = n59515 & n59567;
  assign n59614 = ~n59607 & n59612;
  assign n10416 = n59613 | ~n59614;
  assign n59616 = P2_P3_INSTQUEUE_REG_14__1_ & ~n59558;
  assign n59617 = n59520 & n59554;
  assign n59618 = n59522 & n59547;
  assign n59619 = ~n59617 & ~n59618;
  assign n59620 = n59525 & n59553;
  assign n59621 = n59619 & ~n59620;
  assign n59622 = n59528 & n59567;
  assign n59623 = ~n59616 & n59621;
  assign n10421 = n59622 | ~n59623;
  assign n59625 = P2_P3_INSTQUEUE_REG_14__0_ & ~n59558;
  assign n59626 = n59533 & n59554;
  assign n59627 = n59535 & n59547;
  assign n59628 = ~n59626 & ~n59627;
  assign n59629 = n59538 & n59553;
  assign n59630 = n59628 & ~n59629;
  assign n59631 = n59541 & n59567;
  assign n59632 = ~n59625 & n59630;
  assign n10426 = n59631 | ~n59632;
  assign n59634 = P2_P3_INSTQUEUEWR_ADDR_REG_3_ & P2_P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n59635 = n59393 & n59634;
  assign n59636 = P2_P3_STATE2_REG_3_ & ~n59635;
  assign n59637 = n59384 & ~n59636;
  assign n59638 = n59392 & n59403;
  assign n59639 = ~n59635 & ~n59638;
  assign n59640 = ~P2_P3_INSTQUEUEWR_ADDR_REG_0_ & n59407;
  assign n59641 = n59427 & n59640;
  assign n59642 = n59406 & n59429;
  assign n59643 = ~n59641 & ~n59642;
  assign n59644 = n59401 & ~n59643;
  assign n59645 = n59639 & ~n59644;
  assign n59646 = n59637 & ~n59645;
  assign n59647 = P2_P3_INSTQUEUE_REG_13__7_ & ~n59646;
  assign n59648 = n59438 & n59642;
  assign n59649 = n59441 & n59635;
  assign n59650 = ~n59648 & ~n59649;
  assign n59651 = n59444 & n59641;
  assign n59652 = n59650 & ~n59651;
  assign n59653 = n59436 & n59643;
  assign n59654 = n59401 & ~n59653;
  assign n59655 = ~n59639 & ~n59654;
  assign n59656 = n59450 & n59655;
  assign n59657 = ~n59647 & n59652;
  assign n10431 = n59656 | ~n59657;
  assign n59659 = P2_P3_INSTQUEUE_REG_13__6_ & ~n59646;
  assign n59660 = n59455 & n59642;
  assign n59661 = n59457 & n59635;
  assign n59662 = ~n59660 & ~n59661;
  assign n59663 = n59460 & n59641;
  assign n59664 = n59662 & ~n59663;
  assign n59665 = n59463 & n59655;
  assign n59666 = ~n59659 & n59664;
  assign n10436 = n59665 | ~n59666;
  assign n59668 = P2_P3_INSTQUEUE_REG_13__5_ & ~n59646;
  assign n59669 = n59468 & n59642;
  assign n59670 = n59470 & n59635;
  assign n59671 = ~n59669 & ~n59670;
  assign n59672 = n59473 & n59641;
  assign n59673 = n59671 & ~n59672;
  assign n59674 = n59476 & n59655;
  assign n59675 = ~n59668 & n59673;
  assign n10441 = n59674 | ~n59675;
  assign n59677 = P2_P3_INSTQUEUE_REG_13__4_ & ~n59646;
  assign n59678 = n59481 & n59642;
  assign n59679 = n59483 & n59635;
  assign n59680 = ~n59678 & ~n59679;
  assign n59681 = n59486 & n59641;
  assign n59682 = n59680 & ~n59681;
  assign n59683 = n59489 & n59655;
  assign n59684 = ~n59677 & n59682;
  assign n10446 = n59683 | ~n59684;
  assign n59686 = P2_P3_INSTQUEUE_REG_13__3_ & ~n59646;
  assign n59687 = n59494 & n59642;
  assign n59688 = n59496 & n59635;
  assign n59689 = ~n59687 & ~n59688;
  assign n59690 = n59499 & n59641;
  assign n59691 = n59689 & ~n59690;
  assign n59692 = n59502 & n59655;
  assign n59693 = ~n59686 & n59691;
  assign n10451 = n59692 | ~n59693;
  assign n59695 = P2_P3_INSTQUEUE_REG_13__2_ & ~n59646;
  assign n59696 = n59507 & n59642;
  assign n59697 = n59509 & n59635;
  assign n59698 = ~n59696 & ~n59697;
  assign n59699 = n59512 & n59641;
  assign n59700 = n59698 & ~n59699;
  assign n59701 = n59515 & n59655;
  assign n59702 = ~n59695 & n59700;
  assign n10456 = n59701 | ~n59702;
  assign n59704 = P2_P3_INSTQUEUE_REG_13__1_ & ~n59646;
  assign n59705 = n59520 & n59642;
  assign n59706 = n59522 & n59635;
  assign n59707 = ~n59705 & ~n59706;
  assign n59708 = n59525 & n59641;
  assign n59709 = n59707 & ~n59708;
  assign n59710 = n59528 & n59655;
  assign n59711 = ~n59704 & n59709;
  assign n10461 = n59710 | ~n59711;
  assign n59713 = P2_P3_INSTQUEUE_REG_13__0_ & ~n59646;
  assign n59714 = n59533 & n59642;
  assign n59715 = n59535 & n59635;
  assign n59716 = ~n59714 & ~n59715;
  assign n59717 = n59538 & n59641;
  assign n59718 = n59716 & ~n59717;
  assign n59719 = n59541 & n59655;
  assign n59720 = ~n59713 & n59718;
  assign n10466 = n59719 | ~n59720;
  assign n59722 = P2_P3_INSTQUEUEWR_ADDR_REG_3_ & ~P2_P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n59723 = n59546 & n59722;
  assign n59724 = P2_P3_STATE2_REG_3_ & ~n59723;
  assign n59725 = n59384 & ~n59724;
  assign n59726 = P2_P3_INSTQUEUEWR_ADDR_REG_0_ & n59407;
  assign n59727 = n59427 & n59726;
  assign n59728 = ~P2_P3_INSTQUEUEWR_ADDR_REG_0_ & n59404;
  assign n59729 = n59429 & n59728;
  assign n59730 = ~n59727 & ~n59729;
  assign n59731 = n59401 & ~n59730;
  assign n59732 = n59392 & n59395;
  assign n59733 = ~n59731 & ~n59732;
  assign n59734 = n59725 & ~n59733;
  assign n59735 = P2_P3_INSTQUEUE_REG_12__7_ & ~n59734;
  assign n59736 = n59438 & n59729;
  assign n59737 = n59441 & n59723;
  assign n59738 = ~n59736 & ~n59737;
  assign n59739 = n59444 & n59727;
  assign n59740 = n59738 & ~n59739;
  assign n59741 = n59436 & n59730;
  assign n59742 = n59401 & ~n59741;
  assign n59743 = n59732 & ~n59742;
  assign n59744 = n59450 & n59743;
  assign n59745 = ~n59735 & n59740;
  assign n10471 = n59744 | ~n59745;
  assign n59747 = P2_P3_INSTQUEUE_REG_12__6_ & ~n59734;
  assign n59748 = n59455 & n59729;
  assign n59749 = n59457 & n59723;
  assign n59750 = ~n59748 & ~n59749;
  assign n59751 = n59460 & n59727;
  assign n59752 = n59750 & ~n59751;
  assign n59753 = n59463 & n59743;
  assign n59754 = ~n59747 & n59752;
  assign n10476 = n59753 | ~n59754;
  assign n59756 = P2_P3_INSTQUEUE_REG_12__5_ & ~n59734;
  assign n59757 = n59468 & n59729;
  assign n59758 = n59470 & n59723;
  assign n59759 = ~n59757 & ~n59758;
  assign n59760 = n59473 & n59727;
  assign n59761 = n59759 & ~n59760;
  assign n59762 = n59476 & n59743;
  assign n59763 = ~n59756 & n59761;
  assign n10481 = n59762 | ~n59763;
  assign n59765 = P2_P3_INSTQUEUE_REG_12__4_ & ~n59734;
  assign n59766 = n59481 & n59729;
  assign n59767 = n59483 & n59723;
  assign n59768 = ~n59766 & ~n59767;
  assign n59769 = n59486 & n59727;
  assign n59770 = n59768 & ~n59769;
  assign n59771 = n59489 & n59743;
  assign n59772 = ~n59765 & n59770;
  assign n10486 = n59771 | ~n59772;
  assign n59774 = P2_P3_INSTQUEUE_REG_12__3_ & ~n59734;
  assign n59775 = n59494 & n59729;
  assign n59776 = n59496 & n59723;
  assign n59777 = ~n59775 & ~n59776;
  assign n59778 = n59499 & n59727;
  assign n59779 = n59777 & ~n59778;
  assign n59780 = n59502 & n59743;
  assign n59781 = ~n59774 & n59779;
  assign n10491 = n59780 | ~n59781;
  assign n59783 = P2_P3_INSTQUEUE_REG_12__2_ & ~n59734;
  assign n59784 = n59507 & n59729;
  assign n59785 = n59509 & n59723;
  assign n59786 = ~n59784 & ~n59785;
  assign n59787 = n59512 & n59727;
  assign n59788 = n59786 & ~n59787;
  assign n59789 = n59515 & n59743;
  assign n59790 = ~n59783 & n59788;
  assign n10496 = n59789 | ~n59790;
  assign n59792 = P2_P3_INSTQUEUE_REG_12__1_ & ~n59734;
  assign n59793 = n59520 & n59729;
  assign n59794 = n59522 & n59723;
  assign n59795 = ~n59793 & ~n59794;
  assign n59796 = n59525 & n59727;
  assign n59797 = n59795 & ~n59796;
  assign n59798 = n59528 & n59743;
  assign n59799 = ~n59792 & n59797;
  assign n10501 = n59798 | ~n59799;
  assign n59801 = P2_P3_INSTQUEUE_REG_12__0_ & ~n59734;
  assign n59802 = n59533 & n59729;
  assign n59803 = n59535 & n59723;
  assign n59804 = ~n59802 & ~n59803;
  assign n59805 = n59538 & n59727;
  assign n59806 = n59804 & ~n59805;
  assign n59807 = n59541 & n59743;
  assign n59808 = ~n59801 & n59806;
  assign n10506 = n59807 | ~n59808;
  assign n59810 = P2_P3_INSTQUEUEWR_ADDR_REG_3_ & ~P2_P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n59811 = n59377 & n59810;
  assign n59812 = P2_P3_STATE2_REG_3_ & ~n59811;
  assign n59813 = n59384 & ~n59812;
  assign n59814 = n59388 & ~n59391;
  assign n59815 = n59396 & n59814;
  assign n59816 = ~n59811 & ~n59815;
  assign n59817 = n59415 & ~n59426;
  assign n59818 = n59408 & n59817;
  assign n59819 = n59412 & n59421;
  assign n59820 = ~n59818 & ~n59819;
  assign n59821 = n59401 & ~n59820;
  assign n59822 = n59816 & ~n59821;
  assign n59823 = n59813 & ~n59822;
  assign n59824 = P2_P3_INSTQUEUE_REG_11__7_ & ~n59823;
  assign n59825 = n59438 & n59819;
  assign n59826 = n59441 & n59811;
  assign n59827 = ~n59825 & ~n59826;
  assign n59828 = n59444 & n59818;
  assign n59829 = n59827 & ~n59828;
  assign n59830 = n59436 & n59820;
  assign n59831 = n59401 & ~n59830;
  assign n59832 = ~n59816 & ~n59831;
  assign n59833 = n59450 & n59832;
  assign n59834 = ~n59824 & n59829;
  assign n10511 = n59833 | ~n59834;
  assign n59836 = P2_P3_INSTQUEUE_REG_11__6_ & ~n59823;
  assign n59837 = n59455 & n59819;
  assign n59838 = n59457 & n59811;
  assign n59839 = ~n59837 & ~n59838;
  assign n59840 = n59460 & n59818;
  assign n59841 = n59839 & ~n59840;
  assign n59842 = n59463 & n59832;
  assign n59843 = ~n59836 & n59841;
  assign n10516 = n59842 | ~n59843;
  assign n59845 = P2_P3_INSTQUEUE_REG_11__5_ & ~n59823;
  assign n59846 = n59468 & n59819;
  assign n59847 = n59470 & n59811;
  assign n59848 = ~n59846 & ~n59847;
  assign n59849 = n59473 & n59818;
  assign n59850 = n59848 & ~n59849;
  assign n59851 = n59476 & n59832;
  assign n59852 = ~n59845 & n59850;
  assign n10521 = n59851 | ~n59852;
  assign n59854 = P2_P3_INSTQUEUE_REG_11__4_ & ~n59823;
  assign n59855 = n59481 & n59819;
  assign n59856 = n59483 & n59811;
  assign n59857 = ~n59855 & ~n59856;
  assign n59858 = n59486 & n59818;
  assign n59859 = n59857 & ~n59858;
  assign n59860 = n59489 & n59832;
  assign n59861 = ~n59854 & n59859;
  assign n10526 = n59860 | ~n59861;
  assign n59863 = P2_P3_INSTQUEUE_REG_11__3_ & ~n59823;
  assign n59864 = n59494 & n59819;
  assign n59865 = n59496 & n59811;
  assign n59866 = ~n59864 & ~n59865;
  assign n59867 = n59499 & n59818;
  assign n59868 = n59866 & ~n59867;
  assign n59869 = n59502 & n59832;
  assign n59870 = ~n59863 & n59868;
  assign n10531 = n59869 | ~n59870;
  assign n59872 = P2_P3_INSTQUEUE_REG_11__2_ & ~n59823;
  assign n59873 = n59507 & n59819;
  assign n59874 = n59509 & n59811;
  assign n59875 = ~n59873 & ~n59874;
  assign n59876 = n59512 & n59818;
  assign n59877 = n59875 & ~n59876;
  assign n59878 = n59515 & n59832;
  assign n59879 = ~n59872 & n59877;
  assign n10536 = n59878 | ~n59879;
  assign n59881 = P2_P3_INSTQUEUE_REG_11__1_ & ~n59823;
  assign n59882 = n59520 & n59819;
  assign n59883 = n59522 & n59811;
  assign n59884 = ~n59882 & ~n59883;
  assign n59885 = n59525 & n59818;
  assign n59886 = n59884 & ~n59885;
  assign n59887 = n59528 & n59832;
  assign n59888 = ~n59881 & n59886;
  assign n10541 = n59887 | ~n59888;
  assign n59890 = P2_P3_INSTQUEUE_REG_11__0_ & ~n59823;
  assign n59891 = n59533 & n59819;
  assign n59892 = n59535 & n59811;
  assign n59893 = ~n59891 & ~n59892;
  assign n59894 = n59538 & n59818;
  assign n59895 = n59893 & ~n59894;
  assign n59896 = n59541 & n59832;
  assign n59897 = ~n59890 & n59895;
  assign n10546 = n59896 | ~n59897;
  assign n59899 = ~P2_P3_INSTQUEUEWR_ADDR_REG_2_ & ~P2_P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n59900 = n59545 & n59899;
  assign n59901 = P2_P3_STATE2_REG_3_ & ~n59900;
  assign n59902 = n59384 & ~n59901;
  assign n59903 = n59402 & n59814;
  assign n59904 = ~n59900 & ~n59903;
  assign n59905 = n59552 & n59817;
  assign n59906 = n59405 & n59421;
  assign n59907 = ~n59905 & ~n59906;
  assign n59908 = n59401 & ~n59907;
  assign n59909 = n59904 & ~n59908;
  assign n59910 = n59902 & ~n59909;
  assign n59911 = P2_P3_INSTQUEUE_REG_10__7_ & ~n59910;
  assign n59912 = n59438 & n59906;
  assign n59913 = n59441 & n59900;
  assign n59914 = ~n59912 & ~n59913;
  assign n59915 = n59444 & n59905;
  assign n59916 = n59914 & ~n59915;
  assign n59917 = n59436 & n59907;
  assign n59918 = n59401 & ~n59917;
  assign n59919 = ~n59904 & ~n59918;
  assign n59920 = n59450 & n59919;
  assign n59921 = ~n59911 & n59916;
  assign n10551 = n59920 | ~n59921;
  assign n59923 = P2_P3_INSTQUEUE_REG_10__6_ & ~n59910;
  assign n59924 = n59455 & n59906;
  assign n59925 = n59457 & n59900;
  assign n59926 = ~n59924 & ~n59925;
  assign n59927 = n59460 & n59905;
  assign n59928 = n59926 & ~n59927;
  assign n59929 = n59463 & n59919;
  assign n59930 = ~n59923 & n59928;
  assign n10556 = n59929 | ~n59930;
  assign n59932 = P2_P3_INSTQUEUE_REG_10__5_ & ~n59910;
  assign n59933 = n59468 & n59906;
  assign n59934 = n59470 & n59900;
  assign n59935 = ~n59933 & ~n59934;
  assign n59936 = n59473 & n59905;
  assign n59937 = n59935 & ~n59936;
  assign n59938 = n59476 & n59919;
  assign n59939 = ~n59932 & n59937;
  assign n10561 = n59938 | ~n59939;
  assign n59941 = P2_P3_INSTQUEUE_REG_10__4_ & ~n59910;
  assign n59942 = n59481 & n59906;
  assign n59943 = n59483 & n59900;
  assign n59944 = ~n59942 & ~n59943;
  assign n59945 = n59486 & n59905;
  assign n59946 = n59944 & ~n59945;
  assign n59947 = n59489 & n59919;
  assign n59948 = ~n59941 & n59946;
  assign n10566 = n59947 | ~n59948;
  assign n59950 = P2_P3_INSTQUEUE_REG_10__3_ & ~n59910;
  assign n59951 = n59494 & n59906;
  assign n59952 = n59496 & n59900;
  assign n59953 = ~n59951 & ~n59952;
  assign n59954 = n59499 & n59905;
  assign n59955 = n59953 & ~n59954;
  assign n59956 = n59502 & n59919;
  assign n59957 = ~n59950 & n59955;
  assign n10571 = n59956 | ~n59957;
  assign n59959 = P2_P3_INSTQUEUE_REG_10__2_ & ~n59910;
  assign n59960 = n59507 & n59906;
  assign n59961 = n59509 & n59900;
  assign n59962 = ~n59960 & ~n59961;
  assign n59963 = n59512 & n59905;
  assign n59964 = n59962 & ~n59963;
  assign n59965 = n59515 & n59919;
  assign n59966 = ~n59959 & n59964;
  assign n10576 = n59965 | ~n59966;
  assign n59968 = P2_P3_INSTQUEUE_REG_10__1_ & ~n59910;
  assign n59969 = n59520 & n59906;
  assign n59970 = n59522 & n59900;
  assign n59971 = ~n59969 & ~n59970;
  assign n59972 = n59525 & n59905;
  assign n59973 = n59971 & ~n59972;
  assign n59974 = n59528 & n59919;
  assign n59975 = ~n59968 & n59973;
  assign n10581 = n59974 | ~n59975;
  assign n59977 = P2_P3_INSTQUEUE_REG_10__0_ & ~n59910;
  assign n59978 = n59533 & n59906;
  assign n59979 = n59535 & n59900;
  assign n59980 = ~n59978 & ~n59979;
  assign n59981 = n59538 & n59905;
  assign n59982 = n59980 & ~n59981;
  assign n59983 = n59541 & n59919;
  assign n59984 = ~n59977 & n59982;
  assign n10586 = n59983 | ~n59984;
  assign n59986 = n59393 & n59810;
  assign n59987 = P2_P3_STATE2_REG_3_ & ~n59986;
  assign n59988 = n59384 & ~n59987;
  assign n59989 = n59403 & n59814;
  assign n59990 = ~n59986 & ~n59989;
  assign n59991 = n59640 & n59817;
  assign n59992 = n59406 & n59421;
  assign n59993 = ~n59991 & ~n59992;
  assign n59994 = n59401 & ~n59993;
  assign n59995 = n59990 & ~n59994;
  assign n59996 = n59988 & ~n59995;
  assign n59997 = P2_P3_INSTQUEUE_REG_9__7_ & ~n59996;
  assign n59998 = n59438 & n59992;
  assign n59999 = n59441 & n59986;
  assign n60000 = ~n59998 & ~n59999;
  assign n60001 = n59444 & n59991;
  assign n60002 = n60000 & ~n60001;
  assign n60003 = n59436 & n59993;
  assign n60004 = n59401 & ~n60003;
  assign n60005 = ~n59990 & ~n60004;
  assign n60006 = n59450 & n60005;
  assign n60007 = ~n59997 & n60002;
  assign n10591 = n60006 | ~n60007;
  assign n60009 = P2_P3_INSTQUEUE_REG_9__6_ & ~n59996;
  assign n60010 = n59455 & n59992;
  assign n60011 = n59457 & n59986;
  assign n60012 = ~n60010 & ~n60011;
  assign n60013 = n59460 & n59991;
  assign n60014 = n60012 & ~n60013;
  assign n60015 = n59463 & n60005;
  assign n60016 = ~n60009 & n60014;
  assign n10596 = n60015 | ~n60016;
  assign n60018 = P2_P3_INSTQUEUE_REG_9__5_ & ~n59996;
  assign n60019 = n59468 & n59992;
  assign n60020 = n59470 & n59986;
  assign n60021 = ~n60019 & ~n60020;
  assign n60022 = n59473 & n59991;
  assign n60023 = n60021 & ~n60022;
  assign n60024 = n59476 & n60005;
  assign n60025 = ~n60018 & n60023;
  assign n10601 = n60024 | ~n60025;
  assign n60027 = P2_P3_INSTQUEUE_REG_9__4_ & ~n59996;
  assign n60028 = n59481 & n59992;
  assign n60029 = n59483 & n59986;
  assign n60030 = ~n60028 & ~n60029;
  assign n60031 = n59486 & n59991;
  assign n60032 = n60030 & ~n60031;
  assign n60033 = n59489 & n60005;
  assign n60034 = ~n60027 & n60032;
  assign n10606 = n60033 | ~n60034;
  assign n60036 = P2_P3_INSTQUEUE_REG_9__3_ & ~n59996;
  assign n60037 = n59494 & n59992;
  assign n60038 = n59496 & n59986;
  assign n60039 = ~n60037 & ~n60038;
  assign n60040 = n59499 & n59991;
  assign n60041 = n60039 & ~n60040;
  assign n60042 = n59502 & n60005;
  assign n60043 = ~n60036 & n60041;
  assign n10611 = n60042 | ~n60043;
  assign n60045 = P2_P3_INSTQUEUE_REG_9__2_ & ~n59996;
  assign n60046 = n59507 & n59992;
  assign n60047 = n59509 & n59986;
  assign n60048 = ~n60046 & ~n60047;
  assign n60049 = n59512 & n59991;
  assign n60050 = n60048 & ~n60049;
  assign n60051 = n59515 & n60005;
  assign n60052 = ~n60045 & n60050;
  assign n10616 = n60051 | ~n60052;
  assign n60054 = P2_P3_INSTQUEUE_REG_9__1_ & ~n59996;
  assign n60055 = n59520 & n59992;
  assign n60056 = n59522 & n59986;
  assign n60057 = ~n60055 & ~n60056;
  assign n60058 = n59525 & n59991;
  assign n60059 = n60057 & ~n60058;
  assign n60060 = n59528 & n60005;
  assign n60061 = ~n60054 & n60059;
  assign n10621 = n60060 | ~n60061;
  assign n60063 = P2_P3_INSTQUEUE_REG_9__0_ & ~n59996;
  assign n60064 = n59533 & n59992;
  assign n60065 = n59535 & n59986;
  assign n60066 = ~n60064 & ~n60065;
  assign n60067 = n59538 & n59991;
  assign n60068 = n60066 & ~n60067;
  assign n60069 = n59541 & n60005;
  assign n60070 = ~n60063 & n60068;
  assign n10626 = n60069 | ~n60070;
  assign n60072 = n59722 & n59899;
  assign n60073 = P2_P3_STATE2_REG_3_ & ~n60072;
  assign n60074 = n59384 & ~n60073;
  assign n60075 = n59726 & n59817;
  assign n60076 = n59421 & n59728;
  assign n60077 = ~n60075 & ~n60076;
  assign n60078 = n59401 & ~n60077;
  assign n60079 = n59395 & n59814;
  assign n60080 = ~n60078 & ~n60079;
  assign n60081 = n60074 & ~n60080;
  assign n60082 = P2_P3_INSTQUEUE_REG_8__7_ & ~n60081;
  assign n60083 = n59438 & n60076;
  assign n60084 = n59441 & n60072;
  assign n60085 = ~n60083 & ~n60084;
  assign n60086 = n59444 & n60075;
  assign n60087 = n60085 & ~n60086;
  assign n60088 = n59436 & n60077;
  assign n60089 = n59401 & ~n60088;
  assign n60090 = n60079 & ~n60089;
  assign n60091 = n59450 & n60090;
  assign n60092 = ~n60082 & n60087;
  assign n10631 = n60091 | ~n60092;
  assign n60094 = P2_P3_INSTQUEUE_REG_8__6_ & ~n60081;
  assign n60095 = n59455 & n60076;
  assign n60096 = n59457 & n60072;
  assign n60097 = ~n60095 & ~n60096;
  assign n60098 = n59460 & n60075;
  assign n60099 = n60097 & ~n60098;
  assign n60100 = n59463 & n60090;
  assign n60101 = ~n60094 & n60099;
  assign n10636 = n60100 | ~n60101;
  assign n60103 = P2_P3_INSTQUEUE_REG_8__5_ & ~n60081;
  assign n60104 = n59468 & n60076;
  assign n60105 = n59470 & n60072;
  assign n60106 = ~n60104 & ~n60105;
  assign n60107 = n59473 & n60075;
  assign n60108 = n60106 & ~n60107;
  assign n60109 = n59476 & n60090;
  assign n60110 = ~n60103 & n60108;
  assign n10641 = n60109 | ~n60110;
  assign n60112 = P2_P3_INSTQUEUE_REG_8__4_ & ~n60081;
  assign n60113 = n59481 & n60076;
  assign n60114 = n59483 & n60072;
  assign n60115 = ~n60113 & ~n60114;
  assign n60116 = n59486 & n60075;
  assign n60117 = n60115 & ~n60116;
  assign n60118 = n59489 & n60090;
  assign n60119 = ~n60112 & n60117;
  assign n10646 = n60118 | ~n60119;
  assign n60121 = P2_P3_INSTQUEUE_REG_8__3_ & ~n60081;
  assign n60122 = n59494 & n60076;
  assign n60123 = n59496 & n60072;
  assign n60124 = ~n60122 & ~n60123;
  assign n60125 = n59499 & n60075;
  assign n60126 = n60124 & ~n60125;
  assign n60127 = n59502 & n60090;
  assign n60128 = ~n60121 & n60126;
  assign n10651 = n60127 | ~n60128;
  assign n60130 = P2_P3_INSTQUEUE_REG_8__2_ & ~n60081;
  assign n60131 = n59507 & n60076;
  assign n60132 = n59509 & n60072;
  assign n60133 = ~n60131 & ~n60132;
  assign n60134 = n59512 & n60075;
  assign n60135 = n60133 & ~n60134;
  assign n60136 = n59515 & n60090;
  assign n60137 = ~n60130 & n60135;
  assign n10656 = n60136 | ~n60137;
  assign n60139 = P2_P3_INSTQUEUE_REG_8__1_ & ~n60081;
  assign n60140 = n59520 & n60076;
  assign n60141 = n59522 & n60072;
  assign n60142 = ~n60140 & ~n60141;
  assign n60143 = n59525 & n60075;
  assign n60144 = n60142 & ~n60143;
  assign n60145 = n59528 & n60090;
  assign n60146 = ~n60139 & n60144;
  assign n10661 = n60145 | ~n60146;
  assign n60148 = P2_P3_INSTQUEUE_REG_8__0_ & ~n60081;
  assign n60149 = n59533 & n60076;
  assign n60150 = n59535 & n60072;
  assign n60151 = ~n60149 & ~n60150;
  assign n60152 = n59538 & n60075;
  assign n60153 = n60151 & ~n60152;
  assign n60154 = n59541 & n60090;
  assign n60155 = ~n60148 & n60153;
  assign n10666 = n60154 | ~n60155;
  assign n60157 = P2_P3_STATE2_REG_3_ & ~n59389;
  assign n60158 = n59384 & ~n60157;
  assign n60159 = ~n59389 & ~n59417;
  assign n60160 = ~n59415 & n59426;
  assign n60161 = n59408 & n60160;
  assign n60162 = ~n59425 & ~n60161;
  assign n60163 = n59401 & ~n60162;
  assign n60164 = n60159 & ~n60163;
  assign n60165 = n60158 & ~n60164;
  assign n60166 = P2_P3_INSTQUEUE_REG_7__7_ & ~n60165;
  assign n60167 = n59425 & n59438;
  assign n60168 = n59389 & n59441;
  assign n60169 = ~n60167 & ~n60168;
  assign n60170 = n59444 & n60161;
  assign n60171 = n60169 & ~n60170;
  assign n60172 = n59436 & n60162;
  assign n60173 = n59401 & ~n60172;
  assign n60174 = ~n60159 & ~n60173;
  assign n60175 = n59450 & n60174;
  assign n60176 = ~n60166 & n60171;
  assign n10671 = n60175 | ~n60176;
  assign n60178 = P2_P3_INSTQUEUE_REG_7__6_ & ~n60165;
  assign n60179 = n59425 & n59455;
  assign n60180 = n59389 & n59457;
  assign n60181 = ~n60179 & ~n60180;
  assign n60182 = n59460 & n60161;
  assign n60183 = n60181 & ~n60182;
  assign n60184 = n59463 & n60174;
  assign n60185 = ~n60178 & n60183;
  assign n10676 = n60184 | ~n60185;
  assign n60187 = P2_P3_INSTQUEUE_REG_7__5_ & ~n60165;
  assign n60188 = n59425 & n59468;
  assign n60189 = n59389 & n59470;
  assign n60190 = ~n60188 & ~n60189;
  assign n60191 = n59473 & n60161;
  assign n60192 = n60190 & ~n60191;
  assign n60193 = n59476 & n60174;
  assign n60194 = ~n60187 & n60192;
  assign n10681 = n60193 | ~n60194;
  assign n60196 = P2_P3_INSTQUEUE_REG_7__4_ & ~n60165;
  assign n60197 = n59425 & n59481;
  assign n60198 = n59389 & n59483;
  assign n60199 = ~n60197 & ~n60198;
  assign n60200 = n59486 & n60161;
  assign n60201 = n60199 & ~n60200;
  assign n60202 = n59489 & n60174;
  assign n60203 = ~n60196 & n60201;
  assign n10686 = n60202 | ~n60203;
  assign n60205 = P2_P3_INSTQUEUE_REG_7__3_ & ~n60165;
  assign n60206 = n59425 & n59494;
  assign n60207 = n59389 & n59496;
  assign n60208 = ~n60206 & ~n60207;
  assign n60209 = n59499 & n60161;
  assign n60210 = n60208 & ~n60209;
  assign n60211 = n59502 & n60174;
  assign n60212 = ~n60205 & n60210;
  assign n10691 = n60211 | ~n60212;
  assign n60214 = P2_P3_INSTQUEUE_REG_7__2_ & ~n60165;
  assign n60215 = n59425 & n59507;
  assign n60216 = n59389 & n59509;
  assign n60217 = ~n60215 & ~n60216;
  assign n60218 = n59512 & n60161;
  assign n60219 = n60217 & ~n60218;
  assign n60220 = n59515 & n60174;
  assign n60221 = ~n60214 & n60219;
  assign n10696 = n60220 | ~n60221;
  assign n60223 = P2_P3_INSTQUEUE_REG_7__1_ & ~n60165;
  assign n60224 = n59425 & n59520;
  assign n60225 = n59389 & n59522;
  assign n60226 = ~n60224 & ~n60225;
  assign n60227 = n59525 & n60161;
  assign n60228 = n60226 & ~n60227;
  assign n60229 = n59528 & n60174;
  assign n60230 = ~n60223 & n60228;
  assign n10701 = n60229 | ~n60230;
  assign n60232 = P2_P3_INSTQUEUE_REG_7__0_ & ~n60165;
  assign n60233 = n59425 & n59533;
  assign n60234 = n59389 & n59535;
  assign n60235 = ~n60233 & ~n60234;
  assign n60236 = n59538 & n60161;
  assign n60237 = n60235 & ~n60236;
  assign n60238 = n59541 & n60174;
  assign n60239 = ~n60232 & n60237;
  assign n10706 = n60238 | ~n60239;
  assign n60241 = ~P2_P3_INSTQUEUEWR_ADDR_REG_3_ & P2_P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n60242 = n59546 & n60241;
  assign n60243 = P2_P3_STATE2_REG_3_ & ~n60242;
  assign n60244 = n59384 & ~n60243;
  assign n60245 = n59402 & n59416;
  assign n60246 = ~n60242 & ~n60245;
  assign n60247 = n59552 & n60160;
  assign n60248 = n59405 & n59424;
  assign n60249 = ~n60247 & ~n60248;
  assign n60250 = n59401 & ~n60249;
  assign n60251 = n60246 & ~n60250;
  assign n60252 = n60244 & ~n60251;
  assign n60253 = P2_P3_INSTQUEUE_REG_6__7_ & ~n60252;
  assign n60254 = n59438 & n60248;
  assign n60255 = n59441 & n60242;
  assign n60256 = ~n60254 & ~n60255;
  assign n60257 = n59444 & n60247;
  assign n60258 = n60256 & ~n60257;
  assign n60259 = n59436 & n60249;
  assign n60260 = n59401 & ~n60259;
  assign n60261 = ~n60246 & ~n60260;
  assign n60262 = n59450 & n60261;
  assign n60263 = ~n60253 & n60258;
  assign n10711 = n60262 | ~n60263;
  assign n60265 = P2_P3_INSTQUEUE_REG_6__6_ & ~n60252;
  assign n60266 = n59455 & n60248;
  assign n60267 = n59457 & n60242;
  assign n60268 = ~n60266 & ~n60267;
  assign n60269 = n59460 & n60247;
  assign n60270 = n60268 & ~n60269;
  assign n60271 = n59463 & n60261;
  assign n60272 = ~n60265 & n60270;
  assign n10716 = n60271 | ~n60272;
  assign n60274 = P2_P3_INSTQUEUE_REG_6__5_ & ~n60252;
  assign n60275 = n59468 & n60248;
  assign n60276 = n59470 & n60242;
  assign n60277 = ~n60275 & ~n60276;
  assign n60278 = n59473 & n60247;
  assign n60279 = n60277 & ~n60278;
  assign n60280 = n59476 & n60261;
  assign n60281 = ~n60274 & n60279;
  assign n10721 = n60280 | ~n60281;
  assign n60283 = P2_P3_INSTQUEUE_REG_6__4_ & ~n60252;
  assign n60284 = n59481 & n60248;
  assign n60285 = n59483 & n60242;
  assign n60286 = ~n60284 & ~n60285;
  assign n60287 = n59486 & n60247;
  assign n60288 = n60286 & ~n60287;
  assign n60289 = n59489 & n60261;
  assign n60290 = ~n60283 & n60288;
  assign n10726 = n60289 | ~n60290;
  assign n60292 = P2_P3_INSTQUEUE_REG_6__3_ & ~n60252;
  assign n60293 = n59494 & n60248;
  assign n60294 = n59496 & n60242;
  assign n60295 = ~n60293 & ~n60294;
  assign n60296 = n59499 & n60247;
  assign n60297 = n60295 & ~n60296;
  assign n60298 = n59502 & n60261;
  assign n60299 = ~n60292 & n60297;
  assign n10731 = n60298 | ~n60299;
  assign n60301 = P2_P3_INSTQUEUE_REG_6__2_ & ~n60252;
  assign n60302 = n59507 & n60248;
  assign n60303 = n59509 & n60242;
  assign n60304 = ~n60302 & ~n60303;
  assign n60305 = n59512 & n60247;
  assign n60306 = n60304 & ~n60305;
  assign n60307 = n59515 & n60261;
  assign n60308 = ~n60301 & n60306;
  assign n10736 = n60307 | ~n60308;
  assign n60310 = P2_P3_INSTQUEUE_REG_6__1_ & ~n60252;
  assign n60311 = n59520 & n60248;
  assign n60312 = n59522 & n60242;
  assign n60313 = ~n60311 & ~n60312;
  assign n60314 = n59525 & n60247;
  assign n60315 = n60313 & ~n60314;
  assign n60316 = n59528 & n60261;
  assign n60317 = ~n60310 & n60315;
  assign n10741 = n60316 | ~n60317;
  assign n60319 = P2_P3_INSTQUEUE_REG_6__0_ & ~n60252;
  assign n60320 = n59533 & n60248;
  assign n60321 = n59535 & n60242;
  assign n60322 = ~n60320 & ~n60321;
  assign n60323 = n59538 & n60247;
  assign n60324 = n60322 & ~n60323;
  assign n60325 = n59541 & n60261;
  assign n60326 = ~n60319 & n60324;
  assign n10746 = n60325 | ~n60326;
  assign n60328 = ~P2_P3_INSTQUEUEWR_ADDR_REG_3_ & P2_P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n60329 = n59393 & n60328;
  assign n60330 = P2_P3_STATE2_REG_3_ & ~n60329;
  assign n60331 = n59384 & ~n60330;
  assign n60332 = n59403 & n59416;
  assign n60333 = ~n60329 & ~n60332;
  assign n60334 = n59640 & n60160;
  assign n60335 = n59406 & n59424;
  assign n60336 = ~n60334 & ~n60335;
  assign n60337 = n59401 & ~n60336;
  assign n60338 = n60333 & ~n60337;
  assign n60339 = n60331 & ~n60338;
  assign n60340 = P2_P3_INSTQUEUE_REG_5__7_ & ~n60339;
  assign n60341 = n59438 & n60335;
  assign n60342 = n59441 & n60329;
  assign n60343 = ~n60341 & ~n60342;
  assign n60344 = n59444 & n60334;
  assign n60345 = n60343 & ~n60344;
  assign n60346 = n59436 & n60336;
  assign n60347 = n59401 & ~n60346;
  assign n60348 = ~n60333 & ~n60347;
  assign n60349 = n59450 & n60348;
  assign n60350 = ~n60340 & n60345;
  assign n10751 = n60349 | ~n60350;
  assign n60352 = P2_P3_INSTQUEUE_REG_5__6_ & ~n60339;
  assign n60353 = n59455 & n60335;
  assign n60354 = n59457 & n60329;
  assign n60355 = ~n60353 & ~n60354;
  assign n60356 = n59460 & n60334;
  assign n60357 = n60355 & ~n60356;
  assign n60358 = n59463 & n60348;
  assign n60359 = ~n60352 & n60357;
  assign n10756 = n60358 | ~n60359;
  assign n60361 = P2_P3_INSTQUEUE_REG_5__5_ & ~n60339;
  assign n60362 = n59468 & n60335;
  assign n60363 = n59470 & n60329;
  assign n60364 = ~n60362 & ~n60363;
  assign n60365 = n59473 & n60334;
  assign n60366 = n60364 & ~n60365;
  assign n60367 = n59476 & n60348;
  assign n60368 = ~n60361 & n60366;
  assign n10761 = n60367 | ~n60368;
  assign n60370 = P2_P3_INSTQUEUE_REG_5__4_ & ~n60339;
  assign n60371 = n59481 & n60335;
  assign n60372 = n59483 & n60329;
  assign n60373 = ~n60371 & ~n60372;
  assign n60374 = n59486 & n60334;
  assign n60375 = n60373 & ~n60374;
  assign n60376 = n59489 & n60348;
  assign n60377 = ~n60370 & n60375;
  assign n10766 = n60376 | ~n60377;
  assign n60379 = P2_P3_INSTQUEUE_REG_5__3_ & ~n60339;
  assign n60380 = n59494 & n60335;
  assign n60381 = n59496 & n60329;
  assign n60382 = ~n60380 & ~n60381;
  assign n60383 = n59499 & n60334;
  assign n60384 = n60382 & ~n60383;
  assign n60385 = n59502 & n60348;
  assign n60386 = ~n60379 & n60384;
  assign n10771 = n60385 | ~n60386;
  assign n60388 = P2_P3_INSTQUEUE_REG_5__2_ & ~n60339;
  assign n60389 = n59507 & n60335;
  assign n60390 = n59509 & n60329;
  assign n60391 = ~n60389 & ~n60390;
  assign n60392 = n59512 & n60334;
  assign n60393 = n60391 & ~n60392;
  assign n60394 = n59515 & n60348;
  assign n60395 = ~n60388 & n60393;
  assign n10776 = n60394 | ~n60395;
  assign n60397 = P2_P3_INSTQUEUE_REG_5__1_ & ~n60339;
  assign n60398 = n59520 & n60335;
  assign n60399 = n59522 & n60329;
  assign n60400 = ~n60398 & ~n60399;
  assign n60401 = n59525 & n60334;
  assign n60402 = n60400 & ~n60401;
  assign n60403 = n59528 & n60348;
  assign n60404 = ~n60397 & n60402;
  assign n10781 = n60403 | ~n60404;
  assign n60406 = P2_P3_INSTQUEUE_REG_5__0_ & ~n60339;
  assign n60407 = n59533 & n60335;
  assign n60408 = n59535 & n60329;
  assign n60409 = ~n60407 & ~n60408;
  assign n60410 = n59538 & n60334;
  assign n60411 = n60409 & ~n60410;
  assign n60412 = n59541 & n60348;
  assign n60413 = ~n60406 & n60411;
  assign n10786 = n60412 | ~n60413;
  assign n60415 = n59424 & n59728;
  assign n60416 = n59438 & n60415;
  assign n60417 = ~P2_P3_INSTQUEUEWR_ADDR_REG_3_ & ~P2_P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n60418 = n59546 & n60417;
  assign n60419 = n59441 & n60418;
  assign n60420 = n59401 & ~n59436;
  assign n60421 = n59395 & n59416;
  assign n60422 = ~n60420 & n60421;
  assign n60423 = n59450 & n60422;
  assign n60424 = ~n60416 & ~n60419;
  assign n60425 = ~n60423 & n60424;
  assign n60426 = n59726 & n60160;
  assign n60427 = n59444 & n60426;
  assign n60428 = n60425 & ~n60427;
  assign n60429 = P2_P3_STATE2_REG_3_ & ~n60418;
  assign n60430 = n59384 & ~n60429;
  assign n60431 = ~n60415 & ~n60426;
  assign n60432 = n59401 & ~n60431;
  assign n60433 = ~n60421 & ~n60432;
  assign n60434 = n60430 & ~n60433;
  assign n60435 = P2_P3_INSTQUEUE_REG_4__7_ & ~n60434;
  assign n10791 = ~n60428 | n60435;
  assign n60437 = n59455 & n60415;
  assign n60438 = n59457 & n60418;
  assign n60439 = n59463 & n60422;
  assign n60440 = ~n60437 & ~n60438;
  assign n60441 = ~n60439 & n60440;
  assign n60442 = n59460 & n60426;
  assign n60443 = n60441 & ~n60442;
  assign n60444 = P2_P3_INSTQUEUE_REG_4__6_ & ~n60434;
  assign n10796 = ~n60443 | n60444;
  assign n60446 = n59468 & n60415;
  assign n60447 = n59470 & n60418;
  assign n60448 = n59476 & n60422;
  assign n60449 = ~n60446 & ~n60447;
  assign n60450 = ~n60448 & n60449;
  assign n60451 = n59473 & n60426;
  assign n60452 = n60450 & ~n60451;
  assign n60453 = P2_P3_INSTQUEUE_REG_4__5_ & ~n60434;
  assign n10801 = ~n60452 | n60453;
  assign n60455 = n59481 & n60415;
  assign n60456 = n59483 & n60418;
  assign n60457 = n59489 & n60422;
  assign n60458 = ~n60455 & ~n60456;
  assign n60459 = ~n60457 & n60458;
  assign n60460 = n59486 & n60426;
  assign n60461 = n60459 & ~n60460;
  assign n60462 = P2_P3_INSTQUEUE_REG_4__4_ & ~n60434;
  assign n10806 = ~n60461 | n60462;
  assign n60464 = n59494 & n60415;
  assign n60465 = n59496 & n60418;
  assign n60466 = n59502 & n60422;
  assign n60467 = ~n60464 & ~n60465;
  assign n60468 = ~n60466 & n60467;
  assign n60469 = n59499 & n60426;
  assign n60470 = n60468 & ~n60469;
  assign n60471 = P2_P3_INSTQUEUE_REG_4__3_ & ~n60434;
  assign n10811 = ~n60470 | n60471;
  assign n60473 = n59507 & n60415;
  assign n60474 = n59509 & n60418;
  assign n60475 = n59515 & n60422;
  assign n60476 = ~n60473 & ~n60474;
  assign n60477 = ~n60475 & n60476;
  assign n60478 = n59512 & n60426;
  assign n60479 = n60477 & ~n60478;
  assign n60480 = P2_P3_INSTQUEUE_REG_4__2_ & ~n60434;
  assign n10816 = ~n60479 | n60480;
  assign n60482 = n59520 & n60415;
  assign n60483 = n59522 & n60418;
  assign n60484 = n59528 & n60422;
  assign n60485 = ~n60482 & ~n60483;
  assign n60486 = ~n60484 & n60485;
  assign n60487 = n59525 & n60426;
  assign n60488 = n60486 & ~n60487;
  assign n60489 = P2_P3_INSTQUEUE_REG_4__1_ & ~n60434;
  assign n10821 = ~n60488 | n60489;
  assign n60491 = n59533 & n60415;
  assign n60492 = n59535 & n60418;
  assign n60493 = n59541 & n60422;
  assign n60494 = ~n60491 & ~n60492;
  assign n60495 = ~n60493 & n60494;
  assign n60496 = n59538 & n60426;
  assign n60497 = n60495 & ~n60496;
  assign n60498 = P2_P3_INSTQUEUE_REG_4__0_ & ~n60434;
  assign n10826 = ~n60497 | n60498;
  assign n60500 = n59411 & n59420;
  assign n60501 = n59412 & n60500;
  assign n60502 = n59438 & n60501;
  assign n60503 = ~P2_P3_INSTQUEUEWR_ADDR_REG_3_ & ~P2_P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n60504 = n59377 & n60503;
  assign n60505 = n59441 & n60504;
  assign n60506 = n59388 & n59391;
  assign n60507 = n59396 & n60506;
  assign n60508 = ~n60504 & ~n60507;
  assign n60509 = ~n60420 & ~n60508;
  assign n60510 = n59450 & n60509;
  assign n60511 = ~n60502 & ~n60505;
  assign n60512 = ~n60510 & n60511;
  assign n60513 = n59415 & n59426;
  assign n60514 = n59408 & n60513;
  assign n60515 = n59444 & n60514;
  assign n60516 = n60512 & ~n60515;
  assign n60517 = P2_P3_STATE2_REG_3_ & ~n60504;
  assign n60518 = n59384 & ~n60517;
  assign n60519 = ~n60501 & ~n60514;
  assign n60520 = n59401 & ~n60519;
  assign n60521 = n60508 & ~n60520;
  assign n60522 = n60518 & ~n60521;
  assign n60523 = P2_P3_INSTQUEUE_REG_3__7_ & ~n60522;
  assign n10831 = ~n60516 | n60523;
  assign n60525 = n59455 & n60501;
  assign n60526 = n59457 & n60504;
  assign n60527 = n59463 & n60509;
  assign n60528 = ~n60525 & ~n60526;
  assign n60529 = ~n60527 & n60528;
  assign n60530 = n59460 & n60514;
  assign n60531 = n60529 & ~n60530;
  assign n60532 = P2_P3_INSTQUEUE_REG_3__6_ & ~n60522;
  assign n10836 = ~n60531 | n60532;
  assign n60534 = n59468 & n60501;
  assign n60535 = n59470 & n60504;
  assign n60536 = n59476 & n60509;
  assign n60537 = ~n60534 & ~n60535;
  assign n60538 = ~n60536 & n60537;
  assign n60539 = n59473 & n60514;
  assign n60540 = n60538 & ~n60539;
  assign n60541 = P2_P3_INSTQUEUE_REG_3__5_ & ~n60522;
  assign n10841 = ~n60540 | n60541;
  assign n60543 = n59481 & n60501;
  assign n60544 = n59483 & n60504;
  assign n60545 = n59489 & n60509;
  assign n60546 = ~n60543 & ~n60544;
  assign n60547 = ~n60545 & n60546;
  assign n60548 = n59486 & n60514;
  assign n60549 = n60547 & ~n60548;
  assign n60550 = P2_P3_INSTQUEUE_REG_3__4_ & ~n60522;
  assign n10846 = ~n60549 | n60550;
  assign n60552 = n59494 & n60501;
  assign n60553 = n59496 & n60504;
  assign n60554 = n59502 & n60509;
  assign n60555 = ~n60552 & ~n60553;
  assign n60556 = ~n60554 & n60555;
  assign n60557 = n59499 & n60514;
  assign n60558 = n60556 & ~n60557;
  assign n60559 = P2_P3_INSTQUEUE_REG_3__3_ & ~n60522;
  assign n10851 = ~n60558 | n60559;
  assign n60561 = n59507 & n60501;
  assign n60562 = n59509 & n60504;
  assign n60563 = n59515 & n60509;
  assign n60564 = ~n60561 & ~n60562;
  assign n60565 = ~n60563 & n60564;
  assign n60566 = n59512 & n60514;
  assign n60567 = n60565 & ~n60566;
  assign n60568 = P2_P3_INSTQUEUE_REG_3__2_ & ~n60522;
  assign n10856 = ~n60567 | n60568;
  assign n60570 = n59520 & n60501;
  assign n60571 = n59522 & n60504;
  assign n60572 = n59528 & n60509;
  assign n60573 = ~n60570 & ~n60571;
  assign n60574 = ~n60572 & n60573;
  assign n60575 = n59525 & n60514;
  assign n60576 = n60574 & ~n60575;
  assign n60577 = P2_P3_INSTQUEUE_REG_3__1_ & ~n60522;
  assign n10861 = ~n60576 | n60577;
  assign n60579 = n59533 & n60501;
  assign n60580 = n59535 & n60504;
  assign n60581 = n59541 & n60509;
  assign n60582 = ~n60579 & ~n60580;
  assign n60583 = ~n60581 & n60582;
  assign n60584 = n59538 & n60514;
  assign n60585 = n60583 & ~n60584;
  assign n60586 = P2_P3_INSTQUEUE_REG_3__0_ & ~n60522;
  assign n10866 = ~n60585 | n60586;
  assign n60588 = n59405 & n60500;
  assign n60589 = n59438 & n60588;
  assign n60590 = n59899 & n60241;
  assign n60591 = n59441 & n60590;
  assign n60592 = n59402 & n60506;
  assign n60593 = ~n60590 & ~n60592;
  assign n60594 = ~n60420 & ~n60593;
  assign n60595 = n59450 & n60594;
  assign n60596 = ~n60589 & ~n60591;
  assign n60597 = ~n60595 & n60596;
  assign n60598 = n59552 & n60513;
  assign n60599 = n59444 & n60598;
  assign n60600 = n60597 & ~n60599;
  assign n60601 = P2_P3_STATE2_REG_3_ & ~n60590;
  assign n60602 = n59384 & ~n60601;
  assign n60603 = ~n60588 & ~n60598;
  assign n60604 = n59401 & ~n60603;
  assign n60605 = n60593 & ~n60604;
  assign n60606 = n60602 & ~n60605;
  assign n60607 = P2_P3_INSTQUEUE_REG_2__7_ & ~n60606;
  assign n10871 = ~n60600 | n60607;
  assign n60609 = n59455 & n60588;
  assign n60610 = n59457 & n60590;
  assign n60611 = n59463 & n60594;
  assign n60612 = ~n60609 & ~n60610;
  assign n60613 = ~n60611 & n60612;
  assign n60614 = n59460 & n60598;
  assign n60615 = n60613 & ~n60614;
  assign n60616 = P2_P3_INSTQUEUE_REG_2__6_ & ~n60606;
  assign n10876 = ~n60615 | n60616;
  assign n60618 = n59468 & n60588;
  assign n60619 = n59470 & n60590;
  assign n60620 = n59476 & n60594;
  assign n60621 = ~n60618 & ~n60619;
  assign n60622 = ~n60620 & n60621;
  assign n60623 = n59473 & n60598;
  assign n60624 = n60622 & ~n60623;
  assign n60625 = P2_P3_INSTQUEUE_REG_2__5_ & ~n60606;
  assign n10881 = ~n60624 | n60625;
  assign n60627 = n59481 & n60588;
  assign n60628 = n59483 & n60590;
  assign n60629 = n59489 & n60594;
  assign n60630 = ~n60627 & ~n60628;
  assign n60631 = ~n60629 & n60630;
  assign n60632 = n59486 & n60598;
  assign n60633 = n60631 & ~n60632;
  assign n60634 = P2_P3_INSTQUEUE_REG_2__4_ & ~n60606;
  assign n10886 = ~n60633 | n60634;
  assign n60636 = n59494 & n60588;
  assign n60637 = n59496 & n60590;
  assign n60638 = n59502 & n60594;
  assign n60639 = ~n60636 & ~n60637;
  assign n60640 = ~n60638 & n60639;
  assign n60641 = n59499 & n60598;
  assign n60642 = n60640 & ~n60641;
  assign n60643 = P2_P3_INSTQUEUE_REG_2__3_ & ~n60606;
  assign n10891 = ~n60642 | n60643;
  assign n60645 = n59507 & n60588;
  assign n60646 = n59509 & n60590;
  assign n60647 = n59515 & n60594;
  assign n60648 = ~n60645 & ~n60646;
  assign n60649 = ~n60647 & n60648;
  assign n60650 = n59512 & n60598;
  assign n60651 = n60649 & ~n60650;
  assign n60652 = P2_P3_INSTQUEUE_REG_2__2_ & ~n60606;
  assign n10896 = ~n60651 | n60652;
  assign n60654 = n59520 & n60588;
  assign n60655 = n59522 & n60590;
  assign n60656 = n59528 & n60594;
  assign n60657 = ~n60654 & ~n60655;
  assign n60658 = ~n60656 & n60657;
  assign n60659 = n59525 & n60598;
  assign n60660 = n60658 & ~n60659;
  assign n60661 = P2_P3_INSTQUEUE_REG_2__1_ & ~n60606;
  assign n10901 = ~n60660 | n60661;
  assign n60663 = n59533 & n60588;
  assign n60664 = n59535 & n60590;
  assign n60665 = n59541 & n60594;
  assign n60666 = ~n60663 & ~n60664;
  assign n60667 = ~n60665 & n60666;
  assign n60668 = n59538 & n60598;
  assign n60669 = n60667 & ~n60668;
  assign n60670 = P2_P3_INSTQUEUE_REG_2__0_ & ~n60606;
  assign n10906 = ~n60669 | n60670;
  assign n60672 = n59406 & n60500;
  assign n60673 = n59438 & n60672;
  assign n60674 = n59393 & n60503;
  assign n60675 = n59441 & n60674;
  assign n60676 = n59403 & n60506;
  assign n60677 = ~n60674 & ~n60676;
  assign n60678 = ~n60420 & ~n60677;
  assign n60679 = n59450 & n60678;
  assign n60680 = ~n60673 & ~n60675;
  assign n60681 = ~n60679 & n60680;
  assign n60682 = n59640 & n60513;
  assign n60683 = n59444 & n60682;
  assign n60684 = n60681 & ~n60683;
  assign n60685 = P2_P3_STATE2_REG_3_ & ~n60674;
  assign n60686 = n59384 & ~n60685;
  assign n60687 = ~n60672 & ~n60682;
  assign n60688 = n59401 & ~n60687;
  assign n60689 = n60677 & ~n60688;
  assign n60690 = n60686 & ~n60689;
  assign n60691 = P2_P3_INSTQUEUE_REG_1__7_ & ~n60690;
  assign n10911 = ~n60684 | n60691;
  assign n60693 = n59455 & n60672;
  assign n60694 = n59457 & n60674;
  assign n60695 = n59463 & n60678;
  assign n60696 = ~n60693 & ~n60694;
  assign n60697 = ~n60695 & n60696;
  assign n60698 = n59460 & n60682;
  assign n60699 = n60697 & ~n60698;
  assign n60700 = P2_P3_INSTQUEUE_REG_1__6_ & ~n60690;
  assign n10916 = ~n60699 | n60700;
  assign n60702 = n59468 & n60672;
  assign n60703 = n59470 & n60674;
  assign n60704 = n59476 & n60678;
  assign n60705 = ~n60702 & ~n60703;
  assign n60706 = ~n60704 & n60705;
  assign n60707 = n59473 & n60682;
  assign n60708 = n60706 & ~n60707;
  assign n60709 = P2_P3_INSTQUEUE_REG_1__5_ & ~n60690;
  assign n10921 = ~n60708 | n60709;
  assign n60711 = n59481 & n60672;
  assign n60712 = n59483 & n60674;
  assign n60713 = n59489 & n60678;
  assign n60714 = ~n60711 & ~n60712;
  assign n60715 = ~n60713 & n60714;
  assign n60716 = n59486 & n60682;
  assign n60717 = n60715 & ~n60716;
  assign n60718 = P2_P3_INSTQUEUE_REG_1__4_ & ~n60690;
  assign n10926 = ~n60717 | n60718;
  assign n60720 = n59494 & n60672;
  assign n60721 = n59496 & n60674;
  assign n60722 = n59502 & n60678;
  assign n60723 = ~n60720 & ~n60721;
  assign n60724 = ~n60722 & n60723;
  assign n60725 = n59499 & n60682;
  assign n60726 = n60724 & ~n60725;
  assign n60727 = P2_P3_INSTQUEUE_REG_1__3_ & ~n60690;
  assign n10931 = ~n60726 | n60727;
  assign n60729 = n59507 & n60672;
  assign n60730 = n59509 & n60674;
  assign n60731 = n59515 & n60678;
  assign n60732 = ~n60729 & ~n60730;
  assign n60733 = ~n60731 & n60732;
  assign n60734 = n59512 & n60682;
  assign n60735 = n60733 & ~n60734;
  assign n60736 = P2_P3_INSTQUEUE_REG_1__2_ & ~n60690;
  assign n10936 = ~n60735 | n60736;
  assign n60738 = n59520 & n60672;
  assign n60739 = n59522 & n60674;
  assign n60740 = n59528 & n60678;
  assign n60741 = ~n60738 & ~n60739;
  assign n60742 = ~n60740 & n60741;
  assign n60743 = n59525 & n60682;
  assign n60744 = n60742 & ~n60743;
  assign n60745 = P2_P3_INSTQUEUE_REG_1__1_ & ~n60690;
  assign n10941 = ~n60744 | n60745;
  assign n60747 = n59533 & n60672;
  assign n60748 = n59535 & n60674;
  assign n60749 = n59541 & n60678;
  assign n60750 = ~n60747 & ~n60748;
  assign n60751 = ~n60749 & n60750;
  assign n60752 = n59538 & n60682;
  assign n60753 = n60751 & ~n60752;
  assign n60754 = P2_P3_INSTQUEUE_REG_1__0_ & ~n60690;
  assign n10946 = ~n60753 | n60754;
  assign n60756 = n59728 & n60500;
  assign n60757 = n59438 & n60756;
  assign n60758 = n59899 & n60417;
  assign n60759 = n59441 & n60758;
  assign n60760 = n59395 & n60506;
  assign n60761 = ~n60420 & n60760;
  assign n60762 = n59450 & n60761;
  assign n60763 = ~n60757 & ~n60759;
  assign n60764 = ~n60762 & n60763;
  assign n60765 = n59726 & n60513;
  assign n60766 = n59444 & n60765;
  assign n60767 = n60764 & ~n60766;
  assign n60768 = P2_P3_STATE2_REG_3_ & ~n60758;
  assign n60769 = n59384 & ~n60768;
  assign n60770 = ~n60756 & ~n60765;
  assign n60771 = n59401 & ~n60770;
  assign n60772 = ~n60760 & ~n60771;
  assign n60773 = n60769 & ~n60772;
  assign n60774 = P2_P3_INSTQUEUE_REG_0__7_ & ~n60773;
  assign n10951 = ~n60767 | n60774;
  assign n60776 = n59455 & n60756;
  assign n60777 = n59457 & n60758;
  assign n60778 = n59463 & n60761;
  assign n60779 = ~n60776 & ~n60777;
  assign n60780 = ~n60778 & n60779;
  assign n60781 = n59460 & n60765;
  assign n60782 = n60780 & ~n60781;
  assign n60783 = P2_P3_INSTQUEUE_REG_0__6_ & ~n60773;
  assign n10956 = ~n60782 | n60783;
  assign n60785 = n59468 & n60756;
  assign n60786 = n59470 & n60758;
  assign n60787 = n59476 & n60761;
  assign n60788 = ~n60785 & ~n60786;
  assign n60789 = ~n60787 & n60788;
  assign n60790 = n59473 & n60765;
  assign n60791 = n60789 & ~n60790;
  assign n60792 = P2_P3_INSTQUEUE_REG_0__5_ & ~n60773;
  assign n10961 = ~n60791 | n60792;
  assign n60794 = n59481 & n60756;
  assign n60795 = n59483 & n60758;
  assign n60796 = n59489 & n60761;
  assign n60797 = ~n60794 & ~n60795;
  assign n60798 = ~n60796 & n60797;
  assign n60799 = n59486 & n60765;
  assign n60800 = n60798 & ~n60799;
  assign n60801 = P2_P3_INSTQUEUE_REG_0__4_ & ~n60773;
  assign n10966 = ~n60800 | n60801;
  assign n60803 = n59494 & n60756;
  assign n60804 = n59496 & n60758;
  assign n60805 = n59502 & n60761;
  assign n60806 = ~n60803 & ~n60804;
  assign n60807 = ~n60805 & n60806;
  assign n60808 = n59499 & n60765;
  assign n60809 = n60807 & ~n60808;
  assign n60810 = P2_P3_INSTQUEUE_REG_0__3_ & ~n60773;
  assign n10971 = ~n60809 | n60810;
  assign n60812 = n59507 & n60756;
  assign n60813 = n59509 & n60758;
  assign n60814 = n59515 & n60761;
  assign n60815 = ~n60812 & ~n60813;
  assign n60816 = ~n60814 & n60815;
  assign n60817 = n59512 & n60765;
  assign n60818 = n60816 & ~n60817;
  assign n60819 = P2_P3_INSTQUEUE_REG_0__2_ & ~n60773;
  assign n10976 = ~n60818 | n60819;
  assign n60821 = n59520 & n60756;
  assign n60822 = n59522 & n60758;
  assign n60823 = n59528 & n60761;
  assign n60824 = ~n60821 & ~n60822;
  assign n60825 = ~n60823 & n60824;
  assign n60826 = n59525 & n60765;
  assign n60827 = n60825 & ~n60826;
  assign n60828 = P2_P3_INSTQUEUE_REG_0__1_ & ~n60773;
  assign n10981 = ~n60827 | n60828;
  assign n60830 = n59533 & n60756;
  assign n60831 = n59535 & n60758;
  assign n60832 = n59541 & n60761;
  assign n60833 = ~n60830 & ~n60831;
  assign n60834 = ~n60832 & n60833;
  assign n60835 = n59538 & n60765;
  assign n60836 = n60834 & ~n60835;
  assign n60837 = P2_P3_INSTQUEUE_REG_0__0_ & ~n60773;
  assign n10986 = ~n60836 | n60837;
  assign n60839 = P2_P3_STATE2_REG_3_ & ~P2_P3_STATE2_REG_0_;
  assign n60840 = P2_P3_STATE2_REG_0_ & P2_P3_FLUSH_REG;
  assign n60841 = n58679 & n60840;
  assign n60842 = ~n60839 & ~n60841;
  assign n60843 = ~n59211 & n59321;
  assign n60844 = n60842 & ~n60843;
  assign n60845 = P2_P3_INSTQUEUERD_ADDR_REG_4_ & n60844;
  assign n60846 = ~n59254 & n59327;
  assign n60847 = n59046 & n60846;
  assign n60848 = ~n60844 & n60847;
  assign n10991 = n60845 | n60848;
  assign n60850 = ~n59245 & n59327;
  assign n60851 = ~n58718 & ~n59218;
  assign n60852 = n59336 & ~n60851;
  assign n60853 = ~n60850 & ~n60852;
  assign n60854 = ~n60844 & ~n60853;
  assign n60855 = P2_P3_INSTQUEUERD_ADDR_REG_3_ & n60844;
  assign n10996 = n60854 | n60855;
  assign n60857 = ~n59169 & n59336;
  assign n60858 = P2_P3_STATE2_REG_1_ & ~n59343;
  assign n60859 = ~n59352 & n60858;
  assign n60860 = ~n60857 & ~n60859;
  assign n60861 = ~n59185 & n59327;
  assign n60862 = n60860 & ~n60861;
  assign n60863 = ~n60844 & ~n60862;
  assign n60864 = P2_P3_INSTQUEUERD_ADDR_REG_2_ & n60844;
  assign n11001 = n60863 | n60864;
  assign n60866 = n59281 & n59336;
  assign n60867 = n59352 & n60858;
  assign n60868 = ~n60866 & ~n60867;
  assign n60869 = ~n59286 & n59327;
  assign n60870 = n60868 & ~n60869;
  assign n60871 = ~n60844 & ~n60870;
  assign n60872 = P2_P3_INSTQUEUERD_ADDR_REG_1_ & n60844;
  assign n11006 = n60871 | n60872;
  assign n60874 = P2_P3_STATE2_REG_1_ & n59343;
  assign n60875 = ~P2_P3_INSTQUEUERD_ADDR_REG_0_ & n59336;
  assign n60876 = ~n60874 & ~n60875;
  assign n60877 = ~n59272 & n59327;
  assign n60878 = n60876 & ~n60877;
  assign n60879 = ~n60844 & ~n60878;
  assign n60880 = P2_P3_INSTQUEUERD_ADDR_REG_0_ & n60844;
  assign n11011 = n60879 | n60880;
  assign n60882 = P2_P3_STATE2_REG_0_ & n58679;
  assign n60883 = ~n59366 & n60882;
  assign n60884 = ~n59384 & ~n60841;
  assign n60885 = ~n60883 & n60884;
  assign n11016 = P2_P3_INSTQUEUEWR_ADDR_REG_4_ & n60885;
  assign n60887 = P2_P3_STATE2_REG_3_ & ~n59378;
  assign n60888 = ~n60885 & ~n60887;
  assign n60889 = P2_P3_INSTQUEUEWR_ADDR_REG_3_ & ~n60888;
  assign n60890 = ~n59327 & ~n59400;
  assign n60891 = ~n59420 & ~n60890;
  assign n60892 = P2_P3_STATE2_REG_3_ & n59389;
  assign n60893 = ~n60891 & ~n60892;
  assign n60894 = n59408 & ~n59415;
  assign n60895 = ~n59426 & ~n60894;
  assign n60896 = ~n60161 & ~n60895;
  assign n60897 = n59436 & ~n60896;
  assign n60898 = n60893 & ~n60897;
  assign n60899 = ~n60885 & ~n60898;
  assign n11021 = n60889 | n60899;
  assign n60901 = ~n59411 & ~n60890;
  assign n60902 = P2_P3_STATE2_REG_3_ & ~P2_P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n60903 = n59377 & n60902;
  assign n60904 = ~n60901 & ~n60903;
  assign n60905 = ~n59408 & ~n59415;
  assign n60906 = n59408 & n59415;
  assign n60907 = ~n60905 & ~n60906;
  assign n60908 = n59436 & ~n60907;
  assign n60909 = n60904 & ~n60908;
  assign n60910 = ~n60885 & ~n60909;
  assign n60911 = P2_P3_STATE2_REG_3_ & ~n59377;
  assign n60912 = ~n60885 & ~n60911;
  assign n60913 = P2_P3_INSTQUEUEWR_ADDR_REG_2_ & ~n60912;
  assign n11026 = n60910 | n60913;
  assign n60915 = ~n59404 & ~n60890;
  assign n60916 = P2_P3_STATE2_REG_3_ & ~P2_P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n60917 = ~n59407 & n59436;
  assign n60918 = ~n60916 & ~n60917;
  assign n60919 = P2_P3_INSTQUEUEWR_ADDR_REG_0_ & ~n60918;
  assign n60920 = n59436 & n59640;
  assign n60921 = ~n60915 & ~n60919;
  assign n60922 = ~n60920 & n60921;
  assign n60923 = ~n60885 & ~n60922;
  assign n60924 = P2_P3_STATE2_REG_3_ & ~P2_P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n60925 = ~n60885 & ~n60924;
  assign n60926 = P2_P3_INSTQUEUEWR_ADDR_REG_1_ & ~n60925;
  assign n11031 = n60923 | n60926;
  assign n60928 = ~n59327 & ~n59399;
  assign n60929 = ~n60885 & n60928;
  assign n60930 = P2_P3_INSTQUEUEWR_ADDR_REG_0_ & ~n60929;
  assign n60931 = ~n59367 & ~n60924;
  assign n60932 = ~n60885 & ~n60931;
  assign n11036 = n60930 | n60932;
  assign n60934 = ~P2_P3_STATE2_REG_1_ & n59399;
  assign n60935 = ~P2_P3_STATE2_REG_0_ & n60934;
  assign n60936 = n58975 & n59019;
  assign n60937 = ~n58807 & ~n58966;
  assign n60938 = n59064 & n60937;
  assign n60939 = n58973 & n59019;
  assign n60940 = ~n59203 & ~n60938;
  assign n60941 = ~n60939 & n60940;
  assign n60942 = n59024 & n59072;
  assign n60943 = n58776 & n58971;
  assign n60944 = n59019 & n60943;
  assign n60945 = ~n60942 & ~n60944;
  assign n60946 = n58935 & ~n60945;
  assign n60947 = ~n58775 & n59078;
  assign n60948 = ~n58594 & n58744;
  assign n60949 = n59019 & n60948;
  assign n60950 = ~n60947 & ~n60949;
  assign n60951 = ~n58935 & ~n60950;
  assign n60952 = n58966 & n59064;
  assign n60953 = ~n60946 & ~n60951;
  assign n60954 = ~n60952 & n60953;
  assign n60955 = n58900 & ~n60954;
  assign n60956 = n59195 & ~n60936;
  assign n60957 = n60941 & n60956;
  assign n60958 = ~n60955 & n60957;
  assign n60959 = n59321 & ~n60958;
  assign n60960 = ~n60935 & ~n60959;
  assign n60961 = P2_P3_STATE2_REG_2_ & ~n60960;
  assign n60962 = ~P2_P3_INSTADDRPOINTER_REG_0_ & n59265;
  assign n60963 = ~P2_P3_INSTADDRPOINTER_REG_0_ & n59108;
  assign n60964 = ~n60962 & ~n60963;
  assign n60965 = ~P2_P3_INSTADDRPOINTER_REG_0_ & ~n59155;
  assign n60966 = P2_P3_INSTADDRPOINTER_REG_0_ & n59226;
  assign n60967 = P2_P3_INSTADDRPOINTER_REG_0_ & n59227;
  assign n60968 = n58967 & n59098;
  assign n60969 = n59104 & n60968;
  assign n60970 = ~P2_P3_INSTADDRPOINTER_REG_0_ & n60969;
  assign n60971 = n59044 & n59098;
  assign n60972 = n59104 & n60971;
  assign n60973 = ~P2_P3_INSTADDRPOINTER_REG_0_ & n60972;
  assign n60974 = ~n60970 & ~n60973;
  assign n60975 = P2_P3_INSTADDRPOINTER_REG_0_ & n59042;
  assign n60976 = n60974 & ~n60975;
  assign n60977 = n59169 & n60851;
  assign n60978 = P2_P3_INSTQUEUERD_ADDR_REG_0_ & ~n59281;
  assign n60979 = n60977 & n60978;
  assign n60980 = P2_P3_INSTQUEUE_REG_0__0_ & n60979;
  assign n60981 = ~P2_P3_INSTQUEUERD_ADDR_REG_0_ & ~n59281;
  assign n60982 = n60977 & n60981;
  assign n60983 = P2_P3_INSTQUEUE_REG_1__0_ & n60982;
  assign n60984 = P2_P3_INSTQUEUERD_ADDR_REG_0_ & n59281;
  assign n60985 = n60977 & n60984;
  assign n60986 = P2_P3_INSTQUEUE_REG_2__0_ & n60985;
  assign n60987 = ~P2_P3_INSTQUEUERD_ADDR_REG_0_ & n59281;
  assign n60988 = n60977 & n60987;
  assign n60989 = P2_P3_INSTQUEUE_REG_3__0_ & n60988;
  assign n60990 = ~n60980 & ~n60983;
  assign n60991 = ~n60986 & n60990;
  assign n60992 = ~n60989 & n60991;
  assign n60993 = ~n59169 & n60851;
  assign n60994 = n60978 & n60993;
  assign n60995 = P2_P3_INSTQUEUE_REG_4__0_ & n60994;
  assign n60996 = n60981 & n60993;
  assign n60997 = P2_P3_INSTQUEUE_REG_5__0_ & n60996;
  assign n60998 = n60984 & n60993;
  assign n60999 = P2_P3_INSTQUEUE_REG_6__0_ & n60998;
  assign n61000 = n60987 & n60993;
  assign n61001 = P2_P3_INSTQUEUE_REG_7__0_ & n61000;
  assign n61002 = ~n60995 & ~n60997;
  assign n61003 = ~n60999 & n61002;
  assign n61004 = ~n61001 & n61003;
  assign n61005 = n59169 & ~n60851;
  assign n61006 = n60978 & n61005;
  assign n61007 = P2_P3_INSTQUEUE_REG_8__0_ & n61006;
  assign n61008 = n60981 & n61005;
  assign n61009 = P2_P3_INSTQUEUE_REG_9__0_ & n61008;
  assign n61010 = n60984 & n61005;
  assign n61011 = P2_P3_INSTQUEUE_REG_10__0_ & n61010;
  assign n61012 = n60987 & n61005;
  assign n61013 = P2_P3_INSTQUEUE_REG_11__0_ & n61012;
  assign n61014 = ~n61007 & ~n61009;
  assign n61015 = ~n61011 & n61014;
  assign n61016 = ~n61013 & n61015;
  assign n61017 = ~n59169 & ~n60851;
  assign n61018 = n60978 & n61017;
  assign n61019 = P2_P3_INSTQUEUE_REG_12__0_ & n61018;
  assign n61020 = n60981 & n61017;
  assign n61021 = P2_P3_INSTQUEUE_REG_13__0_ & n61020;
  assign n61022 = n60984 & n61017;
  assign n61023 = P2_P3_INSTQUEUE_REG_14__0_ & n61022;
  assign n61024 = n60987 & n61017;
  assign n61025 = P2_P3_INSTQUEUE_REG_15__0_ & n61024;
  assign n61026 = ~n61019 & ~n61021;
  assign n61027 = ~n61023 & n61026;
  assign n61028 = ~n61025 & n61027;
  assign n61029 = n60992 & n61004;
  assign n61030 = n61016 & n61029;
  assign n61031 = n61028 & n61030;
  assign n61032 = P2_P3_INSTADDRPOINTER_REG_0_ & n61031;
  assign n61033 = ~P2_P3_INSTADDRPOINTER_REG_0_ & ~n61031;
  assign n61034 = ~n61032 & ~n61033;
  assign n61035 = P2_P3_INSTQUEUE_REG_0__7_ & n60979;
  assign n61036 = P2_P3_INSTQUEUE_REG_1__7_ & n60982;
  assign n61037 = P2_P3_INSTQUEUE_REG_2__7_ & n60985;
  assign n61038 = P2_P3_INSTQUEUE_REG_3__7_ & n60988;
  assign n61039 = ~n61035 & ~n61036;
  assign n61040 = ~n61037 & n61039;
  assign n61041 = ~n61038 & n61040;
  assign n61042 = P2_P3_INSTQUEUE_REG_4__7_ & n60994;
  assign n61043 = P2_P3_INSTQUEUE_REG_5__7_ & n60996;
  assign n61044 = P2_P3_INSTQUEUE_REG_6__7_ & n60998;
  assign n61045 = P2_P3_INSTQUEUE_REG_7__7_ & n61000;
  assign n61046 = ~n61042 & ~n61043;
  assign n61047 = ~n61044 & n61046;
  assign n61048 = ~n61045 & n61047;
  assign n61049 = P2_P3_INSTQUEUE_REG_8__7_ & n61006;
  assign n61050 = P2_P3_INSTQUEUE_REG_9__7_ & n61008;
  assign n61051 = P2_P3_INSTQUEUE_REG_10__7_ & n61010;
  assign n61052 = P2_P3_INSTQUEUE_REG_11__7_ & n61012;
  assign n61053 = ~n61049 & ~n61050;
  assign n61054 = ~n61051 & n61053;
  assign n61055 = ~n61052 & n61054;
  assign n61056 = P2_P3_INSTQUEUE_REG_12__7_ & n61018;
  assign n61057 = P2_P3_INSTQUEUE_REG_13__7_ & n61020;
  assign n61058 = P2_P3_INSTQUEUE_REG_14__7_ & n61022;
  assign n61059 = P2_P3_INSTQUEUE_REG_15__7_ & n61024;
  assign n61060 = ~n61056 & ~n61057;
  assign n61061 = ~n61058 & n61060;
  assign n61062 = ~n61059 & n61061;
  assign n61063 = n61041 & n61048;
  assign n61064 = n61055 & n61063;
  assign n61065 = n61062 & n61064;
  assign n61066 = n59074 & ~n61065;
  assign n61067 = ~n61034 & n61066;
  assign n61068 = n59074 & n61065;
  assign n61069 = ~n61034 & n61068;
  assign n61070 = ~n60966 & ~n60967;
  assign n61071 = n60976 & n61070;
  assign n61072 = ~n61067 & n61071;
  assign n61073 = ~n61069 & n61072;
  assign n61074 = n59040 & n59068;
  assign n61075 = ~P2_P3_INSTADDRPOINTER_REG_0_ & n61074;
  assign n61076 = ~P2_P3_INSTADDRPOINTER_REG_0_ & n59112;
  assign n61077 = n58869 & n59055;
  assign n61078 = n59101 & n61077;
  assign n61079 = ~P2_P3_INSTADDRPOINTER_REG_0_ & n61078;
  assign n61080 = ~P2_P3_INSTADDRPOINTER_REG_0_ & n61031;
  assign n61081 = P2_P3_INSTADDRPOINTER_REG_0_ & ~n61031;
  assign n61082 = ~n61080 & ~n61081;
  assign n61083 = n59069 & ~n61082;
  assign n61084 = n58744 & n59098;
  assign n61085 = n59101 & n61084;
  assign n61086 = ~P2_P3_INSTADDRPOINTER_REG_0_ & n61085;
  assign n61087 = ~n61075 & ~n61076;
  assign n61088 = ~n61079 & n61087;
  assign n61089 = ~n61083 & n61088;
  assign n61090 = ~n61086 & n61089;
  assign n61091 = P2_P3_INSTADDRPOINTER_REG_0_ & n58968;
  assign n61092 = P2_P3_INSTADDRPOINTER_REG_0_ & n59046;
  assign n61093 = P2_P3_INSTADDRPOINTER_REG_0_ & n59050;
  assign n61094 = ~P2_P3_INSTADDRPOINTER_REG_0_ & n59066;
  assign n61095 = ~P2_P3_INSTADDRPOINTER_REG_0_ & n59058;
  assign n61096 = ~n61091 & ~n61092;
  assign n61097 = ~n61093 & n61096;
  assign n61098 = ~n61094 & n61097;
  assign n61099 = ~n61095 & n61098;
  assign n61100 = n61090 & n61099;
  assign n61101 = n60964 & ~n60965;
  assign n61102 = n61073 & n61101;
  assign n61103 = n61100 & n61102;
  assign n61104 = n60961 & ~n61103;
  assign n61105 = ~P2_P3_STATE2_REG_2_ & ~n60960;
  assign n61106 = P2_P3_REIP_REG_0_ & n61105;
  assign n61107 = P2_P3_INSTADDRPOINTER_REG_0_ & n60960;
  assign n61108 = ~n61104 & ~n61106;
  assign n11041 = n61107 | ~n61108;
  assign n61110 = P2_P3_INSTADDRPOINTER_REG_1_ & n60960;
  assign n61111 = P2_P3_REIP_REG_1_ & n61105;
  assign n61112 = ~n59155 & ~n59349;
  assign n61113 = n59265 & ~n59349;
  assign n61114 = n59108 & ~n59349;
  assign n61115 = ~n61113 & ~n61114;
  assign n61116 = ~P2_P3_INSTADDRPOINTER_REG_1_ & n61081;
  assign n61117 = P2_P3_INSTADDRPOINTER_REG_1_ & ~n61081;
  assign n61118 = ~n61116 & ~n61117;
  assign n61119 = P2_P3_INSTQUEUE_REG_0__1_ & n60979;
  assign n61120 = P2_P3_INSTQUEUE_REG_1__1_ & n60982;
  assign n61121 = P2_P3_INSTQUEUE_REG_2__1_ & n60985;
  assign n61122 = P2_P3_INSTQUEUE_REG_3__1_ & n60988;
  assign n61123 = ~n61119 & ~n61120;
  assign n61124 = ~n61121 & n61123;
  assign n61125 = ~n61122 & n61124;
  assign n61126 = P2_P3_INSTQUEUE_REG_4__1_ & n60994;
  assign n61127 = P2_P3_INSTQUEUE_REG_5__1_ & n60996;
  assign n61128 = P2_P3_INSTQUEUE_REG_6__1_ & n60998;
  assign n61129 = P2_P3_INSTQUEUE_REG_7__1_ & n61000;
  assign n61130 = ~n61126 & ~n61127;
  assign n61131 = ~n61128 & n61130;
  assign n61132 = ~n61129 & n61131;
  assign n61133 = P2_P3_INSTQUEUE_REG_8__1_ & n61006;
  assign n61134 = P2_P3_INSTQUEUE_REG_9__1_ & n61008;
  assign n61135 = P2_P3_INSTQUEUE_REG_10__1_ & n61010;
  assign n61136 = P2_P3_INSTQUEUE_REG_11__1_ & n61012;
  assign n61137 = ~n61133 & ~n61134;
  assign n61138 = ~n61135 & n61137;
  assign n61139 = ~n61136 & n61138;
  assign n61140 = P2_P3_INSTQUEUE_REG_12__1_ & n61018;
  assign n61141 = P2_P3_INSTQUEUE_REG_13__1_ & n61020;
  assign n61142 = P2_P3_INSTQUEUE_REG_14__1_ & n61022;
  assign n61143 = P2_P3_INSTQUEUE_REG_15__1_ & n61024;
  assign n61144 = ~n61140 & ~n61141;
  assign n61145 = ~n61142 & n61144;
  assign n61146 = ~n61143 & n61145;
  assign n61147 = n61125 & n61132;
  assign n61148 = n61139 & n61147;
  assign n61149 = n61146 & n61148;
  assign n61150 = ~n61118 & ~n61149;
  assign n61151 = ~P2_P3_INSTADDRPOINTER_REG_1_ & ~n61081;
  assign n61152 = n61149 & n61151;
  assign n61153 = n61081 & n61149;
  assign n61154 = P2_P3_INSTADDRPOINTER_REG_1_ & n61153;
  assign n61155 = ~n61150 & ~n61152;
  assign n61156 = ~n61154 & n61155;
  assign n61157 = n61068 & ~n61156;
  assign n61158 = ~n59349 & n61085;
  assign n61159 = ~n59349 & n61078;
  assign n61160 = ~n59349 & n61074;
  assign n61161 = n59112 & ~n59349;
  assign n61162 = ~n61158 & ~n61159;
  assign n61163 = ~n61160 & n61162;
  assign n61164 = ~n61161 & n61163;
  assign n61165 = ~P2_P3_INSTADDRPOINTER_REG_1_ & n58968;
  assign n61166 = ~P2_P3_INSTADDRPOINTER_REG_1_ & n59046;
  assign n61167 = ~P2_P3_INSTADDRPOINTER_REG_1_ & n59050;
  assign n61168 = n59066 & ~n59349;
  assign n61169 = n59058 & ~n59349;
  assign n61170 = ~n61165 & ~n61166;
  assign n61171 = ~n61167 & n61170;
  assign n61172 = ~n61168 & n61171;
  assign n61173 = ~n61169 & n61172;
  assign n61174 = ~P2_P3_INSTADDRPOINTER_REG_1_ & n61032;
  assign n61175 = P2_P3_INSTADDRPOINTER_REG_1_ & ~n61032;
  assign n61176 = ~n61174 & ~n61175;
  assign n61177 = ~n61031 & n61149;
  assign n61178 = n61031 & ~n61149;
  assign n61179 = ~n61177 & ~n61178;
  assign n61180 = ~n61176 & n61179;
  assign n61181 = ~P2_P3_INSTADDRPOINTER_REG_1_ & ~n61032;
  assign n61182 = ~n61179 & n61181;
  assign n61183 = n61032 & ~n61179;
  assign n61184 = P2_P3_INSTADDRPOINTER_REG_1_ & n61183;
  assign n61185 = ~n61180 & ~n61182;
  assign n61186 = ~n61184 & n61185;
  assign n61187 = n59069 & ~n61186;
  assign n61188 = n61164 & n61173;
  assign n61189 = ~n61187 & n61188;
  assign n61190 = ~P2_P3_INSTADDRPOINTER_REG_1_ & n59226;
  assign n61191 = ~P2_P3_INSTADDRPOINTER_REG_1_ & n59227;
  assign n61192 = ~n59349 & n60969;
  assign n61193 = ~n59349 & n60972;
  assign n61194 = ~n61192 & ~n61193;
  assign n61195 = ~P2_P3_INSTADDRPOINTER_REG_1_ & n59042;
  assign n61196 = n61194 & ~n61195;
  assign n61197 = n61081 & ~n61149;
  assign n61198 = ~n61081 & n61149;
  assign n61199 = ~n61197 & ~n61198;
  assign n61200 = ~P2_P3_INSTADDRPOINTER_REG_1_ & ~n61199;
  assign n61201 = ~n61081 & ~n61149;
  assign n61202 = P2_P3_INSTADDRPOINTER_REG_1_ & n61201;
  assign n61203 = P2_P3_INSTADDRPOINTER_REG_1_ & n61081;
  assign n61204 = n61149 & n61203;
  assign n61205 = ~n61200 & ~n61202;
  assign n61206 = ~n61204 & n61205;
  assign n61207 = n61066 & ~n61206;
  assign n61208 = ~n61190 & ~n61191;
  assign n61209 = n61196 & n61208;
  assign n61210 = ~n61207 & n61209;
  assign n61211 = ~n61112 & n61115;
  assign n61212 = ~n61157 & n61211;
  assign n61213 = n61189 & n61212;
  assign n61214 = n61210 & n61213;
  assign n61215 = n60961 & ~n61214;
  assign n61216 = ~n61110 & ~n61111;
  assign n11046 = n61215 | ~n61216;
  assign n61218 = P2_P3_INSTADDRPOINTER_REG_2_ & n60960;
  assign n61219 = P2_P3_REIP_REG_2_ & n61105;
  assign n61220 = P2_P3_INSTADDRPOINTER_REG_0_ & P2_P3_INSTADDRPOINTER_REG_1_;
  assign n61221 = ~P2_P3_INSTADDRPOINTER_REG_2_ & n61220;
  assign n61222 = P2_P3_INSTADDRPOINTER_REG_2_ & ~n61220;
  assign n61223 = ~n61221 & ~n61222;
  assign n61224 = ~n59155 & ~n61223;
  assign n61225 = P2_P3_INSTADDRPOINTER_REG_1_ & ~P2_P3_INSTADDRPOINTER_REG_2_;
  assign n61226 = ~P2_P3_INSTADDRPOINTER_REG_1_ & P2_P3_INSTADDRPOINTER_REG_2_;
  assign n61227 = ~n61225 & ~n61226;
  assign n61228 = n59226 & ~n61227;
  assign n61229 = n59227 & ~n61227;
  assign n61230 = n60969 & ~n61223;
  assign n61231 = n60972 & ~n61223;
  assign n61232 = ~n61230 & ~n61231;
  assign n61233 = n59042 & ~n61227;
  assign n61234 = n61232 & ~n61233;
  assign n61235 = ~n61228 & ~n61229;
  assign n61236 = n61234 & n61235;
  assign n61237 = P2_P3_INSTADDRPOINTER_REG_1_ & ~n61201;
  assign n61238 = ~n61153 & ~n61237;
  assign n61239 = P2_P3_INSTQUEUE_REG_0__2_ & n60979;
  assign n61240 = P2_P3_INSTQUEUE_REG_1__2_ & n60982;
  assign n61241 = P2_P3_INSTQUEUE_REG_2__2_ & n60985;
  assign n61242 = P2_P3_INSTQUEUE_REG_3__2_ & n60988;
  assign n61243 = ~n61239 & ~n61240;
  assign n61244 = ~n61241 & n61243;
  assign n61245 = ~n61242 & n61244;
  assign n61246 = P2_P3_INSTQUEUE_REG_4__2_ & n60994;
  assign n61247 = P2_P3_INSTQUEUE_REG_5__2_ & n60996;
  assign n61248 = P2_P3_INSTQUEUE_REG_6__2_ & n60998;
  assign n61249 = P2_P3_INSTQUEUE_REG_7__2_ & n61000;
  assign n61250 = ~n61246 & ~n61247;
  assign n61251 = ~n61248 & n61250;
  assign n61252 = ~n61249 & n61251;
  assign n61253 = P2_P3_INSTQUEUE_REG_8__2_ & n61006;
  assign n61254 = P2_P3_INSTQUEUE_REG_9__2_ & n61008;
  assign n61255 = P2_P3_INSTQUEUE_REG_10__2_ & n61010;
  assign n61256 = P2_P3_INSTQUEUE_REG_11__2_ & n61012;
  assign n61257 = ~n61253 & ~n61254;
  assign n61258 = ~n61255 & n61257;
  assign n61259 = ~n61256 & n61258;
  assign n61260 = P2_P3_INSTQUEUE_REG_12__2_ & n61018;
  assign n61261 = P2_P3_INSTQUEUE_REG_13__2_ & n61020;
  assign n61262 = P2_P3_INSTQUEUE_REG_14__2_ & n61022;
  assign n61263 = P2_P3_INSTQUEUE_REG_15__2_ & n61024;
  assign n61264 = ~n61260 & ~n61261;
  assign n61265 = ~n61262 & n61264;
  assign n61266 = ~n61263 & n61265;
  assign n61267 = n61245 & n61252;
  assign n61268 = n61259 & n61267;
  assign n61269 = n61266 & n61268;
  assign n61270 = ~n61149 & n61269;
  assign n61271 = n61149 & ~n61269;
  assign n61272 = ~n61270 & ~n61271;
  assign n61273 = ~P2_P3_INSTADDRPOINTER_REG_2_ & ~n61272;
  assign n61274 = P2_P3_INSTADDRPOINTER_REG_2_ & n61272;
  assign n61275 = ~n61273 & ~n61274;
  assign n61276 = n61238 & ~n61275;
  assign n61277 = ~n61238 & n61275;
  assign n61278 = ~n61276 & ~n61277;
  assign n61279 = n61068 & ~n61278;
  assign n61280 = n59265 & ~n61223;
  assign n61281 = n59108 & ~n61223;
  assign n61282 = ~n61280 & ~n61281;
  assign n61283 = P2_P3_INSTADDRPOINTER_REG_1_ & n61149;
  assign n61284 = ~n61153 & ~n61203;
  assign n61285 = ~n61283 & n61284;
  assign n61286 = ~n61275 & n61285;
  assign n61287 = ~P2_P3_INSTADDRPOINTER_REG_2_ & n61272;
  assign n61288 = P2_P3_INSTADDRPOINTER_REG_2_ & ~n61272;
  assign n61289 = ~n61287 & ~n61288;
  assign n61290 = ~n61285 & ~n61289;
  assign n61291 = ~n61286 & ~n61290;
  assign n61292 = n61066 & ~n61291;
  assign n61293 = n61282 & ~n61292;
  assign n61294 = n61085 & ~n61223;
  assign n61295 = n61078 & ~n61223;
  assign n61296 = n61074 & ~n61223;
  assign n61297 = n59112 & ~n61223;
  assign n61298 = ~n61294 & ~n61295;
  assign n61299 = ~n61296 & n61298;
  assign n61300 = ~n61297 & n61299;
  assign n61301 = n58968 & ~n61227;
  assign n61302 = n59046 & ~n61227;
  assign n61303 = n59050 & ~n61227;
  assign n61304 = ~P2_P3_INSTADDRPOINTER_REG_2_ & ~n61220;
  assign n61305 = P2_P3_INSTADDRPOINTER_REG_2_ & n61220;
  assign n61306 = ~n61304 & ~n61305;
  assign n61307 = n59066 & ~n61306;
  assign n61308 = n59058 & ~n61306;
  assign n61309 = ~n61301 & ~n61302;
  assign n61310 = ~n61303 & n61309;
  assign n61311 = ~n61307 & n61310;
  assign n61312 = ~n61308 & n61311;
  assign n61313 = ~n61031 & ~n61149;
  assign n61314 = n61269 & ~n61313;
  assign n61315 = ~n61269 & n61313;
  assign n61316 = ~n61314 & ~n61315;
  assign n61317 = ~P2_P3_INSTADDRPOINTER_REG_2_ & ~n61316;
  assign n61318 = P2_P3_INSTADDRPOINTER_REG_2_ & n61316;
  assign n61319 = ~n61317 & ~n61318;
  assign n61320 = ~n61032 & n61179;
  assign n61321 = P2_P3_INSTADDRPOINTER_REG_1_ & ~n61320;
  assign n61322 = ~n61183 & ~n61321;
  assign n61323 = ~n61319 & n61322;
  assign n61324 = ~P2_P3_INSTADDRPOINTER_REG_2_ & n61316;
  assign n61325 = P2_P3_INSTADDRPOINTER_REG_2_ & ~n61316;
  assign n61326 = ~n61324 & ~n61325;
  assign n61327 = ~n61322 & ~n61326;
  assign n61328 = ~n61323 & ~n61327;
  assign n61329 = n59069 & ~n61328;
  assign n61330 = n61300 & n61312;
  assign n61331 = ~n61329 & n61330;
  assign n61332 = ~n61224 & n61236;
  assign n61333 = ~n61279 & n61332;
  assign n61334 = n61293 & n61333;
  assign n61335 = n61331 & n61334;
  assign n61336 = n60961 & ~n61335;
  assign n61337 = ~n61218 & ~n61219;
  assign n11051 = n61336 | ~n61337;
  assign n61339 = P2_P3_INSTADDRPOINTER_REG_3_ & n60960;
  assign n61340 = P2_P3_REIP_REG_3_ & n61105;
  assign n61341 = ~P2_P3_INSTADDRPOINTER_REG_3_ & n61305;
  assign n61342 = P2_P3_INSTADDRPOINTER_REG_3_ & ~n61305;
  assign n61343 = ~n61341 & ~n61342;
  assign n61344 = n59265 & ~n61343;
  assign n61345 = n59108 & ~n61343;
  assign n61346 = ~n61344 & ~n61345;
  assign n61347 = ~n59155 & ~n61343;
  assign n61348 = P2_P3_INSTADDRPOINTER_REG_1_ & P2_P3_INSTADDRPOINTER_REG_2_;
  assign n61349 = ~P2_P3_INSTADDRPOINTER_REG_3_ & n61348;
  assign n61350 = P2_P3_INSTADDRPOINTER_REG_3_ & ~n61348;
  assign n61351 = ~n61349 & ~n61350;
  assign n61352 = n59226 & ~n61351;
  assign n61353 = n59227 & ~n61351;
  assign n61354 = n60969 & ~n61343;
  assign n61355 = n60972 & ~n61343;
  assign n61356 = ~n61354 & ~n61355;
  assign n61357 = n59042 & ~n61351;
  assign n61358 = n61356 & ~n61357;
  assign n61359 = ~n61352 & ~n61353;
  assign n61360 = n61358 & n61359;
  assign n61361 = ~n61285 & ~n61287;
  assign n61362 = ~n61288 & ~n61361;
  assign n61363 = P2_P3_INSTQUEUE_REG_0__3_ & n60979;
  assign n61364 = P2_P3_INSTQUEUE_REG_1__3_ & n60982;
  assign n61365 = P2_P3_INSTQUEUE_REG_2__3_ & n60985;
  assign n61366 = P2_P3_INSTQUEUE_REG_3__3_ & n60988;
  assign n61367 = ~n61363 & ~n61364;
  assign n61368 = ~n61365 & n61367;
  assign n61369 = ~n61366 & n61368;
  assign n61370 = P2_P3_INSTQUEUE_REG_4__3_ & n60994;
  assign n61371 = P2_P3_INSTQUEUE_REG_5__3_ & n60996;
  assign n61372 = P2_P3_INSTQUEUE_REG_6__3_ & n60998;
  assign n61373 = P2_P3_INSTQUEUE_REG_7__3_ & n61000;
  assign n61374 = ~n61370 & ~n61371;
  assign n61375 = ~n61372 & n61374;
  assign n61376 = ~n61373 & n61375;
  assign n61377 = P2_P3_INSTQUEUE_REG_8__3_ & n61006;
  assign n61378 = P2_P3_INSTQUEUE_REG_9__3_ & n61008;
  assign n61379 = P2_P3_INSTQUEUE_REG_10__3_ & n61010;
  assign n61380 = P2_P3_INSTQUEUE_REG_11__3_ & n61012;
  assign n61381 = ~n61377 & ~n61378;
  assign n61382 = ~n61379 & n61381;
  assign n61383 = ~n61380 & n61382;
  assign n61384 = P2_P3_INSTQUEUE_REG_12__3_ & n61018;
  assign n61385 = P2_P3_INSTQUEUE_REG_13__3_ & n61020;
  assign n61386 = P2_P3_INSTQUEUE_REG_14__3_ & n61022;
  assign n61387 = P2_P3_INSTQUEUE_REG_15__3_ & n61024;
  assign n61388 = ~n61384 & ~n61385;
  assign n61389 = ~n61386 & n61388;
  assign n61390 = ~n61387 & n61389;
  assign n61391 = n61369 & n61376;
  assign n61392 = n61383 & n61391;
  assign n61393 = n61390 & n61392;
  assign n61394 = ~n61149 & ~n61269;
  assign n61395 = n61393 & ~n61394;
  assign n61396 = ~n61393 & n61394;
  assign n61397 = ~n61395 & ~n61396;
  assign n61398 = P2_P3_INSTADDRPOINTER_REG_3_ & ~n61397;
  assign n61399 = ~P2_P3_INSTADDRPOINTER_REG_3_ & n61397;
  assign n61400 = ~n61398 & ~n61399;
  assign n61401 = n61362 & ~n61400;
  assign n61402 = P2_P3_INSTADDRPOINTER_REG_3_ & n61397;
  assign n61403 = ~P2_P3_INSTADDRPOINTER_REG_3_ & ~n61397;
  assign n61404 = ~n61402 & ~n61403;
  assign n61405 = ~n61362 & ~n61404;
  assign n61406 = ~n61401 & ~n61405;
  assign n61407 = n61066 & ~n61406;
  assign n61408 = ~n61238 & ~n61287;
  assign n61409 = ~n61288 & ~n61408;
  assign n61410 = n61393 & n61394;
  assign n61411 = ~n61393 & ~n61394;
  assign n61412 = ~n61410 & ~n61411;
  assign n61413 = ~P2_P3_INSTADDRPOINTER_REG_3_ & n61412;
  assign n61414 = ~n61409 & ~n61413;
  assign n61415 = P2_P3_INSTADDRPOINTER_REG_3_ & ~n61412;
  assign n61416 = n61414 & ~n61415;
  assign n61417 = ~P2_P3_INSTADDRPOINTER_REG_3_ & ~n61412;
  assign n61418 = P2_P3_INSTADDRPOINTER_REG_3_ & n61412;
  assign n61419 = ~n61417 & ~n61418;
  assign n61420 = n61409 & n61419;
  assign n61421 = ~n61416 & ~n61420;
  assign n61422 = n61068 & n61421;
  assign n61423 = ~n61407 & ~n61422;
  assign n61424 = n61085 & ~n61343;
  assign n61425 = n61078 & ~n61343;
  assign n61426 = n61074 & ~n61343;
  assign n61427 = n59112 & ~n61343;
  assign n61428 = ~n61424 & ~n61425;
  assign n61429 = ~n61426 & n61428;
  assign n61430 = ~n61427 & n61429;
  assign n61431 = n58968 & ~n61351;
  assign n61432 = n59046 & ~n61351;
  assign n61433 = n59050 & ~n61351;
  assign n61434 = ~P2_P3_INSTADDRPOINTER_REG_3_ & n61304;
  assign n61435 = P2_P3_INSTADDRPOINTER_REG_3_ & ~n61304;
  assign n61436 = ~n61434 & ~n61435;
  assign n61437 = n59066 & n61436;
  assign n61438 = n59058 & n61436;
  assign n61439 = ~n61431 & ~n61432;
  assign n61440 = ~n61433 & n61439;
  assign n61441 = ~n61437 & n61440;
  assign n61442 = ~n61438 & n61441;
  assign n61443 = n61322 & ~n61325;
  assign n61444 = n61314 & n61393;
  assign n61445 = ~n61314 & ~n61393;
  assign n61446 = ~n61444 & ~n61445;
  assign n61447 = P2_P3_INSTADDRPOINTER_REG_3_ & n61446;
  assign n61448 = ~n61324 & n61446;
  assign n61449 = P2_P3_INSTADDRPOINTER_REG_3_ & ~n61324;
  assign n61450 = ~n61448 & ~n61449;
  assign n61451 = ~n61443 & ~n61447;
  assign n61452 = ~n61450 & n61451;
  assign n61453 = ~P2_P3_INSTADDRPOINTER_REG_3_ & n61446;
  assign n61454 = P2_P3_INSTADDRPOINTER_REG_3_ & ~n61446;
  assign n61455 = ~n61453 & ~n61454;
  assign n61456 = ~n61325 & n61455;
  assign n61457 = ~n61322 & ~n61324;
  assign n61458 = n61456 & ~n61457;
  assign n61459 = ~n61452 & ~n61458;
  assign n61460 = n59069 & n61459;
  assign n61461 = n61430 & n61442;
  assign n61462 = ~n61460 & n61461;
  assign n61463 = n61346 & ~n61347;
  assign n61464 = n61360 & n61463;
  assign n61465 = n61423 & n61464;
  assign n61466 = n61462 & n61465;
  assign n61467 = n60961 & ~n61466;
  assign n61468 = ~n61339 & ~n61340;
  assign n11056 = n61467 | ~n61468;
  assign n61470 = P2_P3_INSTADDRPOINTER_REG_4_ & n60960;
  assign n61471 = P2_P3_REIP_REG_4_ & n61105;
  assign n61472 = P2_P3_INSTADDRPOINTER_REG_3_ & n61305;
  assign n61473 = ~P2_P3_INSTADDRPOINTER_REG_4_ & n61472;
  assign n61474 = P2_P3_INSTADDRPOINTER_REG_4_ & ~n61472;
  assign n61475 = ~n61473 & ~n61474;
  assign n61476 = ~n59155 & ~n61475;
  assign n61477 = P2_P3_INSTADDRPOINTER_REG_3_ & n61348;
  assign n61478 = ~P2_P3_INSTADDRPOINTER_REG_4_ & n61477;
  assign n61479 = P2_P3_INSTADDRPOINTER_REG_4_ & ~n61477;
  assign n61480 = ~n61478 & ~n61479;
  assign n61481 = n59226 & ~n61480;
  assign n61482 = n59227 & ~n61480;
  assign n61483 = n60969 & ~n61475;
  assign n61484 = n60972 & ~n61475;
  assign n61485 = ~n61483 & ~n61484;
  assign n61486 = n59042 & ~n61480;
  assign n61487 = n61485 & ~n61486;
  assign n61488 = ~n61481 & ~n61482;
  assign n61489 = n61487 & n61488;
  assign n61490 = P2_P3_INSTQUEUE_REG_0__4_ & n60979;
  assign n61491 = P2_P3_INSTQUEUE_REG_1__4_ & n60982;
  assign n61492 = P2_P3_INSTQUEUE_REG_2__4_ & n60985;
  assign n61493 = P2_P3_INSTQUEUE_REG_3__4_ & n60988;
  assign n61494 = ~n61490 & ~n61491;
  assign n61495 = ~n61492 & n61494;
  assign n61496 = ~n61493 & n61495;
  assign n61497 = P2_P3_INSTQUEUE_REG_4__4_ & n60994;
  assign n61498 = P2_P3_INSTQUEUE_REG_5__4_ & n60996;
  assign n61499 = P2_P3_INSTQUEUE_REG_6__4_ & n60998;
  assign n61500 = P2_P3_INSTQUEUE_REG_7__4_ & n61000;
  assign n61501 = ~n61497 & ~n61498;
  assign n61502 = ~n61499 & n61501;
  assign n61503 = ~n61500 & n61502;
  assign n61504 = P2_P3_INSTQUEUE_REG_8__4_ & n61006;
  assign n61505 = P2_P3_INSTQUEUE_REG_9__4_ & n61008;
  assign n61506 = P2_P3_INSTQUEUE_REG_10__4_ & n61010;
  assign n61507 = P2_P3_INSTQUEUE_REG_11__4_ & n61012;
  assign n61508 = ~n61504 & ~n61505;
  assign n61509 = ~n61506 & n61508;
  assign n61510 = ~n61507 & n61509;
  assign n61511 = P2_P3_INSTQUEUE_REG_12__4_ & n61018;
  assign n61512 = P2_P3_INSTQUEUE_REG_13__4_ & n61020;
  assign n61513 = P2_P3_INSTQUEUE_REG_14__4_ & n61022;
  assign n61514 = P2_P3_INSTQUEUE_REG_15__4_ & n61024;
  assign n61515 = ~n61511 & ~n61512;
  assign n61516 = ~n61513 & n61515;
  assign n61517 = ~n61514 & n61516;
  assign n61518 = n61496 & n61503;
  assign n61519 = n61510 & n61518;
  assign n61520 = n61517 & n61519;
  assign n61521 = n61396 & n61520;
  assign n61522 = ~n61396 & ~n61520;
  assign n61523 = ~n61521 & ~n61522;
  assign n61524 = P2_P3_INSTADDRPOINTER_REG_4_ & ~n61523;
  assign n61525 = ~P2_P3_INSTADDRPOINTER_REG_4_ & n61523;
  assign n61526 = ~n61524 & ~n61525;
  assign n61527 = ~n61414 & ~n61415;
  assign n61528 = n61526 & ~n61527;
  assign n61529 = ~P2_P3_INSTADDRPOINTER_REG_4_ & ~n61523;
  assign n61530 = P2_P3_INSTADDRPOINTER_REG_4_ & n61523;
  assign n61531 = ~n61529 & ~n61530;
  assign n61532 = ~n61415 & n61531;
  assign n61533 = ~n61414 & n61532;
  assign n61534 = ~n61528 & ~n61533;
  assign n61535 = n61068 & n61534;
  assign n61536 = n59265 & ~n61475;
  assign n61537 = n59108 & ~n61475;
  assign n61538 = ~n61536 & ~n61537;
  assign n61539 = ~n61287 & ~n61403;
  assign n61540 = ~n61153 & ~n61283;
  assign n61541 = ~n61288 & n61540;
  assign n61542 = ~n61203 & n61541;
  assign n61543 = n61539 & ~n61542;
  assign n61544 = ~n61402 & ~n61543;
  assign n61545 = n61396 & ~n61520;
  assign n61546 = ~n61396 & n61520;
  assign n61547 = ~n61545 & ~n61546;
  assign n61548 = P2_P3_INSTADDRPOINTER_REG_4_ & ~n61547;
  assign n61549 = ~P2_P3_INSTADDRPOINTER_REG_4_ & n61547;
  assign n61550 = ~n61548 & ~n61549;
  assign n61551 = n61544 & ~n61550;
  assign n61552 = P2_P3_INSTADDRPOINTER_REG_4_ & n61547;
  assign n61553 = ~P2_P3_INSTADDRPOINTER_REG_4_ & ~n61547;
  assign n61554 = ~n61552 & ~n61553;
  assign n61555 = ~n61544 & ~n61554;
  assign n61556 = ~n61551 & ~n61555;
  assign n61557 = n61066 & ~n61556;
  assign n61558 = n61538 & ~n61557;
  assign n61559 = n61085 & ~n61475;
  assign n61560 = n61078 & ~n61475;
  assign n61561 = n61074 & ~n61475;
  assign n61562 = n59112 & ~n61475;
  assign n61563 = ~n61559 & ~n61560;
  assign n61564 = ~n61561 & n61563;
  assign n61565 = ~n61562 & n61564;
  assign n61566 = n58968 & ~n61480;
  assign n61567 = n59046 & ~n61480;
  assign n61568 = n59050 & ~n61480;
  assign n61569 = ~P2_P3_INSTADDRPOINTER_REG_4_ & n61435;
  assign n61570 = P2_P3_INSTADDRPOINTER_REG_4_ & ~n61435;
  assign n61571 = ~n61569 & ~n61570;
  assign n61572 = n59066 & ~n61571;
  assign n61573 = n59058 & ~n61571;
  assign n61574 = ~n61566 & ~n61567;
  assign n61575 = ~n61568 & n61574;
  assign n61576 = ~n61572 & n61575;
  assign n61577 = ~n61573 & n61576;
  assign n61578 = n61445 & n61520;
  assign n61579 = ~n61445 & ~n61520;
  assign n61580 = ~n61578 & ~n61579;
  assign n61581 = ~P2_P3_INSTADDRPOINTER_REG_4_ & ~n61580;
  assign n61582 = P2_P3_INSTADDRPOINTER_REG_4_ & n61580;
  assign n61583 = ~n61581 & ~n61582;
  assign n61584 = n61325 & n61446;
  assign n61585 = ~n61325 & ~n61446;
  assign n61586 = P2_P3_INSTADDRPOINTER_REG_3_ & ~n61585;
  assign n61587 = ~n61584 & ~n61586;
  assign n61588 = ~n61322 & ~n61450;
  assign n61589 = n61587 & ~n61588;
  assign n61590 = ~n61583 & n61589;
  assign n61591 = ~P2_P3_INSTADDRPOINTER_REG_4_ & n61580;
  assign n61592 = P2_P3_INSTADDRPOINTER_REG_4_ & ~n61580;
  assign n61593 = ~n61591 & ~n61592;
  assign n61594 = ~n61589 & ~n61593;
  assign n61595 = ~n61590 & ~n61594;
  assign n61596 = n59069 & ~n61595;
  assign n61597 = n61565 & n61577;
  assign n61598 = ~n61596 & n61597;
  assign n61599 = ~n61476 & n61489;
  assign n61600 = ~n61535 & n61599;
  assign n61601 = n61558 & n61600;
  assign n61602 = n61598 & n61601;
  assign n61603 = n60961 & ~n61602;
  assign n61604 = ~n61470 & ~n61471;
  assign n11061 = n61603 | ~n61604;
  assign n61606 = P2_P3_INSTADDRPOINTER_REG_5_ & n60960;
  assign n61607 = P2_P3_REIP_REG_5_ & n61105;
  assign n61608 = P2_P3_INSTADDRPOINTER_REG_4_ & n61477;
  assign n61609 = ~P2_P3_INSTADDRPOINTER_REG_5_ & n61608;
  assign n61610 = P2_P3_INSTADDRPOINTER_REG_5_ & ~n61608;
  assign n61611 = ~n61609 & ~n61610;
  assign n61612 = n59226 & ~n61611;
  assign n61613 = n59227 & ~n61611;
  assign n61614 = P2_P3_INSTADDRPOINTER_REG_4_ & n61472;
  assign n61615 = ~P2_P3_INSTADDRPOINTER_REG_5_ & n61614;
  assign n61616 = P2_P3_INSTADDRPOINTER_REG_5_ & ~n61614;
  assign n61617 = ~n61615 & ~n61616;
  assign n61618 = n60969 & ~n61617;
  assign n61619 = n60972 & ~n61617;
  assign n61620 = ~n61618 & ~n61619;
  assign n61621 = n59042 & ~n61611;
  assign n61622 = n61620 & ~n61621;
  assign n61623 = ~n61612 & ~n61613;
  assign n61624 = n61622 & n61623;
  assign n61625 = ~n59155 & ~n61617;
  assign n61626 = n61402 & ~n61553;
  assign n61627 = ~n61552 & ~n61626;
  assign n61628 = n61539 & ~n61553;
  assign n61629 = ~n61542 & n61628;
  assign n61630 = n61627 & ~n61629;
  assign n61631 = P2_P3_INSTQUEUE_REG_0__5_ & n60979;
  assign n61632 = P2_P3_INSTQUEUE_REG_1__5_ & n60982;
  assign n61633 = P2_P3_INSTQUEUE_REG_2__5_ & n60985;
  assign n61634 = P2_P3_INSTQUEUE_REG_3__5_ & n60988;
  assign n61635 = ~n61631 & ~n61632;
  assign n61636 = ~n61633 & n61635;
  assign n61637 = ~n61634 & n61636;
  assign n61638 = P2_P3_INSTQUEUE_REG_4__5_ & n60994;
  assign n61639 = P2_P3_INSTQUEUE_REG_5__5_ & n60996;
  assign n61640 = P2_P3_INSTQUEUE_REG_6__5_ & n60998;
  assign n61641 = P2_P3_INSTQUEUE_REG_7__5_ & n61000;
  assign n61642 = ~n61638 & ~n61639;
  assign n61643 = ~n61640 & n61642;
  assign n61644 = ~n61641 & n61643;
  assign n61645 = P2_P3_INSTQUEUE_REG_8__5_ & n61006;
  assign n61646 = P2_P3_INSTQUEUE_REG_9__5_ & n61008;
  assign n61647 = P2_P3_INSTQUEUE_REG_10__5_ & n61010;
  assign n61648 = P2_P3_INSTQUEUE_REG_11__5_ & n61012;
  assign n61649 = ~n61645 & ~n61646;
  assign n61650 = ~n61647 & n61649;
  assign n61651 = ~n61648 & n61650;
  assign n61652 = P2_P3_INSTQUEUE_REG_12__5_ & n61018;
  assign n61653 = P2_P3_INSTQUEUE_REG_13__5_ & n61020;
  assign n61654 = P2_P3_INSTQUEUE_REG_14__5_ & n61022;
  assign n61655 = P2_P3_INSTQUEUE_REG_15__5_ & n61024;
  assign n61656 = ~n61652 & ~n61653;
  assign n61657 = ~n61654 & n61656;
  assign n61658 = ~n61655 & n61657;
  assign n61659 = n61637 & n61644;
  assign n61660 = n61651 & n61659;
  assign n61661 = n61658 & n61660;
  assign n61662 = ~n61545 & n61661;
  assign n61663 = ~n61520 & ~n61661;
  assign n61664 = n61396 & n61663;
  assign n61665 = ~n61662 & ~n61664;
  assign n61666 = P2_P3_INSTADDRPOINTER_REG_5_ & ~n61665;
  assign n61667 = ~P2_P3_INSTADDRPOINTER_REG_5_ & n61665;
  assign n61668 = ~n61666 & ~n61667;
  assign n61669 = n61630 & ~n61668;
  assign n61670 = ~n61630 & n61668;
  assign n61671 = ~n61669 & ~n61670;
  assign n61672 = n61066 & ~n61671;
  assign n61673 = n59265 & ~n61617;
  assign n61674 = n59108 & ~n61617;
  assign n61675 = ~n61673 & ~n61674;
  assign n61676 = n61415 & ~n61525;
  assign n61677 = ~n61524 & ~n61676;
  assign n61678 = ~n61413 & ~n61525;
  assign n61679 = ~n61409 & n61678;
  assign n61680 = n61677 & ~n61679;
  assign n61681 = n61545 & n61661;
  assign n61682 = ~n61545 & ~n61661;
  assign n61683 = ~n61681 & ~n61682;
  assign n61684 = ~P2_P3_INSTADDRPOINTER_REG_5_ & ~n61683;
  assign n61685 = P2_P3_INSTADDRPOINTER_REG_5_ & n61683;
  assign n61686 = ~n61684 & ~n61685;
  assign n61687 = n61680 & ~n61686;
  assign n61688 = ~n61680 & n61686;
  assign n61689 = ~n61687 & ~n61688;
  assign n61690 = n61068 & ~n61689;
  assign n61691 = n61675 & ~n61690;
  assign n61692 = n61085 & ~n61617;
  assign n61693 = n61078 & ~n61617;
  assign n61694 = n61074 & ~n61617;
  assign n61695 = n59112 & ~n61617;
  assign n61696 = ~n61692 & ~n61693;
  assign n61697 = ~n61694 & n61696;
  assign n61698 = ~n61695 & n61697;
  assign n61699 = n58968 & ~n61611;
  assign n61700 = n59046 & ~n61611;
  assign n61701 = n59050 & ~n61611;
  assign n61702 = P2_P3_INSTADDRPOINTER_REG_4_ & n61435;
  assign n61703 = ~P2_P3_INSTADDRPOINTER_REG_5_ & n61702;
  assign n61704 = P2_P3_INSTADDRPOINTER_REG_5_ & ~n61702;
  assign n61705 = ~n61703 & ~n61704;
  assign n61706 = n59066 & ~n61705;
  assign n61707 = n59058 & ~n61705;
  assign n61708 = ~n61699 & ~n61700;
  assign n61709 = ~n61701 & n61708;
  assign n61710 = ~n61706 & n61709;
  assign n61711 = ~n61707 & n61710;
  assign n61712 = n61445 & ~n61520;
  assign n61713 = n61661 & n61712;
  assign n61714 = ~n61661 & ~n61712;
  assign n61715 = ~n61713 & ~n61714;
  assign n61716 = P2_P3_INSTADDRPOINTER_REG_5_ & ~n61715;
  assign n61717 = ~P2_P3_INSTADDRPOINTER_REG_5_ & n61715;
  assign n61718 = ~n61591 & ~n61717;
  assign n61719 = ~n61716 & n61718;
  assign n61720 = n61589 & ~n61592;
  assign n61721 = n61719 & ~n61720;
  assign n61722 = ~P2_P3_INSTADDRPOINTER_REG_5_ & ~n61715;
  assign n61723 = P2_P3_INSTADDRPOINTER_REG_5_ & n61715;
  assign n61724 = ~n61722 & ~n61723;
  assign n61725 = ~n61592 & n61724;
  assign n61726 = ~n61589 & ~n61591;
  assign n61727 = n61725 & ~n61726;
  assign n61728 = ~n61721 & ~n61727;
  assign n61729 = n59069 & n61728;
  assign n61730 = n61698 & n61711;
  assign n61731 = ~n61729 & n61730;
  assign n61732 = n61624 & ~n61625;
  assign n61733 = ~n61672 & n61732;
  assign n61734 = n61691 & n61733;
  assign n61735 = n61731 & n61734;
  assign n61736 = n60961 & ~n61735;
  assign n61737 = ~n61606 & ~n61607;
  assign n11066 = n61736 | ~n61737;
  assign n61739 = P2_P3_INSTADDRPOINTER_REG_6_ & n60960;
  assign n61740 = P2_P3_REIP_REG_6_ & n61105;
  assign n61741 = P2_P3_INSTADDRPOINTER_REG_5_ & n61608;
  assign n61742 = ~P2_P3_INSTADDRPOINTER_REG_6_ & n61741;
  assign n61743 = P2_P3_INSTADDRPOINTER_REG_6_ & ~n61741;
  assign n61744 = ~n61742 & ~n61743;
  assign n61745 = n59226 & ~n61744;
  assign n61746 = n59227 & ~n61744;
  assign n61747 = P2_P3_INSTADDRPOINTER_REG_5_ & n61614;
  assign n61748 = ~P2_P3_INSTADDRPOINTER_REG_6_ & n61747;
  assign n61749 = P2_P3_INSTADDRPOINTER_REG_6_ & ~n61747;
  assign n61750 = ~n61748 & ~n61749;
  assign n61751 = n60969 & ~n61750;
  assign n61752 = n60972 & ~n61750;
  assign n61753 = ~n61751 & ~n61752;
  assign n61754 = n59042 & ~n61744;
  assign n61755 = n61753 & ~n61754;
  assign n61756 = ~n61745 & ~n61746;
  assign n61757 = n61755 & n61756;
  assign n61758 = ~n59155 & ~n61750;
  assign n61759 = ~P2_P3_INSTADDRPOINTER_REG_5_ & ~n61665;
  assign n61760 = ~n61630 & ~n61759;
  assign n61761 = P2_P3_INSTADDRPOINTER_REG_5_ & n61665;
  assign n61762 = ~n61760 & ~n61761;
  assign n61763 = P2_P3_INSTQUEUE_REG_0__6_ & n60979;
  assign n61764 = P2_P3_INSTQUEUE_REG_1__6_ & n60982;
  assign n61765 = P2_P3_INSTQUEUE_REG_2__6_ & n60985;
  assign n61766 = P2_P3_INSTQUEUE_REG_3__6_ & n60988;
  assign n61767 = ~n61763 & ~n61764;
  assign n61768 = ~n61765 & n61767;
  assign n61769 = ~n61766 & n61768;
  assign n61770 = P2_P3_INSTQUEUE_REG_4__6_ & n60994;
  assign n61771 = P2_P3_INSTQUEUE_REG_5__6_ & n60996;
  assign n61772 = P2_P3_INSTQUEUE_REG_6__6_ & n60998;
  assign n61773 = P2_P3_INSTQUEUE_REG_7__6_ & n61000;
  assign n61774 = ~n61770 & ~n61771;
  assign n61775 = ~n61772 & n61774;
  assign n61776 = ~n61773 & n61775;
  assign n61777 = P2_P3_INSTQUEUE_REG_8__6_ & n61006;
  assign n61778 = P2_P3_INSTQUEUE_REG_9__6_ & n61008;
  assign n61779 = P2_P3_INSTQUEUE_REG_10__6_ & n61010;
  assign n61780 = P2_P3_INSTQUEUE_REG_11__6_ & n61012;
  assign n61781 = ~n61777 & ~n61778;
  assign n61782 = ~n61779 & n61781;
  assign n61783 = ~n61780 & n61782;
  assign n61784 = P2_P3_INSTQUEUE_REG_12__6_ & n61018;
  assign n61785 = P2_P3_INSTQUEUE_REG_13__6_ & n61020;
  assign n61786 = P2_P3_INSTQUEUE_REG_14__6_ & n61022;
  assign n61787 = P2_P3_INSTQUEUE_REG_15__6_ & n61024;
  assign n61788 = ~n61784 & ~n61785;
  assign n61789 = ~n61786 & n61788;
  assign n61790 = ~n61787 & n61789;
  assign n61791 = n61769 & n61776;
  assign n61792 = n61783 & n61791;
  assign n61793 = n61790 & n61792;
  assign n61794 = n61664 & ~n61793;
  assign n61795 = ~n61664 & n61793;
  assign n61796 = ~n61794 & ~n61795;
  assign n61797 = P2_P3_INSTADDRPOINTER_REG_6_ & ~n61796;
  assign n61798 = ~P2_P3_INSTADDRPOINTER_REG_6_ & n61796;
  assign n61799 = ~n61797 & ~n61798;
  assign n61800 = n61762 & ~n61799;
  assign n61801 = ~n61762 & n61799;
  assign n61802 = ~n61800 & ~n61801;
  assign n61803 = n61066 & ~n61802;
  assign n61804 = n59265 & ~n61750;
  assign n61805 = n59108 & ~n61750;
  assign n61806 = ~n61804 & ~n61805;
  assign n61807 = ~n61680 & ~n61683;
  assign n61808 = P2_P3_INSTADDRPOINTER_REG_5_ & ~n61680;
  assign n61809 = P2_P3_INSTADDRPOINTER_REG_5_ & ~n61683;
  assign n61810 = ~n61807 & ~n61808;
  assign n61811 = ~n61809 & n61810;
  assign n61812 = n61545 & ~n61661;
  assign n61813 = n61793 & n61812;
  assign n61814 = ~n61793 & ~n61812;
  assign n61815 = ~n61813 & ~n61814;
  assign n61816 = ~P2_P3_INSTADDRPOINTER_REG_6_ & ~n61815;
  assign n61817 = P2_P3_INSTADDRPOINTER_REG_6_ & n61815;
  assign n61818 = ~n61816 & ~n61817;
  assign n61819 = n61811 & ~n61818;
  assign n61820 = ~n61811 & n61818;
  assign n61821 = ~n61819 & ~n61820;
  assign n61822 = n61068 & ~n61821;
  assign n61823 = n61806 & ~n61822;
  assign n61824 = n61085 & ~n61750;
  assign n61825 = n61078 & ~n61750;
  assign n61826 = n61074 & ~n61750;
  assign n61827 = n59112 & ~n61750;
  assign n61828 = ~n61824 & ~n61825;
  assign n61829 = ~n61826 & n61828;
  assign n61830 = ~n61827 & n61829;
  assign n61831 = n58968 & ~n61744;
  assign n61832 = n59046 & ~n61744;
  assign n61833 = n59050 & ~n61744;
  assign n61834 = P2_P3_INSTADDRPOINTER_REG_5_ & n61702;
  assign n61835 = ~P2_P3_INSTADDRPOINTER_REG_6_ & n61834;
  assign n61836 = P2_P3_INSTADDRPOINTER_REG_6_ & ~n61834;
  assign n61837 = ~n61835 & ~n61836;
  assign n61838 = n59066 & ~n61837;
  assign n61839 = n59058 & ~n61837;
  assign n61840 = ~n61831 & ~n61832;
  assign n61841 = ~n61833 & n61840;
  assign n61842 = ~n61838 & n61841;
  assign n61843 = ~n61839 & n61842;
  assign n61844 = n61592 & ~n61715;
  assign n61845 = ~n61592 & n61715;
  assign n61846 = P2_P3_INSTADDRPOINTER_REG_5_ & ~n61845;
  assign n61847 = ~n61844 & ~n61846;
  assign n61848 = ~n61589 & n61718;
  assign n61849 = n61847 & ~n61848;
  assign n61850 = ~n61661 & n61712;
  assign n61851 = n61793 & n61850;
  assign n61852 = ~n61793 & ~n61850;
  assign n61853 = ~n61851 & ~n61852;
  assign n61854 = ~P2_P3_INSTADDRPOINTER_REG_6_ & ~n61853;
  assign n61855 = P2_P3_INSTADDRPOINTER_REG_6_ & n61853;
  assign n61856 = ~n61854 & ~n61855;
  assign n61857 = n61849 & ~n61856;
  assign n61858 = ~n61849 & n61856;
  assign n61859 = ~n61857 & ~n61858;
  assign n61860 = n59069 & ~n61859;
  assign n61861 = n61830 & n61843;
  assign n61862 = ~n61860 & n61861;
  assign n61863 = n61757 & ~n61758;
  assign n61864 = ~n61803 & n61863;
  assign n61865 = n61823 & n61864;
  assign n61866 = n61862 & n61865;
  assign n61867 = n60961 & ~n61866;
  assign n61868 = ~n61739 & ~n61740;
  assign n11071 = n61867 | ~n61868;
  assign n61870 = P2_P3_INSTADDRPOINTER_REG_7_ & n60960;
  assign n61871 = P2_P3_REIP_REG_7_ & n61105;
  assign n61872 = P2_P3_INSTADDRPOINTER_REG_6_ & n61741;
  assign n61873 = ~P2_P3_INSTADDRPOINTER_REG_7_ & n61872;
  assign n61874 = P2_P3_INSTADDRPOINTER_REG_7_ & ~n61872;
  assign n61875 = ~n61873 & ~n61874;
  assign n61876 = n59226 & ~n61875;
  assign n61877 = n59227 & ~n61875;
  assign n61878 = P2_P3_INSTADDRPOINTER_REG_6_ & n61747;
  assign n61879 = ~P2_P3_INSTADDRPOINTER_REG_7_ & n61878;
  assign n61880 = P2_P3_INSTADDRPOINTER_REG_7_ & ~n61878;
  assign n61881 = ~n61879 & ~n61880;
  assign n61882 = n60969 & ~n61881;
  assign n61883 = n60972 & ~n61881;
  assign n61884 = ~n61882 & ~n61883;
  assign n61885 = n59042 & ~n61875;
  assign n61886 = n61884 & ~n61885;
  assign n61887 = ~n61876 & ~n61877;
  assign n61888 = n61886 & n61887;
  assign n61889 = ~n59155 & ~n61881;
  assign n61890 = P2_P3_INSTADDRPOINTER_REG_6_ & n61796;
  assign n61891 = ~P2_P3_INSTADDRPOINTER_REG_6_ & ~n61796;
  assign n61892 = ~n61762 & ~n61891;
  assign n61893 = ~n61890 & ~n61892;
  assign n61894 = n61065 & ~n61794;
  assign n61895 = ~n61065 & ~n61793;
  assign n61896 = n61664 & n61895;
  assign n61897 = ~n61894 & ~n61896;
  assign n61898 = P2_P3_INSTADDRPOINTER_REG_7_ & ~n61897;
  assign n61899 = ~P2_P3_INSTADDRPOINTER_REG_7_ & n61897;
  assign n61900 = ~n61898 & ~n61899;
  assign n61901 = n61893 & ~n61900;
  assign n61902 = ~n61893 & n61900;
  assign n61903 = ~n61901 & ~n61902;
  assign n61904 = n61066 & ~n61903;
  assign n61905 = n59265 & ~n61881;
  assign n61906 = n59108 & ~n61881;
  assign n61907 = ~n61905 & ~n61906;
  assign n61908 = P2_P3_INSTADDRPOINTER_REG_6_ & ~n61815;
  assign n61909 = ~P2_P3_INSTADDRPOINTER_REG_6_ & n61815;
  assign n61910 = ~n61811 & ~n61909;
  assign n61911 = ~n61908 & ~n61910;
  assign n61912 = ~n61793 & n61812;
  assign n61913 = n61065 & n61912;
  assign n61914 = ~n61065 & ~n61912;
  assign n61915 = ~n61913 & ~n61914;
  assign n61916 = ~P2_P3_INSTADDRPOINTER_REG_7_ & ~n61915;
  assign n61917 = P2_P3_INSTADDRPOINTER_REG_7_ & n61915;
  assign n61918 = ~n61916 & ~n61917;
  assign n61919 = n61911 & ~n61918;
  assign n61920 = ~n61911 & n61918;
  assign n61921 = ~n61919 & ~n61920;
  assign n61922 = n61068 & ~n61921;
  assign n61923 = n61907 & ~n61922;
  assign n61924 = n61085 & ~n61881;
  assign n61925 = n61078 & ~n61881;
  assign n61926 = n61074 & ~n61881;
  assign n61927 = n59112 & ~n61881;
  assign n61928 = ~n61924 & ~n61925;
  assign n61929 = ~n61926 & n61928;
  assign n61930 = ~n61927 & n61929;
  assign n61931 = n58968 & ~n61875;
  assign n61932 = n59046 & ~n61875;
  assign n61933 = n59050 & ~n61875;
  assign n61934 = P2_P3_INSTADDRPOINTER_REG_6_ & n61834;
  assign n61935 = ~P2_P3_INSTADDRPOINTER_REG_7_ & n61934;
  assign n61936 = P2_P3_INSTADDRPOINTER_REG_7_ & ~n61934;
  assign n61937 = ~n61935 & ~n61936;
  assign n61938 = n59066 & ~n61937;
  assign n61939 = n59058 & ~n61937;
  assign n61940 = ~n61931 & ~n61932;
  assign n61941 = ~n61933 & n61940;
  assign n61942 = ~n61938 & n61941;
  assign n61943 = ~n61939 & n61942;
  assign n61944 = P2_P3_INSTADDRPOINTER_REG_6_ & ~n61853;
  assign n61945 = ~P2_P3_INSTADDRPOINTER_REG_6_ & n61853;
  assign n61946 = ~n61849 & ~n61945;
  assign n61947 = ~n61944 & ~n61946;
  assign n61948 = ~n61793 & n61850;
  assign n61949 = n61065 & n61948;
  assign n61950 = ~n61065 & ~n61948;
  assign n61951 = ~n61949 & ~n61950;
  assign n61952 = ~P2_P3_INSTADDRPOINTER_REG_7_ & ~n61951;
  assign n61953 = P2_P3_INSTADDRPOINTER_REG_7_ & n61951;
  assign n61954 = ~n61952 & ~n61953;
  assign n61955 = n61947 & ~n61954;
  assign n61956 = ~n61947 & n61954;
  assign n61957 = ~n61955 & ~n61956;
  assign n61958 = n59069 & ~n61957;
  assign n61959 = n61930 & n61943;
  assign n61960 = ~n61958 & n61959;
  assign n61961 = n61888 & ~n61889;
  assign n61962 = ~n61904 & n61961;
  assign n61963 = n61923 & n61962;
  assign n61964 = n61960 & n61963;
  assign n61965 = n60961 & ~n61964;
  assign n61966 = ~n61870 & ~n61871;
  assign n11076 = n61965 | ~n61966;
  assign n61968 = P2_P3_INSTADDRPOINTER_REG_8_ & n60960;
  assign n61969 = P2_P3_REIP_REG_8_ & n61105;
  assign n61970 = P2_P3_INSTADDRPOINTER_REG_7_ & n61872;
  assign n61971 = ~P2_P3_INSTADDRPOINTER_REG_8_ & n61970;
  assign n61972 = P2_P3_INSTADDRPOINTER_REG_8_ & ~n61970;
  assign n61973 = ~n61971 & ~n61972;
  assign n61974 = n59226 & ~n61973;
  assign n61975 = n59227 & ~n61973;
  assign n61976 = n59042 & ~n61973;
  assign n61977 = P2_P3_INSTADDRPOINTER_REG_7_ & n61878;
  assign n61978 = ~P2_P3_INSTADDRPOINTER_REG_8_ & n61977;
  assign n61979 = P2_P3_INSTADDRPOINTER_REG_8_ & ~n61977;
  assign n61980 = ~n61978 & ~n61979;
  assign n61981 = n60972 & ~n61980;
  assign n61982 = n60969 & ~n61980;
  assign n61983 = ~n61976 & ~n61981;
  assign n61984 = ~n61982 & n61983;
  assign n61985 = ~n61974 & ~n61975;
  assign n61986 = n61984 & n61985;
  assign n61987 = ~n59155 & ~n61980;
  assign n61988 = ~P2_P3_INSTADDRPOINTER_REG_7_ & ~n61897;
  assign n61989 = ~n61893 & ~n61988;
  assign n61990 = P2_P3_INSTADDRPOINTER_REG_7_ & n61897;
  assign n61991 = ~n61989 & ~n61990;
  assign n61992 = ~P2_P3_INSTADDRPOINTER_REG_8_ & ~n61896;
  assign n61993 = P2_P3_INSTADDRPOINTER_REG_8_ & n61896;
  assign n61994 = ~n61992 & ~n61993;
  assign n61995 = n61991 & ~n61994;
  assign n61996 = ~n61991 & n61994;
  assign n61997 = ~n61995 & ~n61996;
  assign n61998 = n61066 & ~n61997;
  assign n61999 = n59265 & ~n61980;
  assign n62000 = n59108 & ~n61980;
  assign n62001 = ~n61999 & ~n62000;
  assign n62002 = ~n61911 & ~n61915;
  assign n62003 = P2_P3_INSTADDRPOINTER_REG_7_ & ~n61911;
  assign n62004 = P2_P3_INSTADDRPOINTER_REG_7_ & ~n61915;
  assign n62005 = ~n62002 & ~n62003;
  assign n62006 = ~n62004 & n62005;
  assign n62007 = n61812 & n61895;
  assign n62008 = ~P2_P3_INSTADDRPOINTER_REG_8_ & n62007;
  assign n62009 = P2_P3_INSTADDRPOINTER_REG_8_ & ~n62007;
  assign n62010 = ~n62008 & ~n62009;
  assign n62011 = n62006 & ~n62010;
  assign n62012 = ~n62006 & n62010;
  assign n62013 = ~n62011 & ~n62012;
  assign n62014 = n61068 & ~n62013;
  assign n62015 = n62001 & ~n62014;
  assign n62016 = n61085 & ~n61980;
  assign n62017 = n59112 & ~n61980;
  assign n62018 = n61074 & ~n61980;
  assign n62019 = n61078 & ~n61980;
  assign n62020 = ~n62016 & ~n62017;
  assign n62021 = ~n62018 & n62020;
  assign n62022 = ~n62019 & n62021;
  assign n62023 = n58968 & ~n61973;
  assign n62024 = n59046 & ~n61973;
  assign n62025 = n59050 & ~n61973;
  assign n62026 = P2_P3_INSTADDRPOINTER_REG_7_ & n61934;
  assign n62027 = ~P2_P3_INSTADDRPOINTER_REG_8_ & n62026;
  assign n62028 = P2_P3_INSTADDRPOINTER_REG_8_ & ~n62026;
  assign n62029 = ~n62027 & ~n62028;
  assign n62030 = n59066 & ~n62029;
  assign n62031 = n59058 & ~n62029;
  assign n62032 = ~n62023 & ~n62024;
  assign n62033 = ~n62025 & n62032;
  assign n62034 = ~n62030 & n62033;
  assign n62035 = ~n62031 & n62034;
  assign n62036 = ~n61947 & ~n61951;
  assign n62037 = P2_P3_INSTADDRPOINTER_REG_7_ & ~n61947;
  assign n62038 = P2_P3_INSTADDRPOINTER_REG_7_ & ~n61951;
  assign n62039 = ~n62036 & ~n62037;
  assign n62040 = ~n62038 & n62039;
  assign n62041 = n61850 & n61895;
  assign n62042 = ~P2_P3_INSTADDRPOINTER_REG_8_ & n62041;
  assign n62043 = P2_P3_INSTADDRPOINTER_REG_8_ & ~n62041;
  assign n62044 = ~n62042 & ~n62043;
  assign n62045 = n62040 & ~n62044;
  assign n62046 = ~n62040 & n62044;
  assign n62047 = ~n62045 & ~n62046;
  assign n62048 = n59069 & ~n62047;
  assign n62049 = n62022 & n62035;
  assign n62050 = ~n62048 & n62049;
  assign n62051 = n61986 & ~n61987;
  assign n62052 = ~n61998 & n62051;
  assign n62053 = n62015 & n62052;
  assign n62054 = n62050 & n62053;
  assign n62055 = n60961 & ~n62054;
  assign n62056 = ~n61968 & ~n61969;
  assign n11081 = n62055 | ~n62056;
  assign n62058 = P2_P3_INSTADDRPOINTER_REG_9_ & n60960;
  assign n62059 = P2_P3_REIP_REG_9_ & n61105;
  assign n62060 = P2_P3_INSTADDRPOINTER_REG_8_ & n61970;
  assign n62061 = ~P2_P3_INSTADDRPOINTER_REG_9_ & n62060;
  assign n62062 = P2_P3_INSTADDRPOINTER_REG_9_ & ~n62060;
  assign n62063 = ~n62061 & ~n62062;
  assign n62064 = n59226 & ~n62063;
  assign n62065 = n59227 & ~n62063;
  assign n62066 = P2_P3_INSTADDRPOINTER_REG_8_ & n61977;
  assign n62067 = ~P2_P3_INSTADDRPOINTER_REG_9_ & n62066;
  assign n62068 = P2_P3_INSTADDRPOINTER_REG_9_ & ~n62066;
  assign n62069 = ~n62067 & ~n62068;
  assign n62070 = n60969 & ~n62069;
  assign n62071 = n59042 & ~n62063;
  assign n62072 = n60972 & ~n62069;
  assign n62073 = ~n62071 & ~n62072;
  assign n62074 = ~n62064 & ~n62065;
  assign n62075 = ~n62070 & n62074;
  assign n62076 = n62073 & n62075;
  assign n62077 = ~n59155 & ~n62069;
  assign n62078 = ~P2_P3_INSTADDRPOINTER_REG_8_ & n61896;
  assign n62079 = ~n61991 & ~n62078;
  assign n62080 = P2_P3_INSTADDRPOINTER_REG_8_ & ~n61896;
  assign n62081 = ~n62079 & ~n62080;
  assign n62082 = P2_P3_INSTADDRPOINTER_REG_9_ & n61896;
  assign n62083 = ~P2_P3_INSTADDRPOINTER_REG_9_ & ~n61896;
  assign n62084 = ~n62082 & ~n62083;
  assign n62085 = n62081 & ~n62084;
  assign n62086 = P2_P3_INSTADDRPOINTER_REG_9_ & ~n61896;
  assign n62087 = ~P2_P3_INSTADDRPOINTER_REG_9_ & n61896;
  assign n62088 = ~n62086 & ~n62087;
  assign n62089 = ~n62081 & ~n62088;
  assign n62090 = ~n62085 & ~n62089;
  assign n62091 = n61066 & ~n62090;
  assign n62092 = n59265 & ~n62069;
  assign n62093 = n59108 & ~n62069;
  assign n62094 = ~n62092 & ~n62093;
  assign n62095 = P2_P3_INSTADDRPOINTER_REG_8_ & n62007;
  assign n62096 = ~P2_P3_INSTADDRPOINTER_REG_8_ & ~n62007;
  assign n62097 = ~n62006 & ~n62096;
  assign n62098 = ~n62095 & ~n62097;
  assign n62099 = ~P2_P3_INSTADDRPOINTER_REG_9_ & n62098;
  assign n62100 = P2_P3_INSTADDRPOINTER_REG_9_ & ~n62098;
  assign n62101 = ~n62099 & ~n62100;
  assign n62102 = n61068 & n62101;
  assign n62103 = n62094 & ~n62102;
  assign n62104 = n61085 & ~n62069;
  assign n62105 = n59112 & ~n62069;
  assign n62106 = n61074 & ~n62069;
  assign n62107 = n61078 & ~n62069;
  assign n62108 = ~n62104 & ~n62105;
  assign n62109 = ~n62106 & n62108;
  assign n62110 = ~n62107 & n62109;
  assign n62111 = n58968 & ~n62063;
  assign n62112 = n59046 & ~n62063;
  assign n62113 = n59050 & ~n62063;
  assign n62114 = P2_P3_INSTADDRPOINTER_REG_8_ & n62026;
  assign n62115 = ~P2_P3_INSTADDRPOINTER_REG_9_ & n62114;
  assign n62116 = P2_P3_INSTADDRPOINTER_REG_9_ & ~n62114;
  assign n62117 = ~n62115 & ~n62116;
  assign n62118 = n59066 & ~n62117;
  assign n62119 = n59058 & ~n62117;
  assign n62120 = ~n62111 & ~n62112;
  assign n62121 = ~n62113 & n62120;
  assign n62122 = ~n62118 & n62121;
  assign n62123 = ~n62119 & n62122;
  assign n62124 = P2_P3_INSTADDRPOINTER_REG_8_ & n62041;
  assign n62125 = ~P2_P3_INSTADDRPOINTER_REG_8_ & ~n62041;
  assign n62126 = ~n62040 & ~n62125;
  assign n62127 = ~n62124 & ~n62126;
  assign n62128 = ~P2_P3_INSTADDRPOINTER_REG_9_ & n62127;
  assign n62129 = P2_P3_INSTADDRPOINTER_REG_9_ & ~n62127;
  assign n62130 = ~n62128 & ~n62129;
  assign n62131 = n59069 & n62130;
  assign n62132 = n62110 & n62123;
  assign n62133 = ~n62131 & n62132;
  assign n62134 = n62076 & ~n62077;
  assign n62135 = ~n62091 & n62134;
  assign n62136 = n62103 & n62135;
  assign n62137 = n62133 & n62136;
  assign n62138 = n60961 & ~n62137;
  assign n62139 = ~n62058 & ~n62059;
  assign n11086 = n62138 | ~n62139;
  assign n62141 = P2_P3_INSTADDRPOINTER_REG_10_ & n60960;
  assign n62142 = P2_P3_REIP_REG_10_ & n61105;
  assign n62143 = P2_P3_INSTADDRPOINTER_REG_9_ & n62060;
  assign n62144 = ~P2_P3_INSTADDRPOINTER_REG_10_ & n62143;
  assign n62145 = P2_P3_INSTADDRPOINTER_REG_10_ & ~n62143;
  assign n62146 = ~n62144 & ~n62145;
  assign n62147 = n59226 & ~n62146;
  assign n62148 = n59227 & ~n62146;
  assign n62149 = P2_P3_INSTADDRPOINTER_REG_9_ & n62066;
  assign n62150 = ~P2_P3_INSTADDRPOINTER_REG_10_ & n62149;
  assign n62151 = P2_P3_INSTADDRPOINTER_REG_10_ & ~n62149;
  assign n62152 = ~n62150 & ~n62151;
  assign n62153 = n60969 & ~n62152;
  assign n62154 = n59042 & ~n62146;
  assign n62155 = n60972 & ~n62152;
  assign n62156 = ~n62154 & ~n62155;
  assign n62157 = ~n62147 & ~n62148;
  assign n62158 = ~n62153 & n62157;
  assign n62159 = n62156 & n62158;
  assign n62160 = ~n59155 & ~n62152;
  assign n62161 = ~n62078 & ~n62087;
  assign n62162 = ~n61991 & n62161;
  assign n62163 = ~n62080 & ~n62086;
  assign n62164 = ~n62162 & n62163;
  assign n62165 = ~P2_P3_INSTADDRPOINTER_REG_10_ & ~n61896;
  assign n62166 = P2_P3_INSTADDRPOINTER_REG_10_ & n61896;
  assign n62167 = ~n62165 & ~n62166;
  assign n62168 = n62164 & ~n62167;
  assign n62169 = P2_P3_INSTADDRPOINTER_REG_10_ & ~n61896;
  assign n62170 = ~P2_P3_INSTADDRPOINTER_REG_10_ & n61896;
  assign n62171 = ~n62169 & ~n62170;
  assign n62172 = ~n62164 & ~n62171;
  assign n62173 = ~n62168 & ~n62172;
  assign n62174 = n61066 & ~n62173;
  assign n62175 = n59265 & ~n62152;
  assign n62176 = n59108 & ~n62152;
  assign n62177 = ~n62175 & ~n62176;
  assign n62178 = ~P2_P3_INSTADDRPOINTER_REG_10_ & ~n62100;
  assign n62179 = P2_P3_INSTADDRPOINTER_REG_9_ & P2_P3_INSTADDRPOINTER_REG_10_;
  assign n62180 = ~n62098 & n62179;
  assign n62181 = ~n62178 & ~n62180;
  assign n62182 = n61068 & n62181;
  assign n62183 = n62177 & ~n62182;
  assign n62184 = n61085 & ~n62152;
  assign n62185 = n59112 & ~n62152;
  assign n62186 = n61074 & ~n62152;
  assign n62187 = n61078 & ~n62152;
  assign n62188 = ~n62184 & ~n62185;
  assign n62189 = ~n62186 & n62188;
  assign n62190 = ~n62187 & n62189;
  assign n62191 = n58968 & ~n62146;
  assign n62192 = n59046 & ~n62146;
  assign n62193 = n59050 & ~n62146;
  assign n62194 = P2_P3_INSTADDRPOINTER_REG_9_ & n62114;
  assign n62195 = ~P2_P3_INSTADDRPOINTER_REG_10_ & n62194;
  assign n62196 = P2_P3_INSTADDRPOINTER_REG_10_ & ~n62194;
  assign n62197 = ~n62195 & ~n62196;
  assign n62198 = n59066 & ~n62197;
  assign n62199 = n59058 & ~n62197;
  assign n62200 = ~n62191 & ~n62192;
  assign n62201 = ~n62193 & n62200;
  assign n62202 = ~n62198 & n62201;
  assign n62203 = ~n62199 & n62202;
  assign n62204 = ~P2_P3_INSTADDRPOINTER_REG_10_ & ~n62129;
  assign n62205 = ~n62127 & n62179;
  assign n62206 = ~n62204 & ~n62205;
  assign n62207 = n59069 & n62206;
  assign n62208 = n62190 & n62203;
  assign n62209 = ~n62207 & n62208;
  assign n62210 = n62159 & ~n62160;
  assign n62211 = ~n62174 & n62210;
  assign n62212 = n62183 & n62211;
  assign n62213 = n62209 & n62212;
  assign n62214 = n60961 & ~n62213;
  assign n62215 = ~n62141 & ~n62142;
  assign n11091 = n62214 | ~n62215;
  assign n62217 = P2_P3_INSTADDRPOINTER_REG_11_ & n60960;
  assign n62218 = P2_P3_REIP_REG_11_ & n61105;
  assign n62219 = ~n62217 & ~n62218;
  assign n62220 = P2_P3_INSTADDRPOINTER_REG_10_ & n62149;
  assign n62221 = ~P2_P3_INSTADDRPOINTER_REG_11_ & n62220;
  assign n62222 = P2_P3_INSTADDRPOINTER_REG_11_ & ~n62220;
  assign n62223 = ~n62221 & ~n62222;
  assign n62224 = n61085 & ~n62223;
  assign n62225 = n59112 & ~n62223;
  assign n62226 = n61074 & ~n62223;
  assign n62227 = n61078 & ~n62223;
  assign n62228 = ~n62224 & ~n62225;
  assign n62229 = ~n62226 & n62228;
  assign n62230 = ~n62227 & n62229;
  assign n62231 = P2_P3_INSTADDRPOINTER_REG_10_ & n62143;
  assign n62232 = ~P2_P3_INSTADDRPOINTER_REG_11_ & n62231;
  assign n62233 = P2_P3_INSTADDRPOINTER_REG_11_ & ~n62231;
  assign n62234 = ~n62232 & ~n62233;
  assign n62235 = n58968 & ~n62234;
  assign n62236 = n59046 & ~n62234;
  assign n62237 = n59050 & ~n62234;
  assign n62238 = P2_P3_INSTADDRPOINTER_REG_10_ & n62194;
  assign n62239 = ~P2_P3_INSTADDRPOINTER_REG_11_ & n62238;
  assign n62240 = P2_P3_INSTADDRPOINTER_REG_11_ & ~n62238;
  assign n62241 = ~n62239 & ~n62240;
  assign n62242 = n59066 & ~n62241;
  assign n62243 = n59058 & ~n62241;
  assign n62244 = ~n62235 & ~n62236;
  assign n62245 = ~n62237 & n62244;
  assign n62246 = ~n62242 & n62245;
  assign n62247 = ~n62243 & n62246;
  assign n62248 = P2_P3_INSTADDRPOINTER_REG_11_ & ~n62205;
  assign n62249 = ~P2_P3_INSTADDRPOINTER_REG_11_ & n62205;
  assign n62250 = ~n62248 & ~n62249;
  assign n62251 = n59069 & ~n62250;
  assign n62252 = n62230 & n62247;
  assign n62253 = ~n62251 & n62252;
  assign n62254 = n59265 & ~n62223;
  assign n62255 = n59108 & ~n62223;
  assign n62256 = ~n62254 & ~n62255;
  assign n62257 = ~n59155 & ~n62223;
  assign n62258 = n62163 & ~n62169;
  assign n62259 = n62161 & ~n62170;
  assign n62260 = ~n61991 & n62259;
  assign n62261 = n62258 & ~n62260;
  assign n62262 = ~P2_P3_INSTADDRPOINTER_REG_11_ & ~n61896;
  assign n62263 = P2_P3_INSTADDRPOINTER_REG_11_ & n61896;
  assign n62264 = ~n62262 & ~n62263;
  assign n62265 = n62261 & ~n62264;
  assign n62266 = ~n62261 & n62264;
  assign n62267 = ~n62265 & ~n62266;
  assign n62268 = n61066 & ~n62267;
  assign n62269 = n59226 & ~n62234;
  assign n62270 = n59227 & ~n62234;
  assign n62271 = n60969 & ~n62223;
  assign n62272 = n59042 & ~n62234;
  assign n62273 = n60972 & ~n62223;
  assign n62274 = ~n62272 & ~n62273;
  assign n62275 = ~n62269 & ~n62270;
  assign n62276 = ~n62271 & n62275;
  assign n62277 = n62274 & n62276;
  assign n62278 = P2_P3_INSTADDRPOINTER_REG_11_ & ~n62180;
  assign n62279 = ~P2_P3_INSTADDRPOINTER_REG_11_ & n62180;
  assign n62280 = ~n62278 & ~n62279;
  assign n62281 = n61068 & ~n62280;
  assign n62282 = n62256 & ~n62257;
  assign n62283 = ~n62268 & n62282;
  assign n62284 = n62277 & n62283;
  assign n62285 = ~n62281 & n62284;
  assign n62286 = n62253 & n62285;
  assign n62287 = n60961 & ~n62286;
  assign n11096 = ~n62219 | n62287;
  assign n62289 = P2_P3_INSTADDRPOINTER_REG_12_ & n60960;
  assign n62290 = P2_P3_REIP_REG_12_ & n61105;
  assign n62291 = P2_P3_INSTADDRPOINTER_REG_11_ & n62231;
  assign n62292 = ~P2_P3_INSTADDRPOINTER_REG_12_ & n62291;
  assign n62293 = P2_P3_INSTADDRPOINTER_REG_12_ & ~n62291;
  assign n62294 = ~n62292 & ~n62293;
  assign n62295 = n59226 & ~n62294;
  assign n62296 = n59227 & ~n62294;
  assign n62297 = P2_P3_INSTADDRPOINTER_REG_11_ & n62220;
  assign n62298 = ~P2_P3_INSTADDRPOINTER_REG_12_ & n62297;
  assign n62299 = P2_P3_INSTADDRPOINTER_REG_12_ & ~n62297;
  assign n62300 = ~n62298 & ~n62299;
  assign n62301 = n60969 & ~n62300;
  assign n62302 = n59042 & ~n62294;
  assign n62303 = n60972 & ~n62300;
  assign n62304 = ~n62302 & ~n62303;
  assign n62305 = ~n62295 & ~n62296;
  assign n62306 = ~n62301 & n62305;
  assign n62307 = n62304 & n62306;
  assign n62308 = ~n59155 & ~n62300;
  assign n62309 = ~P2_P3_INSTADDRPOINTER_REG_12_ & ~n61896;
  assign n62310 = P2_P3_INSTADDRPOINTER_REG_12_ & n61896;
  assign n62311 = ~n62309 & ~n62310;
  assign n62312 = P2_P3_INSTADDRPOINTER_REG_11_ & ~n61896;
  assign n62313 = ~P2_P3_INSTADDRPOINTER_REG_11_ & n61896;
  assign n62314 = ~n62261 & ~n62313;
  assign n62315 = ~n62312 & ~n62314;
  assign n62316 = ~n62311 & n62315;
  assign n62317 = ~P2_P3_INSTADDRPOINTER_REG_12_ & n61896;
  assign n62318 = P2_P3_INSTADDRPOINTER_REG_12_ & ~n61896;
  assign n62319 = ~n62317 & ~n62318;
  assign n62320 = ~n62315 & ~n62319;
  assign n62321 = ~n62316 & ~n62320;
  assign n62322 = n61066 & ~n62321;
  assign n62323 = n59265 & ~n62300;
  assign n62324 = n59108 & ~n62300;
  assign n62325 = ~n62323 & ~n62324;
  assign n62326 = P2_P3_INSTADDRPOINTER_REG_11_ & n62180;
  assign n62327 = ~P2_P3_INSTADDRPOINTER_REG_12_ & ~n62326;
  assign n62328 = P2_P3_INSTADDRPOINTER_REG_11_ & P2_P3_INSTADDRPOINTER_REG_12_;
  assign n62329 = n62180 & n62328;
  assign n62330 = ~n62327 & ~n62329;
  assign n62331 = n61068 & n62330;
  assign n62332 = n62325 & ~n62331;
  assign n62333 = n61085 & ~n62300;
  assign n62334 = n59112 & ~n62300;
  assign n62335 = n61074 & ~n62300;
  assign n62336 = n61078 & ~n62300;
  assign n62337 = ~n62333 & ~n62334;
  assign n62338 = ~n62335 & n62337;
  assign n62339 = ~n62336 & n62338;
  assign n62340 = n58968 & ~n62294;
  assign n62341 = n59046 & ~n62294;
  assign n62342 = n59050 & ~n62294;
  assign n62343 = P2_P3_INSTADDRPOINTER_REG_11_ & n62238;
  assign n62344 = ~P2_P3_INSTADDRPOINTER_REG_12_ & n62343;
  assign n62345 = P2_P3_INSTADDRPOINTER_REG_12_ & ~n62343;
  assign n62346 = ~n62344 & ~n62345;
  assign n62347 = n59066 & ~n62346;
  assign n62348 = n59058 & ~n62346;
  assign n62349 = ~n62340 & ~n62341;
  assign n62350 = ~n62342 & n62349;
  assign n62351 = ~n62347 & n62350;
  assign n62352 = ~n62348 & n62351;
  assign n62353 = P2_P3_INSTADDRPOINTER_REG_11_ & n62205;
  assign n62354 = ~P2_P3_INSTADDRPOINTER_REG_12_ & ~n62353;
  assign n62355 = n62205 & n62328;
  assign n62356 = ~n62354 & ~n62355;
  assign n62357 = n59069 & n62356;
  assign n62358 = n62339 & n62352;
  assign n62359 = ~n62357 & n62358;
  assign n62360 = n62307 & ~n62308;
  assign n62361 = ~n62322 & n62360;
  assign n62362 = n62332 & n62361;
  assign n62363 = n62359 & n62362;
  assign n62364 = n60961 & ~n62363;
  assign n62365 = ~n62289 & ~n62290;
  assign n11101 = n62364 | ~n62365;
  assign n62367 = P2_P3_INSTADDRPOINTER_REG_13_ & n60960;
  assign n62368 = P2_P3_REIP_REG_13_ & n61105;
  assign n62369 = P2_P3_INSTADDRPOINTER_REG_12_ & n62291;
  assign n62370 = ~P2_P3_INSTADDRPOINTER_REG_13_ & n62369;
  assign n62371 = P2_P3_INSTADDRPOINTER_REG_13_ & ~n62369;
  assign n62372 = ~n62370 & ~n62371;
  assign n62373 = n59226 & ~n62372;
  assign n62374 = n59227 & ~n62372;
  assign n62375 = P2_P3_INSTADDRPOINTER_REG_12_ & n62297;
  assign n62376 = ~P2_P3_INSTADDRPOINTER_REG_13_ & n62375;
  assign n62377 = P2_P3_INSTADDRPOINTER_REG_13_ & ~n62375;
  assign n62378 = ~n62376 & ~n62377;
  assign n62379 = n60969 & ~n62378;
  assign n62380 = n59042 & ~n62372;
  assign n62381 = n60972 & ~n62378;
  assign n62382 = ~n62380 & ~n62381;
  assign n62383 = ~n62373 & ~n62374;
  assign n62384 = ~n62379 & n62383;
  assign n62385 = n62382 & n62384;
  assign n62386 = ~n59155 & ~n62378;
  assign n62387 = P2_P3_INSTADDRPOINTER_REG_13_ & ~n61896;
  assign n62388 = P2_P3_INSTADDRPOINTER_REG_12_ & P2_P3_INSTADDRPOINTER_REG_13_;
  assign n62389 = n61896 & ~n62388;
  assign n62390 = ~n62387 & ~n62389;
  assign n62391 = n62315 & ~n62318;
  assign n62392 = n62390 & ~n62391;
  assign n62393 = ~P2_P3_INSTADDRPOINTER_REG_13_ & ~n61896;
  assign n62394 = P2_P3_INSTADDRPOINTER_REG_13_ & n61896;
  assign n62395 = ~n62393 & ~n62394;
  assign n62396 = ~n62318 & n62395;
  assign n62397 = ~n62315 & ~n62317;
  assign n62398 = n62396 & ~n62397;
  assign n62399 = ~n62392 & ~n62398;
  assign n62400 = n61066 & n62399;
  assign n62401 = n59265 & ~n62378;
  assign n62402 = n59108 & ~n62378;
  assign n62403 = ~n62401 & ~n62402;
  assign n62404 = ~P2_P3_INSTADDRPOINTER_REG_13_ & ~n62329;
  assign n62405 = P2_P3_INSTADDRPOINTER_REG_13_ & n62329;
  assign n62406 = ~n62404 & ~n62405;
  assign n62407 = n61068 & n62406;
  assign n62408 = n62403 & ~n62407;
  assign n62409 = n61085 & ~n62378;
  assign n62410 = n59112 & ~n62378;
  assign n62411 = n61074 & ~n62378;
  assign n62412 = n61078 & ~n62378;
  assign n62413 = ~n62409 & ~n62410;
  assign n62414 = ~n62411 & n62413;
  assign n62415 = ~n62412 & n62414;
  assign n62416 = n58968 & ~n62372;
  assign n62417 = n59046 & ~n62372;
  assign n62418 = n59050 & ~n62372;
  assign n62419 = P2_P3_INSTADDRPOINTER_REG_12_ & n62343;
  assign n62420 = ~P2_P3_INSTADDRPOINTER_REG_13_ & n62419;
  assign n62421 = P2_P3_INSTADDRPOINTER_REG_13_ & ~n62419;
  assign n62422 = ~n62420 & ~n62421;
  assign n62423 = n59066 & ~n62422;
  assign n62424 = n59058 & ~n62422;
  assign n62425 = ~n62416 & ~n62417;
  assign n62426 = ~n62418 & n62425;
  assign n62427 = ~n62423 & n62426;
  assign n62428 = ~n62424 & n62427;
  assign n62429 = ~P2_P3_INSTADDRPOINTER_REG_13_ & ~n62355;
  assign n62430 = P2_P3_INSTADDRPOINTER_REG_13_ & n62355;
  assign n62431 = ~n62429 & ~n62430;
  assign n62432 = n59069 & n62431;
  assign n62433 = n62415 & n62428;
  assign n62434 = ~n62432 & n62433;
  assign n62435 = n62385 & ~n62386;
  assign n62436 = ~n62400 & n62435;
  assign n62437 = n62408 & n62436;
  assign n62438 = n62434 & n62437;
  assign n62439 = n60961 & ~n62438;
  assign n62440 = ~n62367 & ~n62368;
  assign n11106 = n62439 | ~n62440;
  assign n62442 = P2_P3_INSTADDRPOINTER_REG_14_ & n60960;
  assign n62443 = P2_P3_REIP_REG_14_ & n61105;
  assign n62444 = ~n62442 & ~n62443;
  assign n62445 = P2_P3_INSTADDRPOINTER_REG_13_ & n62375;
  assign n62446 = ~P2_P3_INSTADDRPOINTER_REG_14_ & n62445;
  assign n62447 = P2_P3_INSTADDRPOINTER_REG_14_ & ~n62445;
  assign n62448 = ~n62446 & ~n62447;
  assign n62449 = n61085 & ~n62448;
  assign n62450 = n59112 & ~n62448;
  assign n62451 = n61074 & ~n62448;
  assign n62452 = n61078 & ~n62448;
  assign n62453 = ~n62449 & ~n62450;
  assign n62454 = ~n62451 & n62453;
  assign n62455 = ~n62452 & n62454;
  assign n62456 = P2_P3_INSTADDRPOINTER_REG_13_ & n62369;
  assign n62457 = ~P2_P3_INSTADDRPOINTER_REG_14_ & n62456;
  assign n62458 = P2_P3_INSTADDRPOINTER_REG_14_ & ~n62456;
  assign n62459 = ~n62457 & ~n62458;
  assign n62460 = n58968 & ~n62459;
  assign n62461 = n59046 & ~n62459;
  assign n62462 = n59050 & ~n62459;
  assign n62463 = P2_P3_INSTADDRPOINTER_REG_13_ & n62419;
  assign n62464 = ~P2_P3_INSTADDRPOINTER_REG_14_ & n62463;
  assign n62465 = P2_P3_INSTADDRPOINTER_REG_14_ & ~n62463;
  assign n62466 = ~n62464 & ~n62465;
  assign n62467 = n59066 & ~n62466;
  assign n62468 = n59058 & ~n62466;
  assign n62469 = ~n62460 & ~n62461;
  assign n62470 = ~n62462 & n62469;
  assign n62471 = ~n62467 & n62470;
  assign n62472 = ~n62468 & n62471;
  assign n62473 = ~P2_P3_INSTADDRPOINTER_REG_14_ & n62430;
  assign n62474 = P2_P3_INSTADDRPOINTER_REG_14_ & ~n62430;
  assign n62475 = ~n62473 & ~n62474;
  assign n62476 = n59069 & ~n62475;
  assign n62477 = n62455 & n62472;
  assign n62478 = ~n62476 & n62477;
  assign n62479 = n59265 & ~n62448;
  assign n62480 = n59108 & ~n62448;
  assign n62481 = ~n62479 & ~n62480;
  assign n62482 = ~n59155 & ~n62448;
  assign n62483 = n59226 & ~n62459;
  assign n62484 = n59227 & ~n62459;
  assign n62485 = n60969 & ~n62448;
  assign n62486 = n59042 & ~n62459;
  assign n62487 = n60972 & ~n62448;
  assign n62488 = ~n62486 & ~n62487;
  assign n62489 = ~n62483 & ~n62484;
  assign n62490 = ~n62485 & n62489;
  assign n62491 = n62488 & n62490;
  assign n62492 = ~n62318 & ~n62387;
  assign n62493 = ~n62312 & n62492;
  assign n62494 = ~n62313 & ~n62389;
  assign n62495 = ~n62261 & n62494;
  assign n62496 = n62493 & ~n62495;
  assign n62497 = ~P2_P3_INSTADDRPOINTER_REG_14_ & ~n61896;
  assign n62498 = P2_P3_INSTADDRPOINTER_REG_14_ & n61896;
  assign n62499 = ~n62497 & ~n62498;
  assign n62500 = n62496 & ~n62499;
  assign n62501 = ~n62496 & n62499;
  assign n62502 = ~n62500 & ~n62501;
  assign n62503 = n61066 & ~n62502;
  assign n62504 = ~P2_P3_INSTADDRPOINTER_REG_14_ & n62405;
  assign n62505 = P2_P3_INSTADDRPOINTER_REG_14_ & ~n62405;
  assign n62506 = ~n62504 & ~n62505;
  assign n62507 = n61068 & ~n62506;
  assign n62508 = n62481 & ~n62482;
  assign n62509 = n62491 & n62508;
  assign n62510 = ~n62503 & n62509;
  assign n62511 = ~n62507 & n62510;
  assign n62512 = n62478 & n62511;
  assign n62513 = n60961 & ~n62512;
  assign n11111 = ~n62444 | n62513;
  assign n62515 = P2_P3_INSTADDRPOINTER_REG_15_ & n60960;
  assign n62516 = P2_P3_REIP_REG_15_ & n61105;
  assign n62517 = ~n62515 & ~n62516;
  assign n62518 = P2_P3_INSTADDRPOINTER_REG_14_ & n62445;
  assign n62519 = ~P2_P3_INSTADDRPOINTER_REG_15_ & n62518;
  assign n62520 = P2_P3_INSTADDRPOINTER_REG_15_ & ~n62518;
  assign n62521 = ~n62519 & ~n62520;
  assign n62522 = n61085 & ~n62521;
  assign n62523 = n59112 & ~n62521;
  assign n62524 = n61074 & ~n62521;
  assign n62525 = n61078 & ~n62521;
  assign n62526 = ~n62522 & ~n62523;
  assign n62527 = ~n62524 & n62526;
  assign n62528 = ~n62525 & n62527;
  assign n62529 = P2_P3_INSTADDRPOINTER_REG_14_ & n62456;
  assign n62530 = ~P2_P3_INSTADDRPOINTER_REG_15_ & n62529;
  assign n62531 = P2_P3_INSTADDRPOINTER_REG_15_ & ~n62529;
  assign n62532 = ~n62530 & ~n62531;
  assign n62533 = n58968 & ~n62532;
  assign n62534 = n59046 & ~n62532;
  assign n62535 = n59050 & ~n62532;
  assign n62536 = P2_P3_INSTADDRPOINTER_REG_14_ & n62463;
  assign n62537 = ~P2_P3_INSTADDRPOINTER_REG_15_ & n62536;
  assign n62538 = P2_P3_INSTADDRPOINTER_REG_15_ & ~n62536;
  assign n62539 = ~n62537 & ~n62538;
  assign n62540 = n59066 & ~n62539;
  assign n62541 = n59058 & ~n62539;
  assign n62542 = ~n62533 & ~n62534;
  assign n62543 = ~n62535 & n62542;
  assign n62544 = ~n62540 & n62543;
  assign n62545 = ~n62541 & n62544;
  assign n62546 = P2_P3_INSTADDRPOINTER_REG_14_ & n62430;
  assign n62547 = ~P2_P3_INSTADDRPOINTER_REG_15_ & ~n62546;
  assign n62548 = P2_P3_INSTADDRPOINTER_REG_14_ & P2_P3_INSTADDRPOINTER_REG_15_;
  assign n62549 = P2_P3_INSTADDRPOINTER_REG_13_ & n62548;
  assign n62550 = n62355 & n62549;
  assign n62551 = ~n62547 & ~n62550;
  assign n62552 = n59069 & n62551;
  assign n62553 = n62528 & n62545;
  assign n62554 = ~n62552 & n62553;
  assign n62555 = n59265 & ~n62521;
  assign n62556 = n59108 & ~n62521;
  assign n62557 = ~n62555 & ~n62556;
  assign n62558 = ~n59155 & ~n62521;
  assign n62559 = n59226 & ~n62532;
  assign n62560 = n59227 & ~n62532;
  assign n62561 = n60969 & ~n62521;
  assign n62562 = n59042 & ~n62532;
  assign n62563 = n60972 & ~n62521;
  assign n62564 = ~n62562 & ~n62563;
  assign n62565 = ~n62559 & ~n62560;
  assign n62566 = ~n62561 & n62565;
  assign n62567 = n62564 & n62566;
  assign n62568 = P2_P3_INSTADDRPOINTER_REG_14_ & ~n61896;
  assign n62569 = n62493 & ~n62568;
  assign n62570 = ~P2_P3_INSTADDRPOINTER_REG_14_ & n61896;
  assign n62571 = n62494 & ~n62570;
  assign n62572 = ~n62261 & n62571;
  assign n62573 = n62569 & ~n62572;
  assign n62574 = ~P2_P3_INSTADDRPOINTER_REG_15_ & ~n61896;
  assign n62575 = P2_P3_INSTADDRPOINTER_REG_15_ & n61896;
  assign n62576 = ~n62574 & ~n62575;
  assign n62577 = n62573 & ~n62576;
  assign n62578 = ~n62573 & n62576;
  assign n62579 = ~n62577 & ~n62578;
  assign n62580 = n61066 & ~n62579;
  assign n62581 = P2_P3_INSTADDRPOINTER_REG_14_ & n62405;
  assign n62582 = ~P2_P3_INSTADDRPOINTER_REG_15_ & ~n62581;
  assign n62583 = n62329 & n62549;
  assign n62584 = ~n62582 & ~n62583;
  assign n62585 = n61068 & n62584;
  assign n62586 = n62557 & ~n62558;
  assign n62587 = n62567 & n62586;
  assign n62588 = ~n62580 & n62587;
  assign n62589 = ~n62585 & n62588;
  assign n62590 = n62554 & n62589;
  assign n62591 = n60961 & ~n62590;
  assign n11116 = ~n62517 | n62591;
  assign n62593 = P2_P3_INSTADDRPOINTER_REG_16_ & n60960;
  assign n62594 = P2_P3_REIP_REG_16_ & n61105;
  assign n62595 = ~n62593 & ~n62594;
  assign n62596 = P2_P3_INSTADDRPOINTER_REG_15_ & n62518;
  assign n62597 = ~P2_P3_INSTADDRPOINTER_REG_16_ & n62596;
  assign n62598 = P2_P3_INSTADDRPOINTER_REG_16_ & ~n62596;
  assign n62599 = ~n62597 & ~n62598;
  assign n62600 = n61085 & ~n62599;
  assign n62601 = n59112 & ~n62599;
  assign n62602 = n61074 & ~n62599;
  assign n62603 = n61078 & ~n62599;
  assign n62604 = ~n62600 & ~n62601;
  assign n62605 = ~n62602 & n62604;
  assign n62606 = ~n62603 & n62605;
  assign n62607 = P2_P3_INSTADDRPOINTER_REG_15_ & n62529;
  assign n62608 = ~P2_P3_INSTADDRPOINTER_REG_16_ & n62607;
  assign n62609 = P2_P3_INSTADDRPOINTER_REG_16_ & ~n62607;
  assign n62610 = ~n62608 & ~n62609;
  assign n62611 = n58968 & ~n62610;
  assign n62612 = n59046 & ~n62610;
  assign n62613 = n59050 & ~n62610;
  assign n62614 = P2_P3_INSTADDRPOINTER_REG_15_ & n62536;
  assign n62615 = ~P2_P3_INSTADDRPOINTER_REG_16_ & n62614;
  assign n62616 = P2_P3_INSTADDRPOINTER_REG_16_ & ~n62614;
  assign n62617 = ~n62615 & ~n62616;
  assign n62618 = n59066 & ~n62617;
  assign n62619 = n59058 & ~n62617;
  assign n62620 = ~n62611 & ~n62612;
  assign n62621 = ~n62613 & n62620;
  assign n62622 = ~n62618 & n62621;
  assign n62623 = ~n62619 & n62622;
  assign n62624 = ~P2_P3_INSTADDRPOINTER_REG_16_ & n62550;
  assign n62625 = P2_P3_INSTADDRPOINTER_REG_16_ & ~n62550;
  assign n62626 = ~n62624 & ~n62625;
  assign n62627 = n59069 & ~n62626;
  assign n62628 = n62606 & n62623;
  assign n62629 = ~n62627 & n62628;
  assign n62630 = n59265 & ~n62599;
  assign n62631 = n59108 & ~n62599;
  assign n62632 = ~n62630 & ~n62631;
  assign n62633 = ~n59155 & ~n62599;
  assign n62634 = P2_P3_INSTADDRPOINTER_REG_15_ & ~n61896;
  assign n62635 = ~P2_P3_INSTADDRPOINTER_REG_15_ & n61896;
  assign n62636 = ~n62573 & ~n62635;
  assign n62637 = ~n62634 & ~n62636;
  assign n62638 = ~P2_P3_INSTADDRPOINTER_REG_16_ & ~n61896;
  assign n62639 = P2_P3_INSTADDRPOINTER_REG_16_ & n61896;
  assign n62640 = ~n62638 & ~n62639;
  assign n62641 = n62637 & ~n62640;
  assign n62642 = ~n62637 & n62640;
  assign n62643 = ~n62641 & ~n62642;
  assign n62644 = n61066 & ~n62643;
  assign n62645 = n59226 & ~n62610;
  assign n62646 = n59227 & ~n62610;
  assign n62647 = n60969 & ~n62599;
  assign n62648 = n59042 & ~n62610;
  assign n62649 = n60972 & ~n62599;
  assign n62650 = ~n62648 & ~n62649;
  assign n62651 = ~n62645 & ~n62646;
  assign n62652 = ~n62647 & n62651;
  assign n62653 = n62650 & n62652;
  assign n62654 = ~P2_P3_INSTADDRPOINTER_REG_16_ & n62583;
  assign n62655 = P2_P3_INSTADDRPOINTER_REG_16_ & ~n62583;
  assign n62656 = ~n62654 & ~n62655;
  assign n62657 = n61068 & ~n62656;
  assign n62658 = n62632 & ~n62633;
  assign n62659 = ~n62644 & n62658;
  assign n62660 = n62653 & n62659;
  assign n62661 = ~n62657 & n62660;
  assign n62662 = n62629 & n62661;
  assign n62663 = n60961 & ~n62662;
  assign n11121 = ~n62595 | n62663;
  assign n62665 = P2_P3_INSTADDRPOINTER_REG_17_ & n60960;
  assign n62666 = P2_P3_REIP_REG_17_ & n61105;
  assign n62667 = P2_P3_INSTADDRPOINTER_REG_16_ & n62607;
  assign n62668 = ~P2_P3_INSTADDRPOINTER_REG_17_ & n62667;
  assign n62669 = P2_P3_INSTADDRPOINTER_REG_17_ & ~n62667;
  assign n62670 = ~n62668 & ~n62669;
  assign n62671 = n59226 & ~n62670;
  assign n62672 = n59227 & ~n62670;
  assign n62673 = P2_P3_INSTADDRPOINTER_REG_16_ & n62596;
  assign n62674 = ~P2_P3_INSTADDRPOINTER_REG_17_ & n62673;
  assign n62675 = P2_P3_INSTADDRPOINTER_REG_17_ & ~n62673;
  assign n62676 = ~n62674 & ~n62675;
  assign n62677 = n60969 & ~n62676;
  assign n62678 = n59042 & ~n62670;
  assign n62679 = n60972 & ~n62676;
  assign n62680 = ~n62678 & ~n62679;
  assign n62681 = ~n62671 & ~n62672;
  assign n62682 = ~n62677 & n62681;
  assign n62683 = n62680 & n62682;
  assign n62684 = ~n59155 & ~n62676;
  assign n62685 = P2_P3_INSTADDRPOINTER_REG_16_ & P2_P3_INSTADDRPOINTER_REG_17_;
  assign n62686 = ~n62637 & n62685;
  assign n62687 = n61896 & ~n62686;
  assign n62688 = P2_P3_INSTADDRPOINTER_REG_17_ & ~n61896;
  assign n62689 = ~P2_P3_INSTADDRPOINTER_REG_16_ & ~n62634;
  assign n62690 = ~n62636 & n62689;
  assign n62691 = ~n62687 & ~n62688;
  assign n62692 = ~n62690 & n62691;
  assign n62693 = P2_P3_INSTADDRPOINTER_REG_17_ & n62690;
  assign n62694 = ~n61896 & ~n62693;
  assign n62695 = P2_P3_INSTADDRPOINTER_REG_17_ & n61896;
  assign n62696 = P2_P3_INSTADDRPOINTER_REG_16_ & ~n62637;
  assign n62697 = ~n62694 & ~n62695;
  assign n62698 = ~n62696 & n62697;
  assign n62699 = ~n62692 & ~n62698;
  assign n62700 = n61066 & n62699;
  assign n62701 = n59265 & ~n62676;
  assign n62702 = n59108 & ~n62676;
  assign n62703 = ~n62701 & ~n62702;
  assign n62704 = P2_P3_INSTADDRPOINTER_REG_16_ & n62583;
  assign n62705 = ~P2_P3_INSTADDRPOINTER_REG_17_ & ~n62704;
  assign n62706 = n62583 & n62685;
  assign n62707 = ~n62705 & ~n62706;
  assign n62708 = n61068 & n62707;
  assign n62709 = n62703 & ~n62708;
  assign n62710 = n61085 & ~n62676;
  assign n62711 = n59112 & ~n62676;
  assign n62712 = n61074 & ~n62676;
  assign n62713 = n61078 & ~n62676;
  assign n62714 = ~n62710 & ~n62711;
  assign n62715 = ~n62712 & n62714;
  assign n62716 = ~n62713 & n62715;
  assign n62717 = n58968 & ~n62670;
  assign n62718 = n59046 & ~n62670;
  assign n62719 = n59050 & ~n62670;
  assign n62720 = P2_P3_INSTADDRPOINTER_REG_16_ & n62614;
  assign n62721 = ~P2_P3_INSTADDRPOINTER_REG_17_ & n62720;
  assign n62722 = P2_P3_INSTADDRPOINTER_REG_17_ & ~n62720;
  assign n62723 = ~n62721 & ~n62722;
  assign n62724 = n59066 & ~n62723;
  assign n62725 = n59058 & ~n62723;
  assign n62726 = ~n62717 & ~n62718;
  assign n62727 = ~n62719 & n62726;
  assign n62728 = ~n62724 & n62727;
  assign n62729 = ~n62725 & n62728;
  assign n62730 = P2_P3_INSTADDRPOINTER_REG_16_ & n62550;
  assign n62731 = ~P2_P3_INSTADDRPOINTER_REG_17_ & ~n62730;
  assign n62732 = n62550 & n62685;
  assign n62733 = ~n62731 & ~n62732;
  assign n62734 = n59069 & n62733;
  assign n62735 = n62716 & n62729;
  assign n62736 = ~n62734 & n62735;
  assign n62737 = n62683 & ~n62684;
  assign n62738 = ~n62700 & n62737;
  assign n62739 = n62709 & n62738;
  assign n62740 = n62736 & n62739;
  assign n62741 = n60961 & ~n62740;
  assign n62742 = ~n62665 & ~n62666;
  assign n11126 = n62741 | ~n62742;
  assign n62744 = P2_P3_INSTADDRPOINTER_REG_18_ & n60960;
  assign n62745 = P2_P3_REIP_REG_18_ & n61105;
  assign n62746 = ~n62744 & ~n62745;
  assign n62747 = P2_P3_INSTADDRPOINTER_REG_17_ & n62673;
  assign n62748 = ~P2_P3_INSTADDRPOINTER_REG_18_ & n62747;
  assign n62749 = P2_P3_INSTADDRPOINTER_REG_18_ & ~n62747;
  assign n62750 = ~n62748 & ~n62749;
  assign n62751 = n61085 & ~n62750;
  assign n62752 = n59112 & ~n62750;
  assign n62753 = n61074 & ~n62750;
  assign n62754 = n61078 & ~n62750;
  assign n62755 = ~n62751 & ~n62752;
  assign n62756 = ~n62753 & n62755;
  assign n62757 = ~n62754 & n62756;
  assign n62758 = P2_P3_INSTADDRPOINTER_REG_17_ & n62667;
  assign n62759 = ~P2_P3_INSTADDRPOINTER_REG_18_ & n62758;
  assign n62760 = P2_P3_INSTADDRPOINTER_REG_18_ & ~n62758;
  assign n62761 = ~n62759 & ~n62760;
  assign n62762 = n58968 & ~n62761;
  assign n62763 = n59046 & ~n62761;
  assign n62764 = n59050 & ~n62761;
  assign n62765 = P2_P3_INSTADDRPOINTER_REG_17_ & n62720;
  assign n62766 = ~P2_P3_INSTADDRPOINTER_REG_18_ & n62765;
  assign n62767 = P2_P3_INSTADDRPOINTER_REG_18_ & ~n62765;
  assign n62768 = ~n62766 & ~n62767;
  assign n62769 = n59066 & ~n62768;
  assign n62770 = n59058 & ~n62768;
  assign n62771 = ~n62762 & ~n62763;
  assign n62772 = ~n62764 & n62771;
  assign n62773 = ~n62769 & n62772;
  assign n62774 = ~n62770 & n62773;
  assign n62775 = ~P2_P3_INSTADDRPOINTER_REG_18_ & n62732;
  assign n62776 = P2_P3_INSTADDRPOINTER_REG_18_ & ~n62732;
  assign n62777 = ~n62775 & ~n62776;
  assign n62778 = n59069 & ~n62777;
  assign n62779 = n62757 & n62774;
  assign n62780 = ~n62778 & n62779;
  assign n62781 = n59265 & ~n62750;
  assign n62782 = n59108 & ~n62750;
  assign n62783 = ~n62781 & ~n62782;
  assign n62784 = ~n59155 & ~n62750;
  assign n62785 = ~n61896 & ~n62690;
  assign n62786 = ~n62686 & ~n62785;
  assign n62787 = ~n62688 & n62786;
  assign n62788 = ~P2_P3_INSTADDRPOINTER_REG_18_ & ~n61896;
  assign n62789 = P2_P3_INSTADDRPOINTER_REG_18_ & n61896;
  assign n62790 = ~n62788 & ~n62789;
  assign n62791 = n62787 & ~n62790;
  assign n62792 = ~n62787 & n62790;
  assign n62793 = ~n62791 & ~n62792;
  assign n62794 = n61066 & ~n62793;
  assign n62795 = n59226 & ~n62761;
  assign n62796 = n59227 & ~n62761;
  assign n62797 = n60969 & ~n62750;
  assign n62798 = n59042 & ~n62761;
  assign n62799 = n60972 & ~n62750;
  assign n62800 = ~n62798 & ~n62799;
  assign n62801 = ~n62795 & ~n62796;
  assign n62802 = ~n62797 & n62801;
  assign n62803 = n62800 & n62802;
  assign n62804 = ~P2_P3_INSTADDRPOINTER_REG_18_ & n62706;
  assign n62805 = P2_P3_INSTADDRPOINTER_REG_18_ & ~n62706;
  assign n62806 = ~n62804 & ~n62805;
  assign n62807 = n61068 & ~n62806;
  assign n62808 = n62783 & ~n62784;
  assign n62809 = ~n62794 & n62808;
  assign n62810 = n62803 & n62809;
  assign n62811 = ~n62807 & n62810;
  assign n62812 = n62780 & n62811;
  assign n62813 = n60961 & ~n62812;
  assign n11131 = ~n62746 | n62813;
  assign n62815 = P2_P3_INSTADDRPOINTER_REG_19_ & n60960;
  assign n62816 = P2_P3_REIP_REG_19_ & n61105;
  assign n62817 = P2_P3_INSTADDRPOINTER_REG_18_ & n62758;
  assign n62818 = ~P2_P3_INSTADDRPOINTER_REG_19_ & n62817;
  assign n62819 = P2_P3_INSTADDRPOINTER_REG_19_ & ~n62817;
  assign n62820 = ~n62818 & ~n62819;
  assign n62821 = n59226 & ~n62820;
  assign n62822 = n59227 & ~n62820;
  assign n62823 = P2_P3_INSTADDRPOINTER_REG_18_ & n62747;
  assign n62824 = ~P2_P3_INSTADDRPOINTER_REG_19_ & n62823;
  assign n62825 = P2_P3_INSTADDRPOINTER_REG_19_ & ~n62823;
  assign n62826 = ~n62824 & ~n62825;
  assign n62827 = n60969 & ~n62826;
  assign n62828 = n59042 & ~n62820;
  assign n62829 = n60972 & ~n62826;
  assign n62830 = ~n62828 & ~n62829;
  assign n62831 = ~n62821 & ~n62822;
  assign n62832 = ~n62827 & n62831;
  assign n62833 = n62830 & n62832;
  assign n62834 = ~n59155 & ~n62826;
  assign n62835 = ~P2_P3_INSTADDRPOINTER_REG_19_ & ~n61896;
  assign n62836 = P2_P3_INSTADDRPOINTER_REG_19_ & n61896;
  assign n62837 = ~n62835 & ~n62836;
  assign n62838 = ~P2_P3_INSTADDRPOINTER_REG_18_ & n61896;
  assign n62839 = ~n62787 & ~n62838;
  assign n62840 = P2_P3_INSTADDRPOINTER_REG_18_ & ~n61896;
  assign n62841 = ~n62839 & ~n62840;
  assign n62842 = ~n62837 & n62841;
  assign n62843 = ~P2_P3_INSTADDRPOINTER_REG_19_ & n61896;
  assign n62844 = P2_P3_INSTADDRPOINTER_REG_19_ & ~n61896;
  assign n62845 = ~n62843 & ~n62844;
  assign n62846 = ~n62841 & ~n62845;
  assign n62847 = ~n62842 & ~n62846;
  assign n62848 = n61066 & ~n62847;
  assign n62849 = n59265 & ~n62826;
  assign n62850 = n59108 & ~n62826;
  assign n62851 = ~n62849 & ~n62850;
  assign n62852 = P2_P3_INSTADDRPOINTER_REG_18_ & n62706;
  assign n62853 = ~P2_P3_INSTADDRPOINTER_REG_19_ & ~n62852;
  assign n62854 = P2_P3_INSTADDRPOINTER_REG_18_ & P2_P3_INSTADDRPOINTER_REG_19_;
  assign n62855 = n62706 & n62854;
  assign n62856 = ~n62853 & ~n62855;
  assign n62857 = n61068 & n62856;
  assign n62858 = n62851 & ~n62857;
  assign n62859 = n61085 & ~n62826;
  assign n62860 = n59112 & ~n62826;
  assign n62861 = n61074 & ~n62826;
  assign n62862 = n61078 & ~n62826;
  assign n62863 = ~n62859 & ~n62860;
  assign n62864 = ~n62861 & n62863;
  assign n62865 = ~n62862 & n62864;
  assign n62866 = n58968 & ~n62820;
  assign n62867 = n59046 & ~n62820;
  assign n62868 = n59050 & ~n62820;
  assign n62869 = P2_P3_INSTADDRPOINTER_REG_18_ & n62765;
  assign n62870 = ~P2_P3_INSTADDRPOINTER_REG_19_ & n62869;
  assign n62871 = P2_P3_INSTADDRPOINTER_REG_19_ & ~n62869;
  assign n62872 = ~n62870 & ~n62871;
  assign n62873 = n59066 & ~n62872;
  assign n62874 = n59058 & ~n62872;
  assign n62875 = ~n62866 & ~n62867;
  assign n62876 = ~n62868 & n62875;
  assign n62877 = ~n62873 & n62876;
  assign n62878 = ~n62874 & n62877;
  assign n62879 = P2_P3_INSTADDRPOINTER_REG_18_ & n62732;
  assign n62880 = ~P2_P3_INSTADDRPOINTER_REG_19_ & ~n62879;
  assign n62881 = n62732 & n62854;
  assign n62882 = ~n62880 & ~n62881;
  assign n62883 = n59069 & n62882;
  assign n62884 = n62865 & n62878;
  assign n62885 = ~n62883 & n62884;
  assign n62886 = n62833 & ~n62834;
  assign n62887 = ~n62848 & n62886;
  assign n62888 = n62858 & n62887;
  assign n62889 = n62885 & n62888;
  assign n62890 = n60961 & ~n62889;
  assign n62891 = ~n62815 & ~n62816;
  assign n11136 = n62890 | ~n62891;
  assign n62893 = P2_P3_INSTADDRPOINTER_REG_20_ & n60960;
  assign n62894 = P2_P3_REIP_REG_20_ & n61105;
  assign n62895 = ~n62893 & ~n62894;
  assign n62896 = P2_P3_INSTADDRPOINTER_REG_19_ & P2_P3_INSTADDRPOINTER_REG_20_;
  assign n62897 = n61896 & ~n62896;
  assign n62898 = P2_P3_INSTADDRPOINTER_REG_20_ & ~n61896;
  assign n62899 = ~n62897 & ~n62898;
  assign n62900 = n62841 & ~n62844;
  assign n62901 = n62899 & ~n62900;
  assign n62902 = ~P2_P3_INSTADDRPOINTER_REG_19_ & n62841;
  assign n62903 = P2_P3_INSTADDRPOINTER_REG_20_ & n62902;
  assign n62904 = ~n61896 & ~n62903;
  assign n62905 = P2_P3_INSTADDRPOINTER_REG_20_ & n61896;
  assign n62906 = P2_P3_INSTADDRPOINTER_REG_19_ & ~n62841;
  assign n62907 = ~n62904 & ~n62905;
  assign n62908 = ~n62906 & n62907;
  assign n62909 = ~n62901 & ~n62908;
  assign n62910 = n61066 & n62909;
  assign n62911 = P2_P3_INSTADDRPOINTER_REG_19_ & n62823;
  assign n62912 = ~P2_P3_INSTADDRPOINTER_REG_20_ & n62911;
  assign n62913 = P2_P3_INSTADDRPOINTER_REG_20_ & ~n62911;
  assign n62914 = ~n62912 & ~n62913;
  assign n62915 = ~n59155 & ~n62914;
  assign n62916 = n59265 & ~n62914;
  assign n62917 = n59108 & ~n62914;
  assign n62918 = ~n62916 & ~n62917;
  assign n62919 = P2_P3_INSTADDRPOINTER_REG_19_ & n62817;
  assign n62920 = ~P2_P3_INSTADDRPOINTER_REG_20_ & n62919;
  assign n62921 = P2_P3_INSTADDRPOINTER_REG_20_ & ~n62919;
  assign n62922 = ~n62920 & ~n62921;
  assign n62923 = n59226 & ~n62922;
  assign n62924 = n59227 & ~n62922;
  assign n62925 = n60969 & ~n62914;
  assign n62926 = n59042 & ~n62922;
  assign n62927 = n60972 & ~n62914;
  assign n62928 = ~n62926 & ~n62927;
  assign n62929 = ~n62923 & ~n62924;
  assign n62930 = ~n62925 & n62929;
  assign n62931 = n62928 & n62930;
  assign n62932 = ~P2_P3_INSTADDRPOINTER_REG_20_ & ~n62855;
  assign n62933 = P2_P3_INSTADDRPOINTER_REG_20_ & n62855;
  assign n62934 = ~n62932 & ~n62933;
  assign n62935 = n61068 & n62934;
  assign n62936 = n61085 & ~n62914;
  assign n62937 = n59112 & ~n62914;
  assign n62938 = n61074 & ~n62914;
  assign n62939 = n61078 & ~n62914;
  assign n62940 = ~n62936 & ~n62937;
  assign n62941 = ~n62938 & n62940;
  assign n62942 = ~n62939 & n62941;
  assign n62943 = n58968 & ~n62922;
  assign n62944 = n59046 & ~n62922;
  assign n62945 = n59050 & ~n62922;
  assign n62946 = P2_P3_INSTADDRPOINTER_REG_19_ & n62869;
  assign n62947 = ~P2_P3_INSTADDRPOINTER_REG_20_ & n62946;
  assign n62948 = P2_P3_INSTADDRPOINTER_REG_20_ & ~n62946;
  assign n62949 = ~n62947 & ~n62948;
  assign n62950 = n59066 & ~n62949;
  assign n62951 = n59058 & ~n62949;
  assign n62952 = ~n62943 & ~n62944;
  assign n62953 = ~n62945 & n62952;
  assign n62954 = ~n62950 & n62953;
  assign n62955 = ~n62951 & n62954;
  assign n62956 = ~P2_P3_INSTADDRPOINTER_REG_20_ & ~n62881;
  assign n62957 = P2_P3_INSTADDRPOINTER_REG_20_ & n62881;
  assign n62958 = ~n62956 & ~n62957;
  assign n62959 = n59069 & n62958;
  assign n62960 = n62942 & n62955;
  assign n62961 = ~n62959 & n62960;
  assign n62962 = ~n62915 & n62918;
  assign n62963 = n62931 & n62962;
  assign n62964 = ~n62935 & n62963;
  assign n62965 = n62961 & n62964;
  assign n62966 = ~n62910 & n62965;
  assign n62967 = n60961 & ~n62966;
  assign n11141 = ~n62895 | n62967;
  assign n62969 = P2_P3_INSTADDRPOINTER_REG_21_ & n60960;
  assign n62970 = P2_P3_REIP_REG_21_ & n61105;
  assign n62971 = P2_P3_INSTADDRPOINTER_REG_20_ & n62911;
  assign n62972 = ~P2_P3_INSTADDRPOINTER_REG_21_ & n62971;
  assign n62973 = P2_P3_INSTADDRPOINTER_REG_21_ & ~n62971;
  assign n62974 = ~n62972 & ~n62973;
  assign n62975 = ~n59155 & ~n62974;
  assign n62976 = P2_P3_INSTADDRPOINTER_REG_20_ & n62919;
  assign n62977 = ~P2_P3_INSTADDRPOINTER_REG_21_ & n62976;
  assign n62978 = P2_P3_INSTADDRPOINTER_REG_21_ & ~n62976;
  assign n62979 = ~n62977 & ~n62978;
  assign n62980 = n59226 & ~n62979;
  assign n62981 = n59227 & ~n62979;
  assign n62982 = n60969 & ~n62974;
  assign n62983 = n59042 & ~n62979;
  assign n62984 = n60972 & ~n62974;
  assign n62985 = ~n62983 & ~n62984;
  assign n62986 = ~n62980 & ~n62981;
  assign n62987 = ~n62982 & n62986;
  assign n62988 = n62985 & n62987;
  assign n62989 = ~P2_P3_INSTADDRPOINTER_REG_21_ & ~n62933;
  assign n62990 = P2_P3_INSTADDRPOINTER_REG_21_ & n62933;
  assign n62991 = ~n62989 & ~n62990;
  assign n62992 = n61068 & n62991;
  assign n62993 = n58968 & ~n62979;
  assign n62994 = n59046 & ~n62979;
  assign n62995 = n59050 & ~n62979;
  assign n62996 = P2_P3_INSTADDRPOINTER_REG_20_ & n62946;
  assign n62997 = ~P2_P3_INSTADDRPOINTER_REG_21_ & n62996;
  assign n62998 = P2_P3_INSTADDRPOINTER_REG_21_ & ~n62996;
  assign n62999 = ~n62997 & ~n62998;
  assign n63000 = n59066 & ~n62999;
  assign n63001 = n59058 & ~n62999;
  assign n63002 = ~n62993 & ~n62994;
  assign n63003 = ~n62995 & n63002;
  assign n63004 = ~n63000 & n63003;
  assign n63005 = ~n63001 & n63004;
  assign n63006 = n61085 & ~n62974;
  assign n63007 = n59112 & ~n62974;
  assign n63008 = n61074 & ~n62974;
  assign n63009 = n61078 & ~n62974;
  assign n63010 = ~n63006 & ~n63007;
  assign n63011 = ~n63008 & n63010;
  assign n63012 = ~n63009 & n63011;
  assign n63013 = ~P2_P3_INSTADDRPOINTER_REG_21_ & ~n62957;
  assign n63014 = P2_P3_INSTADDRPOINTER_REG_20_ & P2_P3_INSTADDRPOINTER_REG_21_;
  assign n63015 = n62881 & n63014;
  assign n63016 = ~n63013 & ~n63015;
  assign n63017 = n59069 & n63016;
  assign n63018 = n63005 & n63012;
  assign n63019 = ~n63017 & n63018;
  assign n63020 = n59265 & ~n62974;
  assign n63021 = n59108 & ~n62974;
  assign n63022 = ~n63020 & ~n63021;
  assign n63023 = ~n62841 & n62896;
  assign n63024 = ~n62898 & ~n63023;
  assign n63025 = ~n61896 & ~n62902;
  assign n63026 = n63024 & ~n63025;
  assign n63027 = ~P2_P3_INSTADDRPOINTER_REG_21_ & ~n61896;
  assign n63028 = P2_P3_INSTADDRPOINTER_REG_21_ & n61896;
  assign n63029 = ~n63027 & ~n63028;
  assign n63030 = n63026 & ~n63029;
  assign n63031 = ~n63026 & n63029;
  assign n63032 = ~n63030 & ~n63031;
  assign n63033 = n61066 & ~n63032;
  assign n63034 = n63022 & ~n63033;
  assign n63035 = ~n62975 & n62988;
  assign n63036 = ~n62992 & n63035;
  assign n63037 = n63019 & n63036;
  assign n63038 = n63034 & n63037;
  assign n63039 = n60961 & ~n63038;
  assign n63040 = ~n62969 & ~n62970;
  assign n11146 = n63039 | ~n63040;
  assign n63042 = P2_P3_INSTADDRPOINTER_REG_22_ & n60960;
  assign n63043 = P2_P3_REIP_REG_22_ & n61105;
  assign n63044 = ~n63042 & ~n63043;
  assign n63045 = P2_P3_INSTADDRPOINTER_REG_21_ & n62996;
  assign n63046 = ~P2_P3_INSTADDRPOINTER_REG_22_ & n63045;
  assign n63047 = P2_P3_INSTADDRPOINTER_REG_22_ & ~n63045;
  assign n63048 = ~n63046 & ~n63047;
  assign n63049 = n59066 & ~n63048;
  assign n63050 = n59058 & ~n63048;
  assign n63051 = ~n63049 & ~n63050;
  assign n63052 = P2_P3_INSTADDRPOINTER_REG_21_ & n62976;
  assign n63053 = ~P2_P3_INSTADDRPOINTER_REG_22_ & n63052;
  assign n63054 = P2_P3_INSTADDRPOINTER_REG_22_ & ~n63052;
  assign n63055 = ~n63053 & ~n63054;
  assign n63056 = n58968 & ~n63055;
  assign n63057 = n59046 & ~n63055;
  assign n63058 = n59050 & ~n63055;
  assign n63059 = ~n63056 & ~n63057;
  assign n63060 = ~n63058 & n63059;
  assign n63061 = P2_P3_INSTADDRPOINTER_REG_21_ & n62971;
  assign n63062 = ~P2_P3_INSTADDRPOINTER_REG_22_ & n63061;
  assign n63063 = P2_P3_INSTADDRPOINTER_REG_22_ & ~n63061;
  assign n63064 = ~n63062 & ~n63063;
  assign n63065 = n61074 & ~n63064;
  assign n63066 = n61078 & ~n63064;
  assign n63067 = n59112 & ~n63064;
  assign n63068 = ~n63065 & ~n63066;
  assign n63069 = ~n63067 & n63068;
  assign n63070 = ~P2_P3_INSTADDRPOINTER_REG_22_ & n63015;
  assign n63071 = P2_P3_INSTADDRPOINTER_REG_22_ & ~n63015;
  assign n63072 = ~n63070 & ~n63071;
  assign n63073 = n59069 & ~n63072;
  assign n63074 = n61085 & ~n63064;
  assign n63075 = ~n63073 & ~n63074;
  assign n63076 = n63051 & n63060;
  assign n63077 = n63069 & n63076;
  assign n63078 = n63075 & n63077;
  assign n63079 = P2_P3_INSTADDRPOINTER_REG_21_ & n62896;
  assign n63080 = n61896 & ~n63079;
  assign n63081 = ~n62838 & ~n63080;
  assign n63082 = ~n62787 & n63081;
  assign n63083 = P2_P3_INSTADDRPOINTER_REG_21_ & ~n61896;
  assign n63084 = ~n62840 & ~n63083;
  assign n63085 = ~n62844 & n63084;
  assign n63086 = ~n62898 & n63085;
  assign n63087 = ~n63082 & n63086;
  assign n63088 = ~P2_P3_INSTADDRPOINTER_REG_22_ & ~n61896;
  assign n63089 = P2_P3_INSTADDRPOINTER_REG_22_ & n61896;
  assign n63090 = ~n63088 & ~n63089;
  assign n63091 = n63087 & ~n63090;
  assign n63092 = ~n63087 & n63090;
  assign n63093 = ~n63091 & ~n63092;
  assign n63094 = n61066 & ~n63093;
  assign n63095 = ~n59155 & ~n63064;
  assign n63096 = n59265 & ~n63064;
  assign n63097 = n59108 & ~n63064;
  assign n63098 = ~n63096 & ~n63097;
  assign n63099 = n59226 & ~n63055;
  assign n63100 = n59227 & ~n63055;
  assign n63101 = n60969 & ~n63064;
  assign n63102 = n59042 & ~n63055;
  assign n63103 = n60972 & ~n63064;
  assign n63104 = ~n63102 & ~n63103;
  assign n63105 = ~n63099 & ~n63100;
  assign n63106 = ~n63101 & n63105;
  assign n63107 = n63104 & n63106;
  assign n63108 = ~P2_P3_INSTADDRPOINTER_REG_22_ & n62990;
  assign n63109 = P2_P3_INSTADDRPOINTER_REG_22_ & ~n62990;
  assign n63110 = ~n63108 & ~n63109;
  assign n63111 = n61068 & ~n63110;
  assign n63112 = ~n63094 & ~n63095;
  assign n63113 = n63098 & n63112;
  assign n63114 = n63107 & n63113;
  assign n63115 = ~n63111 & n63114;
  assign n63116 = n63078 & n63115;
  assign n63117 = n60961 & ~n63116;
  assign n11151 = ~n63044 | n63117;
  assign n63119 = P2_P3_INSTADDRPOINTER_REG_23_ & n60960;
  assign n63120 = P2_P3_REIP_REG_23_ & n61105;
  assign n63121 = ~n63119 & ~n63120;
  assign n63122 = P2_P3_INSTADDRPOINTER_REG_22_ & n63045;
  assign n63123 = ~P2_P3_INSTADDRPOINTER_REG_23_ & n63122;
  assign n63124 = P2_P3_INSTADDRPOINTER_REG_23_ & ~n63122;
  assign n63125 = ~n63123 & ~n63124;
  assign n63126 = n59066 & ~n63125;
  assign n63127 = n59058 & ~n63125;
  assign n63128 = ~n63126 & ~n63127;
  assign n63129 = P2_P3_INSTADDRPOINTER_REG_22_ & n63052;
  assign n63130 = ~P2_P3_INSTADDRPOINTER_REG_23_ & n63129;
  assign n63131 = P2_P3_INSTADDRPOINTER_REG_23_ & ~n63129;
  assign n63132 = ~n63130 & ~n63131;
  assign n63133 = n58968 & ~n63132;
  assign n63134 = n59046 & ~n63132;
  assign n63135 = n59050 & ~n63132;
  assign n63136 = ~n63133 & ~n63134;
  assign n63137 = ~n63135 & n63136;
  assign n63138 = P2_P3_INSTADDRPOINTER_REG_22_ & n63061;
  assign n63139 = ~P2_P3_INSTADDRPOINTER_REG_23_ & n63138;
  assign n63140 = P2_P3_INSTADDRPOINTER_REG_23_ & ~n63138;
  assign n63141 = ~n63139 & ~n63140;
  assign n63142 = n61074 & ~n63141;
  assign n63143 = n61078 & ~n63141;
  assign n63144 = n59112 & ~n63141;
  assign n63145 = ~n63142 & ~n63143;
  assign n63146 = ~n63144 & n63145;
  assign n63147 = P2_P3_INSTADDRPOINTER_REG_22_ & n63015;
  assign n63148 = ~P2_P3_INSTADDRPOINTER_REG_23_ & ~n63147;
  assign n63149 = P2_P3_INSTADDRPOINTER_REG_22_ & P2_P3_INSTADDRPOINTER_REG_23_;
  assign n63150 = n63015 & n63149;
  assign n63151 = ~n63148 & ~n63150;
  assign n63152 = n59069 & n63151;
  assign n63153 = n61085 & ~n63141;
  assign n63154 = ~n63152 & ~n63153;
  assign n63155 = n63128 & n63137;
  assign n63156 = n63146 & n63155;
  assign n63157 = n63154 & n63156;
  assign n63158 = ~P2_P3_INSTADDRPOINTER_REG_22_ & n61896;
  assign n63159 = n63081 & ~n63158;
  assign n63160 = ~n62787 & n63159;
  assign n63161 = P2_P3_INSTADDRPOINTER_REG_22_ & ~n61896;
  assign n63162 = n63086 & ~n63161;
  assign n63163 = ~n63160 & n63162;
  assign n63164 = ~P2_P3_INSTADDRPOINTER_REG_23_ & ~n61896;
  assign n63165 = P2_P3_INSTADDRPOINTER_REG_23_ & n61896;
  assign n63166 = ~n63164 & ~n63165;
  assign n63167 = n63163 & ~n63166;
  assign n63168 = ~n63163 & n63166;
  assign n63169 = ~n63167 & ~n63168;
  assign n63170 = n61066 & ~n63169;
  assign n63171 = ~n59155 & ~n63141;
  assign n63172 = n59265 & ~n63141;
  assign n63173 = n59108 & ~n63141;
  assign n63174 = ~n63172 & ~n63173;
  assign n63175 = n59226 & ~n63132;
  assign n63176 = n59227 & ~n63132;
  assign n63177 = n60969 & ~n63141;
  assign n63178 = n59042 & ~n63132;
  assign n63179 = n60972 & ~n63141;
  assign n63180 = ~n63178 & ~n63179;
  assign n63181 = ~n63175 & ~n63176;
  assign n63182 = ~n63177 & n63181;
  assign n63183 = n63180 & n63182;
  assign n63184 = P2_P3_INSTADDRPOINTER_REG_22_ & n62990;
  assign n63185 = ~P2_P3_INSTADDRPOINTER_REG_23_ & ~n63184;
  assign n63186 = n62990 & n63149;
  assign n63187 = ~n63185 & ~n63186;
  assign n63188 = n61068 & n63187;
  assign n63189 = ~n63170 & ~n63171;
  assign n63190 = n63174 & n63189;
  assign n63191 = n63183 & n63190;
  assign n63192 = ~n63188 & n63191;
  assign n63193 = n63157 & n63192;
  assign n63194 = n60961 & ~n63193;
  assign n11156 = ~n63121 | n63194;
  assign n63196 = P2_P3_INSTADDRPOINTER_REG_24_ & n60960;
  assign n63197 = P2_P3_REIP_REG_24_ & n61105;
  assign n63198 = ~n63196 & ~n63197;
  assign n63199 = P2_P3_INSTADDRPOINTER_REG_23_ & n63122;
  assign n63200 = ~P2_P3_INSTADDRPOINTER_REG_24_ & n63199;
  assign n63201 = P2_P3_INSTADDRPOINTER_REG_24_ & ~n63199;
  assign n63202 = ~n63200 & ~n63201;
  assign n63203 = n59066 & ~n63202;
  assign n63204 = n59058 & ~n63202;
  assign n63205 = ~n63203 & ~n63204;
  assign n63206 = P2_P3_INSTADDRPOINTER_REG_23_ & n63129;
  assign n63207 = ~P2_P3_INSTADDRPOINTER_REG_24_ & n63206;
  assign n63208 = P2_P3_INSTADDRPOINTER_REG_24_ & ~n63206;
  assign n63209 = ~n63207 & ~n63208;
  assign n63210 = n58968 & ~n63209;
  assign n63211 = n59046 & ~n63209;
  assign n63212 = n59050 & ~n63209;
  assign n63213 = ~n63210 & ~n63211;
  assign n63214 = ~n63212 & n63213;
  assign n63215 = ~P2_P3_INSTADDRPOINTER_REG_24_ & n63150;
  assign n63216 = P2_P3_INSTADDRPOINTER_REG_24_ & ~n63150;
  assign n63217 = ~n63215 & ~n63216;
  assign n63218 = n59069 & ~n63217;
  assign n63219 = P2_P3_INSTADDRPOINTER_REG_23_ & n63138;
  assign n63220 = ~P2_P3_INSTADDRPOINTER_REG_24_ & n63219;
  assign n63221 = P2_P3_INSTADDRPOINTER_REG_24_ & ~n63219;
  assign n63222 = ~n63220 & ~n63221;
  assign n63223 = n61085 & ~n63222;
  assign n63224 = ~n63218 & ~n63223;
  assign n63225 = n61074 & ~n63222;
  assign n63226 = n61078 & ~n63222;
  assign n63227 = n59112 & ~n63222;
  assign n63228 = ~n63225 & ~n63226;
  assign n63229 = ~n63227 & n63228;
  assign n63230 = n63205 & n63214;
  assign n63231 = n63224 & n63230;
  assign n63232 = n63229 & n63231;
  assign n63233 = P2_P3_INSTADDRPOINTER_REG_23_ & ~n61896;
  assign n63234 = n63162 & ~n63233;
  assign n63235 = ~P2_P3_INSTADDRPOINTER_REG_23_ & n61896;
  assign n63236 = n63159 & ~n63235;
  assign n63237 = ~n62787 & n63236;
  assign n63238 = n63234 & ~n63237;
  assign n63239 = ~P2_P3_INSTADDRPOINTER_REG_24_ & ~n61896;
  assign n63240 = P2_P3_INSTADDRPOINTER_REG_24_ & n61896;
  assign n63241 = ~n63239 & ~n63240;
  assign n63242 = n63238 & ~n63241;
  assign n63243 = ~n63238 & n63241;
  assign n63244 = ~n63242 & ~n63243;
  assign n63245 = n61066 & ~n63244;
  assign n63246 = ~n59155 & ~n63222;
  assign n63247 = n59265 & ~n63222;
  assign n63248 = n59108 & ~n63222;
  assign n63249 = ~n63247 & ~n63248;
  assign n63250 = ~P2_P3_INSTADDRPOINTER_REG_24_ & n63186;
  assign n63251 = P2_P3_INSTADDRPOINTER_REG_24_ & ~n63186;
  assign n63252 = ~n63250 & ~n63251;
  assign n63253 = n61068 & ~n63252;
  assign n63254 = n59226 & ~n63209;
  assign n63255 = n59227 & ~n63209;
  assign n63256 = n60969 & ~n63222;
  assign n63257 = n59042 & ~n63209;
  assign n63258 = n60972 & ~n63222;
  assign n63259 = ~n63257 & ~n63258;
  assign n63260 = ~n63254 & ~n63255;
  assign n63261 = ~n63256 & n63260;
  assign n63262 = n63259 & n63261;
  assign n63263 = ~n63245 & ~n63246;
  assign n63264 = n63249 & n63263;
  assign n63265 = ~n63253 & n63264;
  assign n63266 = n63262 & n63265;
  assign n63267 = n63232 & n63266;
  assign n63268 = n60961 & ~n63267;
  assign n11161 = ~n63198 | n63268;
  assign n63270 = P2_P3_INSTADDRPOINTER_REG_25_ & n60960;
  assign n63271 = P2_P3_REIP_REG_25_ & n61105;
  assign n63272 = ~n63270 & ~n63271;
  assign n63273 = P2_P3_INSTADDRPOINTER_REG_24_ & n63199;
  assign n63274 = ~P2_P3_INSTADDRPOINTER_REG_25_ & n63273;
  assign n63275 = P2_P3_INSTADDRPOINTER_REG_25_ & ~n63273;
  assign n63276 = ~n63274 & ~n63275;
  assign n63277 = n59066 & ~n63276;
  assign n63278 = n59058 & ~n63276;
  assign n63279 = ~n63277 & ~n63278;
  assign n63280 = P2_P3_INSTADDRPOINTER_REG_24_ & n63206;
  assign n63281 = ~P2_P3_INSTADDRPOINTER_REG_25_ & n63280;
  assign n63282 = P2_P3_INSTADDRPOINTER_REG_25_ & ~n63280;
  assign n63283 = ~n63281 & ~n63282;
  assign n63284 = n58968 & ~n63283;
  assign n63285 = n59046 & ~n63283;
  assign n63286 = n59050 & ~n63283;
  assign n63287 = ~n63284 & ~n63285;
  assign n63288 = ~n63286 & n63287;
  assign n63289 = P2_P3_INSTADDRPOINTER_REG_24_ & n63150;
  assign n63290 = ~P2_P3_INSTADDRPOINTER_REG_25_ & ~n63289;
  assign n63291 = P2_P3_INSTADDRPOINTER_REG_24_ & P2_P3_INSTADDRPOINTER_REG_25_;
  assign n63292 = n63150 & n63291;
  assign n63293 = ~n63290 & ~n63292;
  assign n63294 = n59069 & n63293;
  assign n63295 = P2_P3_INSTADDRPOINTER_REG_24_ & n63219;
  assign n63296 = ~P2_P3_INSTADDRPOINTER_REG_25_ & n63295;
  assign n63297 = P2_P3_INSTADDRPOINTER_REG_25_ & ~n63295;
  assign n63298 = ~n63296 & ~n63297;
  assign n63299 = n61085 & ~n63298;
  assign n63300 = ~n63294 & ~n63299;
  assign n63301 = n61074 & ~n63298;
  assign n63302 = n61078 & ~n63298;
  assign n63303 = n59112 & ~n63298;
  assign n63304 = ~n63301 & ~n63302;
  assign n63305 = ~n63303 & n63304;
  assign n63306 = n63279 & n63288;
  assign n63307 = n63300 & n63306;
  assign n63308 = n63305 & n63307;
  assign n63309 = ~P2_P3_INSTADDRPOINTER_REG_25_ & ~n61896;
  assign n63310 = P2_P3_INSTADDRPOINTER_REG_25_ & n61896;
  assign n63311 = ~n63309 & ~n63310;
  assign n63312 = P2_P3_INSTADDRPOINTER_REG_24_ & ~n61896;
  assign n63313 = ~P2_P3_INSTADDRPOINTER_REG_24_ & n61896;
  assign n63314 = ~n63238 & ~n63313;
  assign n63315 = ~n63312 & ~n63314;
  assign n63316 = ~n63311 & n63315;
  assign n63317 = ~P2_P3_INSTADDRPOINTER_REG_25_ & n61896;
  assign n63318 = P2_P3_INSTADDRPOINTER_REG_25_ & ~n61896;
  assign n63319 = ~n63317 & ~n63318;
  assign n63320 = ~n63315 & ~n63319;
  assign n63321 = ~n63316 & ~n63320;
  assign n63322 = n61066 & ~n63321;
  assign n63323 = ~n59155 & ~n63298;
  assign n63324 = P2_P3_INSTADDRPOINTER_REG_24_ & n63186;
  assign n63325 = ~P2_P3_INSTADDRPOINTER_REG_25_ & ~n63324;
  assign n63326 = n63186 & n63291;
  assign n63327 = ~n63325 & ~n63326;
  assign n63328 = n61068 & n63327;
  assign n63329 = n59265 & ~n63298;
  assign n63330 = n59108 & ~n63298;
  assign n63331 = ~n63329 & ~n63330;
  assign n63332 = n59226 & ~n63283;
  assign n63333 = n59227 & ~n63283;
  assign n63334 = n60969 & ~n63298;
  assign n63335 = n59042 & ~n63283;
  assign n63336 = n60972 & ~n63298;
  assign n63337 = ~n63335 & ~n63336;
  assign n63338 = ~n63332 & ~n63333;
  assign n63339 = ~n63334 & n63338;
  assign n63340 = n63337 & n63339;
  assign n63341 = ~n63322 & ~n63323;
  assign n63342 = ~n63328 & n63341;
  assign n63343 = n63331 & n63342;
  assign n63344 = n63340 & n63343;
  assign n63345 = n63308 & n63344;
  assign n63346 = n60961 & ~n63345;
  assign n11166 = ~n63272 | n63346;
  assign n63348 = P2_P3_INSTADDRPOINTER_REG_26_ & n60960;
  assign n63349 = P2_P3_REIP_REG_26_ & n61105;
  assign n63350 = P2_P3_INSTADDRPOINTER_REG_26_ & ~n61896;
  assign n63351 = P2_P3_INSTADDRPOINTER_REG_25_ & P2_P3_INSTADDRPOINTER_REG_26_;
  assign n63352 = n61896 & ~n63351;
  assign n63353 = ~n63350 & ~n63352;
  assign n63354 = n63315 & ~n63318;
  assign n63355 = n63353 & ~n63354;
  assign n63356 = ~P2_P3_INSTADDRPOINTER_REG_26_ & ~n61896;
  assign n63357 = P2_P3_INSTADDRPOINTER_REG_26_ & n61896;
  assign n63358 = ~n63356 & ~n63357;
  assign n63359 = ~n63318 & n63358;
  assign n63360 = ~n63315 & ~n63317;
  assign n63361 = n63359 & ~n63360;
  assign n63362 = ~n63355 & ~n63361;
  assign n63363 = n61066 & n63362;
  assign n63364 = ~P2_P3_INSTADDRPOINTER_REG_26_ & ~n63326;
  assign n63365 = P2_P3_INSTADDRPOINTER_REG_26_ & n63326;
  assign n63366 = ~n63364 & ~n63365;
  assign n63367 = n61068 & n63366;
  assign n63368 = ~n63363 & ~n63367;
  assign n63369 = P2_P3_INSTADDRPOINTER_REG_25_ & n63295;
  assign n63370 = ~P2_P3_INSTADDRPOINTER_REG_26_ & n63369;
  assign n63371 = P2_P3_INSTADDRPOINTER_REG_26_ & ~n63369;
  assign n63372 = ~n63370 & ~n63371;
  assign n63373 = ~n59155 & ~n63372;
  assign n63374 = n59265 & ~n63372;
  assign n63375 = n59108 & ~n63372;
  assign n63376 = ~n63374 & ~n63375;
  assign n63377 = P2_P3_INSTADDRPOINTER_REG_25_ & n63280;
  assign n63378 = ~P2_P3_INSTADDRPOINTER_REG_26_ & n63377;
  assign n63379 = P2_P3_INSTADDRPOINTER_REG_26_ & ~n63377;
  assign n63380 = ~n63378 & ~n63379;
  assign n63381 = n59226 & ~n63380;
  assign n63382 = n59227 & ~n63380;
  assign n63383 = n60969 & ~n63372;
  assign n63384 = n59042 & ~n63380;
  assign n63385 = n60972 & ~n63372;
  assign n63386 = ~n63384 & ~n63385;
  assign n63387 = ~n63381 & ~n63382;
  assign n63388 = ~n63383 & n63387;
  assign n63389 = n63386 & n63388;
  assign n63390 = P2_P3_INSTADDRPOINTER_REG_25_ & n63273;
  assign n63391 = ~P2_P3_INSTADDRPOINTER_REG_26_ & n63390;
  assign n63392 = P2_P3_INSTADDRPOINTER_REG_26_ & ~n63390;
  assign n63393 = ~n63391 & ~n63392;
  assign n63394 = n59066 & ~n63393;
  assign n63395 = n59058 & ~n63393;
  assign n63396 = ~n63394 & ~n63395;
  assign n63397 = n58968 & ~n63380;
  assign n63398 = n59046 & ~n63380;
  assign n63399 = n59050 & ~n63380;
  assign n63400 = ~n63397 & ~n63398;
  assign n63401 = ~n63399 & n63400;
  assign n63402 = ~P2_P3_INSTADDRPOINTER_REG_26_ & ~n63292;
  assign n63403 = P2_P3_INSTADDRPOINTER_REG_26_ & n63292;
  assign n63404 = ~n63402 & ~n63403;
  assign n63405 = n59069 & n63404;
  assign n63406 = n61085 & ~n63372;
  assign n63407 = ~n63405 & ~n63406;
  assign n63408 = n61074 & ~n63372;
  assign n63409 = n61078 & ~n63372;
  assign n63410 = n59112 & ~n63372;
  assign n63411 = ~n63408 & ~n63409;
  assign n63412 = ~n63410 & n63411;
  assign n63413 = n63396 & n63401;
  assign n63414 = n63407 & n63413;
  assign n63415 = n63412 & n63414;
  assign n63416 = n63368 & ~n63373;
  assign n63417 = n63376 & n63416;
  assign n63418 = n63389 & n63417;
  assign n63419 = n63415 & n63418;
  assign n63420 = n60961 & ~n63419;
  assign n63421 = ~n63348 & ~n63349;
  assign n11171 = n63420 | ~n63421;
  assign n63423 = P2_P3_INSTADDRPOINTER_REG_27_ & n60960;
  assign n63424 = P2_P3_REIP_REG_27_ & n61105;
  assign n63425 = ~n63318 & ~n63350;
  assign n63426 = ~n63315 & ~n63352;
  assign n63427 = n63425 & ~n63426;
  assign n63428 = ~P2_P3_INSTADDRPOINTER_REG_27_ & ~n61896;
  assign n63429 = P2_P3_INSTADDRPOINTER_REG_27_ & n61896;
  assign n63430 = ~n63428 & ~n63429;
  assign n63431 = n63427 & ~n63430;
  assign n63432 = ~n63427 & n63430;
  assign n63433 = ~n63431 & ~n63432;
  assign n63434 = n61066 & ~n63433;
  assign n63435 = ~P2_P3_INSTADDRPOINTER_REG_27_ & n63365;
  assign n63436 = P2_P3_INSTADDRPOINTER_REG_27_ & ~n63365;
  assign n63437 = ~n63435 & ~n63436;
  assign n63438 = n61068 & ~n63437;
  assign n63439 = ~n63434 & ~n63438;
  assign n63440 = P2_P3_INSTADDRPOINTER_REG_26_ & n63369;
  assign n63441 = ~P2_P3_INSTADDRPOINTER_REG_27_ & n63440;
  assign n63442 = P2_P3_INSTADDRPOINTER_REG_27_ & ~n63440;
  assign n63443 = ~n63441 & ~n63442;
  assign n63444 = ~n59155 & ~n63443;
  assign n63445 = n59265 & ~n63443;
  assign n63446 = n59108 & ~n63443;
  assign n63447 = ~n63445 & ~n63446;
  assign n63448 = P2_P3_INSTADDRPOINTER_REG_26_ & n63377;
  assign n63449 = ~P2_P3_INSTADDRPOINTER_REG_27_ & n63448;
  assign n63450 = P2_P3_INSTADDRPOINTER_REG_27_ & ~n63448;
  assign n63451 = ~n63449 & ~n63450;
  assign n63452 = n59226 & ~n63451;
  assign n63453 = n59227 & ~n63451;
  assign n63454 = n60969 & ~n63443;
  assign n63455 = n59042 & ~n63451;
  assign n63456 = n60972 & ~n63443;
  assign n63457 = ~n63455 & ~n63456;
  assign n63458 = ~n63452 & ~n63453;
  assign n63459 = ~n63454 & n63458;
  assign n63460 = n63457 & n63459;
  assign n63461 = P2_P3_INSTADDRPOINTER_REG_26_ & n63390;
  assign n63462 = ~P2_P3_INSTADDRPOINTER_REG_27_ & n63461;
  assign n63463 = P2_P3_INSTADDRPOINTER_REG_27_ & ~n63461;
  assign n63464 = ~n63462 & ~n63463;
  assign n63465 = n59066 & ~n63464;
  assign n63466 = n59058 & ~n63464;
  assign n63467 = ~n63465 & ~n63466;
  assign n63468 = n58968 & ~n63451;
  assign n63469 = n59046 & ~n63451;
  assign n63470 = n59050 & ~n63451;
  assign n63471 = ~n63468 & ~n63469;
  assign n63472 = ~n63470 & n63471;
  assign n63473 = ~P2_P3_INSTADDRPOINTER_REG_27_ & n63403;
  assign n63474 = P2_P3_INSTADDRPOINTER_REG_27_ & ~n63403;
  assign n63475 = ~n63473 & ~n63474;
  assign n63476 = n59069 & ~n63475;
  assign n63477 = n61085 & ~n63443;
  assign n63478 = ~n63476 & ~n63477;
  assign n63479 = n61074 & ~n63443;
  assign n63480 = n61078 & ~n63443;
  assign n63481 = n59112 & ~n63443;
  assign n63482 = ~n63479 & ~n63480;
  assign n63483 = ~n63481 & n63482;
  assign n63484 = n63467 & n63472;
  assign n63485 = n63478 & n63484;
  assign n63486 = n63483 & n63485;
  assign n63487 = n63439 & ~n63444;
  assign n63488 = n63447 & n63487;
  assign n63489 = n63460 & n63488;
  assign n63490 = n63486 & n63489;
  assign n63491 = n60961 & ~n63490;
  assign n63492 = ~n63423 & ~n63424;
  assign n11176 = n63491 | ~n63492;
  assign n63494 = P2_P3_INSTADDRPOINTER_REG_28_ & n60960;
  assign n63495 = P2_P3_REIP_REG_28_ & n61105;
  assign n63496 = P2_P3_INSTADDRPOINTER_REG_27_ & P2_P3_INSTADDRPOINTER_REG_28_;
  assign n63497 = ~n63427 & n63496;
  assign n63498 = n61896 & ~n63497;
  assign n63499 = P2_P3_INSTADDRPOINTER_REG_28_ & ~n61896;
  assign n63500 = ~P2_P3_INSTADDRPOINTER_REG_27_ & ~n63318;
  assign n63501 = ~n63350 & n63500;
  assign n63502 = ~n63426 & n63501;
  assign n63503 = ~n63498 & ~n63499;
  assign n63504 = ~n63502 & n63503;
  assign n63505 = P2_P3_INSTADDRPOINTER_REG_28_ & n63502;
  assign n63506 = ~n61896 & ~n63505;
  assign n63507 = P2_P3_INSTADDRPOINTER_REG_28_ & n61896;
  assign n63508 = P2_P3_INSTADDRPOINTER_REG_27_ & ~n63427;
  assign n63509 = ~n63506 & ~n63507;
  assign n63510 = ~n63508 & n63509;
  assign n63511 = ~n63504 & ~n63510;
  assign n63512 = n61066 & n63511;
  assign n63513 = P2_P3_INSTADDRPOINTER_REG_27_ & n63365;
  assign n63514 = ~P2_P3_INSTADDRPOINTER_REG_28_ & ~n63513;
  assign n63515 = n63365 & n63496;
  assign n63516 = ~n63514 & ~n63515;
  assign n63517 = n61068 & n63516;
  assign n63518 = ~n63512 & ~n63517;
  assign n63519 = P2_P3_INSTADDRPOINTER_REG_27_ & n63440;
  assign n63520 = ~P2_P3_INSTADDRPOINTER_REG_28_ & n63519;
  assign n63521 = P2_P3_INSTADDRPOINTER_REG_28_ & ~n63519;
  assign n63522 = ~n63520 & ~n63521;
  assign n63523 = ~n59155 & ~n63522;
  assign n63524 = n59265 & ~n63522;
  assign n63525 = n59108 & ~n63522;
  assign n63526 = ~n63524 & ~n63525;
  assign n63527 = P2_P3_INSTADDRPOINTER_REG_27_ & n63448;
  assign n63528 = ~P2_P3_INSTADDRPOINTER_REG_28_ & n63527;
  assign n63529 = P2_P3_INSTADDRPOINTER_REG_28_ & ~n63527;
  assign n63530 = ~n63528 & ~n63529;
  assign n63531 = n59226 & ~n63530;
  assign n63532 = n59227 & ~n63530;
  assign n63533 = n60969 & ~n63522;
  assign n63534 = n59042 & ~n63530;
  assign n63535 = n60972 & ~n63522;
  assign n63536 = ~n63534 & ~n63535;
  assign n63537 = ~n63531 & ~n63532;
  assign n63538 = ~n63533 & n63537;
  assign n63539 = n63536 & n63538;
  assign n63540 = P2_P3_INSTADDRPOINTER_REG_27_ & n63461;
  assign n63541 = ~P2_P3_INSTADDRPOINTER_REG_28_ & n63540;
  assign n63542 = P2_P3_INSTADDRPOINTER_REG_28_ & ~n63540;
  assign n63543 = ~n63541 & ~n63542;
  assign n63544 = n59066 & ~n63543;
  assign n63545 = n59058 & ~n63543;
  assign n63546 = ~n63544 & ~n63545;
  assign n63547 = n58968 & ~n63530;
  assign n63548 = n59046 & ~n63530;
  assign n63549 = n59050 & ~n63530;
  assign n63550 = ~n63547 & ~n63548;
  assign n63551 = ~n63549 & n63550;
  assign n63552 = P2_P3_INSTADDRPOINTER_REG_27_ & n63403;
  assign n63553 = ~P2_P3_INSTADDRPOINTER_REG_28_ & ~n63552;
  assign n63554 = n63403 & n63496;
  assign n63555 = ~n63553 & ~n63554;
  assign n63556 = n59069 & n63555;
  assign n63557 = n61085 & ~n63522;
  assign n63558 = ~n63556 & ~n63557;
  assign n63559 = n61074 & ~n63522;
  assign n63560 = n61078 & ~n63522;
  assign n63561 = n59112 & ~n63522;
  assign n63562 = ~n63559 & ~n63560;
  assign n63563 = ~n63561 & n63562;
  assign n63564 = n63546 & n63551;
  assign n63565 = n63558 & n63564;
  assign n63566 = n63563 & n63565;
  assign n63567 = n63518 & ~n63523;
  assign n63568 = n63526 & n63567;
  assign n63569 = n63539 & n63568;
  assign n63570 = n63566 & n63569;
  assign n63571 = n60961 & ~n63570;
  assign n63572 = ~n63494 & ~n63495;
  assign n11181 = n63571 | ~n63572;
  assign n63574 = P2_P3_INSTADDRPOINTER_REG_29_ & n60960;
  assign n63575 = P2_P3_REIP_REG_29_ & n61105;
  assign n63576 = ~n61896 & ~n63502;
  assign n63577 = ~n63499 & ~n63576;
  assign n63578 = ~n63497 & n63577;
  assign n63579 = ~P2_P3_INSTADDRPOINTER_REG_29_ & ~n61896;
  assign n63580 = P2_P3_INSTADDRPOINTER_REG_29_ & n61896;
  assign n63581 = ~n63579 & ~n63580;
  assign n63582 = n63578 & ~n63581;
  assign n63583 = ~n63578 & n63581;
  assign n63584 = ~n63582 & ~n63583;
  assign n63585 = n61066 & ~n63584;
  assign n63586 = ~P2_P3_INSTADDRPOINTER_REG_29_ & ~n63515;
  assign n63587 = P2_P3_INSTADDRPOINTER_REG_29_ & n63515;
  assign n63588 = ~n63586 & ~n63587;
  assign n63589 = n61068 & n63588;
  assign n63590 = ~n63585 & ~n63589;
  assign n63591 = P2_P3_INSTADDRPOINTER_REG_28_ & n63519;
  assign n63592 = ~P2_P3_INSTADDRPOINTER_REG_29_ & n63591;
  assign n63593 = P2_P3_INSTADDRPOINTER_REG_29_ & ~n63591;
  assign n63594 = ~n63592 & ~n63593;
  assign n63595 = ~n59155 & ~n63594;
  assign n63596 = n59265 & ~n63594;
  assign n63597 = n59108 & ~n63594;
  assign n63598 = ~n63596 & ~n63597;
  assign n63599 = P2_P3_INSTADDRPOINTER_REG_28_ & n63527;
  assign n63600 = ~P2_P3_INSTADDRPOINTER_REG_29_ & n63599;
  assign n63601 = P2_P3_INSTADDRPOINTER_REG_29_ & ~n63599;
  assign n63602 = ~n63600 & ~n63601;
  assign n63603 = n59226 & ~n63602;
  assign n63604 = n59227 & ~n63602;
  assign n63605 = n60969 & ~n63594;
  assign n63606 = n59042 & ~n63602;
  assign n63607 = n60972 & ~n63594;
  assign n63608 = ~n63606 & ~n63607;
  assign n63609 = ~n63603 & ~n63604;
  assign n63610 = ~n63605 & n63609;
  assign n63611 = n63608 & n63610;
  assign n63612 = P2_P3_INSTADDRPOINTER_REG_28_ & n63540;
  assign n63613 = ~P2_P3_INSTADDRPOINTER_REG_29_ & n63612;
  assign n63614 = P2_P3_INSTADDRPOINTER_REG_29_ & ~n63612;
  assign n63615 = ~n63613 & ~n63614;
  assign n63616 = n59066 & ~n63615;
  assign n63617 = n59058 & ~n63615;
  assign n63618 = ~n63616 & ~n63617;
  assign n63619 = n58968 & ~n63602;
  assign n63620 = n59046 & ~n63602;
  assign n63621 = n59050 & ~n63602;
  assign n63622 = ~n63619 & ~n63620;
  assign n63623 = ~n63621 & n63622;
  assign n63624 = ~P2_P3_INSTADDRPOINTER_REG_29_ & ~n63554;
  assign n63625 = P2_P3_INSTADDRPOINTER_REG_29_ & n63554;
  assign n63626 = ~n63624 & ~n63625;
  assign n63627 = n59069 & n63626;
  assign n63628 = n61085 & ~n63594;
  assign n63629 = ~n63627 & ~n63628;
  assign n63630 = n61074 & ~n63594;
  assign n63631 = n61078 & ~n63594;
  assign n63632 = n59112 & ~n63594;
  assign n63633 = ~n63630 & ~n63631;
  assign n63634 = ~n63632 & n63633;
  assign n63635 = n63618 & n63623;
  assign n63636 = n63629 & n63635;
  assign n63637 = n63634 & n63636;
  assign n63638 = n63590 & ~n63595;
  assign n63639 = n63598 & n63638;
  assign n63640 = n63611 & n63639;
  assign n63641 = n63637 & n63640;
  assign n63642 = n60961 & ~n63641;
  assign n63643 = ~n63574 & ~n63575;
  assign n11186 = n63642 | ~n63643;
  assign n63645 = P2_P3_INSTADDRPOINTER_REG_30_ & n60960;
  assign n63646 = P2_P3_REIP_REG_30_ & n61105;
  assign n63647 = ~P2_P3_INSTADDRPOINTER_REG_30_ & ~n61896;
  assign n63648 = P2_P3_INSTADDRPOINTER_REG_30_ & n61896;
  assign n63649 = ~n63647 & ~n63648;
  assign n63650 = P2_P3_INSTADDRPOINTER_REG_29_ & ~n61896;
  assign n63651 = ~P2_P3_INSTADDRPOINTER_REG_29_ & n61896;
  assign n63652 = ~n63578 & ~n63651;
  assign n63653 = ~n63650 & ~n63652;
  assign n63654 = ~n63649 & n63653;
  assign n63655 = n63649 & ~n63653;
  assign n63656 = ~n63654 & ~n63655;
  assign n63657 = n61066 & ~n63656;
  assign n63658 = ~P2_P3_INSTADDRPOINTER_REG_30_ & n63587;
  assign n63659 = P2_P3_INSTADDRPOINTER_REG_30_ & ~n63587;
  assign n63660 = ~n63658 & ~n63659;
  assign n63661 = n61068 & ~n63660;
  assign n63662 = ~n63657 & ~n63661;
  assign n63663 = P2_P3_INSTADDRPOINTER_REG_29_ & n63591;
  assign n63664 = ~P2_P3_INSTADDRPOINTER_REG_30_ & n63663;
  assign n63665 = P2_P3_INSTADDRPOINTER_REG_30_ & ~n63663;
  assign n63666 = ~n63664 & ~n63665;
  assign n63667 = ~n59155 & ~n63666;
  assign n63668 = n59265 & ~n63666;
  assign n63669 = n59108 & ~n63666;
  assign n63670 = ~n63668 & ~n63669;
  assign n63671 = P2_P3_INSTADDRPOINTER_REG_29_ & n63599;
  assign n63672 = ~P2_P3_INSTADDRPOINTER_REG_30_ & n63671;
  assign n63673 = P2_P3_INSTADDRPOINTER_REG_30_ & ~n63671;
  assign n63674 = ~n63672 & ~n63673;
  assign n63675 = n59226 & ~n63674;
  assign n63676 = n59227 & ~n63674;
  assign n63677 = n60969 & ~n63666;
  assign n63678 = n59042 & ~n63674;
  assign n63679 = n60972 & ~n63666;
  assign n63680 = ~n63678 & ~n63679;
  assign n63681 = ~n63675 & ~n63676;
  assign n63682 = ~n63677 & n63681;
  assign n63683 = n63680 & n63682;
  assign n63684 = P2_P3_INSTADDRPOINTER_REG_29_ & n63612;
  assign n63685 = ~P2_P3_INSTADDRPOINTER_REG_30_ & n63684;
  assign n63686 = P2_P3_INSTADDRPOINTER_REG_30_ & ~n63684;
  assign n63687 = ~n63685 & ~n63686;
  assign n63688 = n59066 & ~n63687;
  assign n63689 = n59058 & ~n63687;
  assign n63690 = ~n63688 & ~n63689;
  assign n63691 = n58968 & ~n63674;
  assign n63692 = n59046 & ~n63674;
  assign n63693 = n59050 & ~n63674;
  assign n63694 = ~n63691 & ~n63692;
  assign n63695 = ~n63693 & n63694;
  assign n63696 = ~P2_P3_INSTADDRPOINTER_REG_30_ & n63625;
  assign n63697 = P2_P3_INSTADDRPOINTER_REG_30_ & ~n63625;
  assign n63698 = ~n63696 & ~n63697;
  assign n63699 = n59069 & ~n63698;
  assign n63700 = n61085 & ~n63666;
  assign n63701 = ~n63699 & ~n63700;
  assign n63702 = n61074 & ~n63666;
  assign n63703 = n61078 & ~n63666;
  assign n63704 = n59112 & ~n63666;
  assign n63705 = ~n63702 & ~n63703;
  assign n63706 = ~n63704 & n63705;
  assign n63707 = n63690 & n63695;
  assign n63708 = n63701 & n63707;
  assign n63709 = n63706 & n63708;
  assign n63710 = n63662 & ~n63667;
  assign n63711 = n63670 & n63710;
  assign n63712 = n63683 & n63711;
  assign n63713 = n63709 & n63712;
  assign n63714 = n60961 & ~n63713;
  assign n63715 = ~n63645 & ~n63646;
  assign n11191 = n63714 | ~n63715;
  assign n63717 = P2_P3_INSTADDRPOINTER_REG_31_ & n60960;
  assign n63718 = P2_P3_REIP_REG_31_ & n61105;
  assign n63719 = P2_P3_INSTADDRPOINTER_REG_30_ & n63625;
  assign n63720 = ~P2_P3_INSTADDRPOINTER_REG_31_ & n63719;
  assign n63721 = P2_P3_INSTADDRPOINTER_REG_31_ & ~n63719;
  assign n63722 = ~n63720 & ~n63721;
  assign n63723 = n59069 & ~n63722;
  assign n63724 = P2_P3_INSTADDRPOINTER_REG_30_ & n63663;
  assign n63725 = ~P2_P3_INSTADDRPOINTER_REG_31_ & n63724;
  assign n63726 = P2_P3_INSTADDRPOINTER_REG_31_ & ~n63724;
  assign n63727 = ~n63725 & ~n63726;
  assign n63728 = n61085 & ~n63727;
  assign n63729 = n59112 & ~n63727;
  assign n63730 = ~n63728 & ~n63729;
  assign n63731 = P2_P3_INSTADDRPOINTER_REG_30_ & n63671;
  assign n63732 = ~P2_P3_INSTADDRPOINTER_REG_31_ & n63731;
  assign n63733 = P2_P3_INSTADDRPOINTER_REG_31_ & ~n63731;
  assign n63734 = ~n63732 & ~n63733;
  assign n63735 = n59050 & ~n63734;
  assign n63736 = n58968 & ~n63734;
  assign n63737 = P2_P3_INSTADDRPOINTER_REG_30_ & n63684;
  assign n63738 = ~P2_P3_INSTADDRPOINTER_REG_31_ & n63737;
  assign n63739 = P2_P3_INSTADDRPOINTER_REG_31_ & ~n63737;
  assign n63740 = ~n63738 & ~n63739;
  assign n63741 = n59058 & ~n63740;
  assign n63742 = ~n63735 & ~n63736;
  assign n63743 = ~n63741 & n63742;
  assign n63744 = n61074 & ~n63727;
  assign n63745 = n61078 & ~n63727;
  assign n63746 = n59066 & ~n63740;
  assign n63747 = ~n63745 & ~n63746;
  assign n63748 = n63743 & ~n63744;
  assign n63749 = n63747 & n63748;
  assign n63750 = ~n63717 & ~n63718;
  assign n63751 = ~n63723 & n63750;
  assign n63752 = n63730 & n63751;
  assign n63753 = n63749 & n63752;
  assign n63754 = P2_P3_INSTADDRPOINTER_REG_30_ & P2_P3_INSTADDRPOINTER_REG_31_;
  assign n63755 = ~n63653 & n63754;
  assign n63756 = n61896 & ~n63755;
  assign n63757 = P2_P3_INSTADDRPOINTER_REG_31_ & ~n61896;
  assign n63758 = ~P2_P3_INSTADDRPOINTER_REG_30_ & n63653;
  assign n63759 = ~n63756 & ~n63757;
  assign n63760 = ~n63758 & n63759;
  assign n63761 = ~P2_P3_INSTADDRPOINTER_REG_30_ & P2_P3_INSTADDRPOINTER_REG_31_;
  assign n63762 = ~n63650 & n63761;
  assign n63763 = ~n63652 & n63762;
  assign n63764 = ~n61896 & ~n63763;
  assign n63765 = P2_P3_INSTADDRPOINTER_REG_31_ & n61896;
  assign n63766 = P2_P3_INSTADDRPOINTER_REG_30_ & ~n63653;
  assign n63767 = ~n63764 & ~n63765;
  assign n63768 = ~n63766 & n63767;
  assign n63769 = ~n63760 & ~n63768;
  assign n63770 = n61066 & n63769;
  assign n63771 = P2_P3_INSTADDRPOINTER_REG_30_ & n63587;
  assign n63772 = ~P2_P3_INSTADDRPOINTER_REG_31_ & n63771;
  assign n63773 = P2_P3_INSTADDRPOINTER_REG_31_ & ~n63771;
  assign n63774 = ~n63772 & ~n63773;
  assign n63775 = n61068 & ~n63774;
  assign n63776 = ~n63770 & ~n63775;
  assign n63777 = ~n59155 & ~n63727;
  assign n63778 = n59265 & ~n63727;
  assign n63779 = n59108 & ~n63727;
  assign n63780 = ~n63778 & ~n63779;
  assign n63781 = n59227 & ~n63734;
  assign n63782 = n63780 & ~n63781;
  assign n63783 = n60969 & ~n63727;
  assign n63784 = n59226 & ~n63734;
  assign n63785 = n59046 & ~n63734;
  assign n63786 = n59042 & ~n63734;
  assign n63787 = n60972 & ~n63727;
  assign n63788 = ~n63785 & ~n63786;
  assign n63789 = ~n63787 & n63788;
  assign n63790 = ~n63783 & ~n63784;
  assign n63791 = n63789 & n63790;
  assign n63792 = n63776 & ~n63777;
  assign n63793 = n63782 & n63792;
  assign n63794 = n63791 & n63793;
  assign n63795 = n63753 & n63794;
  assign n63796 = ~n60961 & ~n63717;
  assign n63797 = ~n63718 & n63796;
  assign n11196 = ~n63795 & ~n63797;
  assign n63799 = P2_P3_STATE2_REG_0_ & ~n58935;
  assign n63800 = ~P2_P3_STATE2_REG_0_ & ~n60928;
  assign n63801 = n59069 & n59072;
  assign n63802 = n59074 & n59078;
  assign n63803 = ~n63801 & ~n63802;
  assign n63804 = n59321 & ~n63803;
  assign n63805 = ~n63800 & ~n63804;
  assign n63806 = n63799 & ~n63805;
  assign n63807 = ~n61065 & n63806;
  assign n63808 = ~n61034 & n63807;
  assign n63809 = n61065 & n63806;
  assign n63810 = ~n61034 & n63809;
  assign n63811 = P2_P3_STATE2_REG_1_ & ~n63805;
  assign n63812 = P2_P3_STATEBS16_REG & n63811;
  assign n63813 = P2_P3_PHYADDRPOINTER_REG_0_ & n63812;
  assign n63814 = ~P2_P3_STATEBS16_REG & n63811;
  assign n63815 = P2_P3_PHYADDRPOINTER_REG_0_ & n63814;
  assign n63816 = P2_P3_PHYADDRPOINTER_REG_0_ & n63805;
  assign n63817 = P2_P3_STATE2_REG_0_ & n58935;
  assign n63818 = ~n63805 & n63817;
  assign n63819 = ~n61082 & n63818;
  assign n63820 = P2_P3_STATE2_REG_2_ & ~P2_P3_STATE2_REG_0_;
  assign n63821 = ~n63805 & n63820;
  assign n63822 = P2_P3_PHYADDRPOINTER_REG_0_ & n63821;
  assign n63823 = n59337 & ~n63805;
  assign n63824 = P2_P3_REIP_REG_0_ & n63823;
  assign n63825 = ~n63816 & ~n63819;
  assign n63826 = ~n63822 & n63825;
  assign n63827 = ~n63824 & n63826;
  assign n63828 = ~n63808 & ~n63810;
  assign n63829 = ~n63813 & n63828;
  assign n63830 = ~n63815 & n63829;
  assign n11201 = ~n63827 | ~n63830;
  assign n63832 = ~n61206 & n63807;
  assign n63833 = ~n61156 & n63809;
  assign n63834 = P2_P3_PHYADDRPOINTER_REG_1_ & n63812;
  assign n63835 = ~P2_P3_PHYADDRPOINTER_REG_1_ & n63814;
  assign n63836 = P2_P3_PHYADDRPOINTER_REG_1_ & n63805;
  assign n63837 = ~n61186 & n63818;
  assign n63838 = ~P2_P3_PHYADDRPOINTER_REG_1_ & n63821;
  assign n63839 = P2_P3_REIP_REG_1_ & n63823;
  assign n63840 = ~n63836 & ~n63837;
  assign n63841 = ~n63838 & n63840;
  assign n63842 = ~n63839 & n63841;
  assign n63843 = ~n63832 & ~n63833;
  assign n63844 = ~n63834 & n63843;
  assign n63845 = ~n63835 & n63844;
  assign n11206 = ~n63842 | ~n63845;
  assign n63847 = ~n61291 & n63807;
  assign n63848 = ~n61278 & n63809;
  assign n63849 = ~P2_P3_PHYADDRPOINTER_REG_2_ & n63812;
  assign n63850 = P2_P3_PHYADDRPOINTER_REG_1_ & ~P2_P3_PHYADDRPOINTER_REG_2_;
  assign n63851 = ~P2_P3_PHYADDRPOINTER_REG_1_ & P2_P3_PHYADDRPOINTER_REG_2_;
  assign n63852 = ~n63850 & ~n63851;
  assign n63853 = n63814 & ~n63852;
  assign n63854 = n63821 & ~n63852;
  assign n63855 = P2_P3_REIP_REG_2_ & n63823;
  assign n63856 = P2_P3_PHYADDRPOINTER_REG_2_ & n63805;
  assign n63857 = ~n61328 & n63818;
  assign n63858 = ~n63854 & ~n63855;
  assign n63859 = ~n63856 & n63858;
  assign n63860 = ~n63857 & n63859;
  assign n63861 = ~n63847 & ~n63848;
  assign n63862 = ~n63849 & n63861;
  assign n63863 = ~n63853 & n63862;
  assign n11211 = ~n63860 | ~n63863;
  assign n63865 = ~n61406 & n63807;
  assign n63866 = n61421 & n63809;
  assign n63867 = P2_P3_PHYADDRPOINTER_REG_2_ & ~P2_P3_PHYADDRPOINTER_REG_3_;
  assign n63868 = ~P2_P3_PHYADDRPOINTER_REG_2_ & P2_P3_PHYADDRPOINTER_REG_3_;
  assign n63869 = ~n63867 & ~n63868;
  assign n63870 = n63812 & ~n63869;
  assign n63871 = P2_P3_PHYADDRPOINTER_REG_1_ & P2_P3_PHYADDRPOINTER_REG_2_;
  assign n63872 = ~P2_P3_PHYADDRPOINTER_REG_3_ & n63871;
  assign n63873 = P2_P3_PHYADDRPOINTER_REG_3_ & ~n63871;
  assign n63874 = ~n63872 & ~n63873;
  assign n63875 = n63814 & ~n63874;
  assign n63876 = n63821 & ~n63874;
  assign n63877 = P2_P3_REIP_REG_3_ & n63823;
  assign n63878 = P2_P3_PHYADDRPOINTER_REG_3_ & n63805;
  assign n63879 = n61459 & n63818;
  assign n63880 = ~n63876 & ~n63877;
  assign n63881 = ~n63878 & n63880;
  assign n63882 = ~n63879 & n63881;
  assign n63883 = ~n63865 & ~n63866;
  assign n63884 = ~n63870 & n63883;
  assign n63885 = ~n63875 & n63884;
  assign n11216 = ~n63882 | ~n63885;
  assign n63887 = P2_P3_PHYADDRPOINTER_REG_2_ & P2_P3_PHYADDRPOINTER_REG_3_;
  assign n63888 = ~P2_P3_PHYADDRPOINTER_REG_4_ & n63887;
  assign n63889 = P2_P3_PHYADDRPOINTER_REG_4_ & ~n63887;
  assign n63890 = ~n63888 & ~n63889;
  assign n63891 = n63812 & ~n63890;
  assign n63892 = P2_P3_PHYADDRPOINTER_REG_3_ & n63871;
  assign n63893 = ~P2_P3_PHYADDRPOINTER_REG_4_ & n63892;
  assign n63894 = P2_P3_PHYADDRPOINTER_REG_4_ & ~n63892;
  assign n63895 = ~n63893 & ~n63894;
  assign n63896 = n63814 & ~n63895;
  assign n63897 = n61534 & n63809;
  assign n63898 = ~n61556 & n63807;
  assign n63899 = n63821 & ~n63895;
  assign n63900 = P2_P3_REIP_REG_4_ & n63823;
  assign n63901 = P2_P3_PHYADDRPOINTER_REG_4_ & n63805;
  assign n63902 = ~n61595 & n63818;
  assign n63903 = ~n63899 & ~n63900;
  assign n63904 = ~n63901 & n63903;
  assign n63905 = ~n63902 & n63904;
  assign n63906 = ~n63891 & ~n63896;
  assign n63907 = ~n63897 & n63906;
  assign n63908 = ~n63898 & n63907;
  assign n11221 = ~n63905 | ~n63908;
  assign n63910 = P2_P3_PHYADDRPOINTER_REG_4_ & n63887;
  assign n63911 = ~P2_P3_PHYADDRPOINTER_REG_5_ & n63910;
  assign n63912 = P2_P3_PHYADDRPOINTER_REG_5_ & ~n63910;
  assign n63913 = ~n63911 & ~n63912;
  assign n63914 = n63812 & ~n63913;
  assign n63915 = P2_P3_PHYADDRPOINTER_REG_4_ & n63892;
  assign n63916 = ~P2_P3_PHYADDRPOINTER_REG_5_ & n63915;
  assign n63917 = P2_P3_PHYADDRPOINTER_REG_5_ & ~n63915;
  assign n63918 = ~n63916 & ~n63917;
  assign n63919 = n63814 & ~n63918;
  assign n63920 = ~n61671 & n63807;
  assign n63921 = ~n61689 & n63809;
  assign n63922 = n63821 & ~n63918;
  assign n63923 = P2_P3_REIP_REG_5_ & n63823;
  assign n63924 = P2_P3_PHYADDRPOINTER_REG_5_ & n63805;
  assign n63925 = n61728 & n63818;
  assign n63926 = ~n63922 & ~n63923;
  assign n63927 = ~n63924 & n63926;
  assign n63928 = ~n63925 & n63927;
  assign n63929 = ~n63914 & ~n63919;
  assign n63930 = ~n63920 & n63929;
  assign n63931 = ~n63921 & n63930;
  assign n11226 = ~n63928 | ~n63931;
  assign n63933 = P2_P3_PHYADDRPOINTER_REG_5_ & n63910;
  assign n63934 = ~P2_P3_PHYADDRPOINTER_REG_6_ & n63933;
  assign n63935 = P2_P3_PHYADDRPOINTER_REG_6_ & ~n63933;
  assign n63936 = ~n63934 & ~n63935;
  assign n63937 = n63812 & ~n63936;
  assign n63938 = P2_P3_PHYADDRPOINTER_REG_5_ & n63915;
  assign n63939 = ~P2_P3_PHYADDRPOINTER_REG_6_ & n63938;
  assign n63940 = P2_P3_PHYADDRPOINTER_REG_6_ & ~n63938;
  assign n63941 = ~n63939 & ~n63940;
  assign n63942 = n63814 & ~n63941;
  assign n63943 = ~n61802 & n63807;
  assign n63944 = ~n61821 & n63809;
  assign n63945 = n63821 & ~n63941;
  assign n63946 = P2_P3_REIP_REG_6_ & n63823;
  assign n63947 = P2_P3_PHYADDRPOINTER_REG_6_ & n63805;
  assign n63948 = ~n61859 & n63818;
  assign n63949 = ~n63945 & ~n63946;
  assign n63950 = ~n63947 & n63949;
  assign n63951 = ~n63948 & n63950;
  assign n63952 = ~n63937 & ~n63942;
  assign n63953 = ~n63943 & n63952;
  assign n63954 = ~n63944 & n63953;
  assign n11231 = ~n63951 | ~n63954;
  assign n63956 = P2_P3_PHYADDRPOINTER_REG_6_ & n63933;
  assign n63957 = ~P2_P3_PHYADDRPOINTER_REG_7_ & n63956;
  assign n63958 = P2_P3_PHYADDRPOINTER_REG_7_ & ~n63956;
  assign n63959 = ~n63957 & ~n63958;
  assign n63960 = n63812 & ~n63959;
  assign n63961 = P2_P3_PHYADDRPOINTER_REG_6_ & n63938;
  assign n63962 = ~P2_P3_PHYADDRPOINTER_REG_7_ & n63961;
  assign n63963 = P2_P3_PHYADDRPOINTER_REG_7_ & ~n63961;
  assign n63964 = ~n63962 & ~n63963;
  assign n63965 = n63814 & ~n63964;
  assign n63966 = ~n61903 & n63807;
  assign n63967 = ~n61921 & n63809;
  assign n63968 = n63821 & ~n63964;
  assign n63969 = P2_P3_REIP_REG_7_ & n63823;
  assign n63970 = P2_P3_PHYADDRPOINTER_REG_7_ & n63805;
  assign n63971 = ~n61957 & n63818;
  assign n63972 = ~n63968 & ~n63969;
  assign n63973 = ~n63970 & n63972;
  assign n63974 = ~n63971 & n63973;
  assign n63975 = ~n63960 & ~n63965;
  assign n63976 = ~n63966 & n63975;
  assign n63977 = ~n63967 & n63976;
  assign n11236 = ~n63974 | ~n63977;
  assign n63979 = P2_P3_PHYADDRPOINTER_REG_7_ & n63956;
  assign n63980 = ~P2_P3_PHYADDRPOINTER_REG_8_ & n63979;
  assign n63981 = P2_P3_PHYADDRPOINTER_REG_8_ & ~n63979;
  assign n63982 = ~n63980 & ~n63981;
  assign n63983 = n63812 & ~n63982;
  assign n63984 = P2_P3_PHYADDRPOINTER_REG_7_ & n63961;
  assign n63985 = ~P2_P3_PHYADDRPOINTER_REG_8_ & n63984;
  assign n63986 = P2_P3_PHYADDRPOINTER_REG_8_ & ~n63984;
  assign n63987 = ~n63985 & ~n63986;
  assign n63988 = n63814 & ~n63987;
  assign n63989 = ~n61997 & n63807;
  assign n63990 = ~n62013 & n63809;
  assign n63991 = n63821 & ~n63987;
  assign n63992 = P2_P3_REIP_REG_8_ & n63823;
  assign n63993 = P2_P3_PHYADDRPOINTER_REG_8_ & n63805;
  assign n63994 = ~n62047 & n63818;
  assign n63995 = ~n63991 & ~n63992;
  assign n63996 = ~n63993 & n63995;
  assign n63997 = ~n63994 & n63996;
  assign n63998 = ~n63983 & ~n63988;
  assign n63999 = ~n63989 & n63998;
  assign n64000 = ~n63990 & n63999;
  assign n11241 = ~n63997 | ~n64000;
  assign n64002 = P2_P3_PHYADDRPOINTER_REG_8_ & n63979;
  assign n64003 = ~P2_P3_PHYADDRPOINTER_REG_9_ & n64002;
  assign n64004 = P2_P3_PHYADDRPOINTER_REG_9_ & ~n64002;
  assign n64005 = ~n64003 & ~n64004;
  assign n64006 = n63812 & ~n64005;
  assign n64007 = P2_P3_PHYADDRPOINTER_REG_8_ & n63984;
  assign n64008 = ~P2_P3_PHYADDRPOINTER_REG_9_ & n64007;
  assign n64009 = P2_P3_PHYADDRPOINTER_REG_9_ & ~n64007;
  assign n64010 = ~n64008 & ~n64009;
  assign n64011 = n63814 & ~n64010;
  assign n64012 = ~n62090 & n63807;
  assign n64013 = n62101 & n63809;
  assign n64014 = n63821 & ~n64010;
  assign n64015 = P2_P3_REIP_REG_9_ & n63823;
  assign n64016 = P2_P3_PHYADDRPOINTER_REG_9_ & n63805;
  assign n64017 = n62130 & n63818;
  assign n64018 = ~n64014 & ~n64015;
  assign n64019 = ~n64016 & n64018;
  assign n64020 = ~n64017 & n64019;
  assign n64021 = ~n64006 & ~n64011;
  assign n64022 = ~n64012 & n64021;
  assign n64023 = ~n64013 & n64022;
  assign n11246 = ~n64020 | ~n64023;
  assign n64025 = P2_P3_PHYADDRPOINTER_REG_9_ & n64002;
  assign n64026 = ~P2_P3_PHYADDRPOINTER_REG_10_ & n64025;
  assign n64027 = P2_P3_PHYADDRPOINTER_REG_10_ & ~n64025;
  assign n64028 = ~n64026 & ~n64027;
  assign n64029 = n63812 & ~n64028;
  assign n64030 = P2_P3_PHYADDRPOINTER_REG_9_ & n64007;
  assign n64031 = ~P2_P3_PHYADDRPOINTER_REG_10_ & n64030;
  assign n64032 = P2_P3_PHYADDRPOINTER_REG_10_ & ~n64030;
  assign n64033 = ~n64031 & ~n64032;
  assign n64034 = n63814 & ~n64033;
  assign n64035 = ~n62173 & n63807;
  assign n64036 = n62181 & n63809;
  assign n64037 = n63821 & ~n64033;
  assign n64038 = P2_P3_REIP_REG_10_ & n63823;
  assign n64039 = P2_P3_PHYADDRPOINTER_REG_10_ & n63805;
  assign n64040 = n62206 & n63818;
  assign n64041 = ~n64037 & ~n64038;
  assign n64042 = ~n64039 & n64041;
  assign n64043 = ~n64040 & n64042;
  assign n64044 = ~n64029 & ~n64034;
  assign n64045 = ~n64035 & n64044;
  assign n64046 = ~n64036 & n64045;
  assign n11251 = ~n64043 | ~n64046;
  assign n64048 = P2_P3_PHYADDRPOINTER_REG_10_ & n64025;
  assign n64049 = ~P2_P3_PHYADDRPOINTER_REG_11_ & n64048;
  assign n64050 = P2_P3_PHYADDRPOINTER_REG_11_ & ~n64048;
  assign n64051 = ~n64049 & ~n64050;
  assign n64052 = n63812 & ~n64051;
  assign n64053 = P2_P3_PHYADDRPOINTER_REG_10_ & n64030;
  assign n64054 = ~P2_P3_PHYADDRPOINTER_REG_11_ & n64053;
  assign n64055 = P2_P3_PHYADDRPOINTER_REG_11_ & ~n64053;
  assign n64056 = ~n64054 & ~n64055;
  assign n64057 = n63814 & ~n64056;
  assign n64058 = ~n62267 & n63807;
  assign n64059 = ~n62280 & n63809;
  assign n64060 = n63821 & ~n64056;
  assign n64061 = P2_P3_REIP_REG_11_ & n63823;
  assign n64062 = P2_P3_PHYADDRPOINTER_REG_11_ & n63805;
  assign n64063 = ~n62250 & n63818;
  assign n64064 = ~n64060 & ~n64061;
  assign n64065 = ~n64062 & n64064;
  assign n64066 = ~n64063 & n64065;
  assign n64067 = ~n64052 & ~n64057;
  assign n64068 = ~n64058 & n64067;
  assign n64069 = ~n64059 & n64068;
  assign n11256 = ~n64066 | ~n64069;
  assign n64071 = P2_P3_PHYADDRPOINTER_REG_11_ & n64048;
  assign n64072 = ~P2_P3_PHYADDRPOINTER_REG_12_ & n64071;
  assign n64073 = P2_P3_PHYADDRPOINTER_REG_12_ & ~n64071;
  assign n64074 = ~n64072 & ~n64073;
  assign n64075 = n63812 & ~n64074;
  assign n64076 = P2_P3_PHYADDRPOINTER_REG_11_ & n64053;
  assign n64077 = ~P2_P3_PHYADDRPOINTER_REG_12_ & n64076;
  assign n64078 = P2_P3_PHYADDRPOINTER_REG_12_ & ~n64076;
  assign n64079 = ~n64077 & ~n64078;
  assign n64080 = n63814 & ~n64079;
  assign n64081 = ~n62321 & n63807;
  assign n64082 = n62330 & n63809;
  assign n64083 = P2_P3_PHYADDRPOINTER_REG_12_ & n63805;
  assign n64084 = P2_P3_REIP_REG_12_ & n63823;
  assign n64085 = n63821 & ~n64079;
  assign n64086 = n62356 & n63818;
  assign n64087 = ~n64083 & ~n64084;
  assign n64088 = ~n64085 & n64087;
  assign n64089 = ~n64086 & n64088;
  assign n64090 = ~n64075 & ~n64080;
  assign n64091 = ~n64081 & n64090;
  assign n64092 = ~n64082 & n64091;
  assign n11261 = ~n64089 | ~n64092;
  assign n64094 = P2_P3_PHYADDRPOINTER_REG_12_ & n64071;
  assign n64095 = ~P2_P3_PHYADDRPOINTER_REG_13_ & n64094;
  assign n64096 = P2_P3_PHYADDRPOINTER_REG_13_ & ~n64094;
  assign n64097 = ~n64095 & ~n64096;
  assign n64098 = n63812 & ~n64097;
  assign n64099 = P2_P3_PHYADDRPOINTER_REG_12_ & n64076;
  assign n64100 = ~P2_P3_PHYADDRPOINTER_REG_13_ & n64099;
  assign n64101 = P2_P3_PHYADDRPOINTER_REG_13_ & ~n64099;
  assign n64102 = ~n64100 & ~n64101;
  assign n64103 = n63814 & ~n64102;
  assign n64104 = n62399 & n63807;
  assign n64105 = n62406 & n63809;
  assign n64106 = P2_P3_PHYADDRPOINTER_REG_13_ & n63805;
  assign n64107 = P2_P3_REIP_REG_13_ & n63823;
  assign n64108 = n63821 & ~n64102;
  assign n64109 = n62431 & n63818;
  assign n64110 = ~n64106 & ~n64107;
  assign n64111 = ~n64108 & n64110;
  assign n64112 = ~n64109 & n64111;
  assign n64113 = ~n64098 & ~n64103;
  assign n64114 = ~n64104 & n64113;
  assign n64115 = ~n64105 & n64114;
  assign n11266 = ~n64112 | ~n64115;
  assign n64117 = P2_P3_PHYADDRPOINTER_REG_13_ & n64094;
  assign n64118 = ~P2_P3_PHYADDRPOINTER_REG_14_ & n64117;
  assign n64119 = P2_P3_PHYADDRPOINTER_REG_14_ & ~n64117;
  assign n64120 = ~n64118 & ~n64119;
  assign n64121 = n63812 & ~n64120;
  assign n64122 = P2_P3_PHYADDRPOINTER_REG_13_ & n64099;
  assign n64123 = ~P2_P3_PHYADDRPOINTER_REG_14_ & n64122;
  assign n64124 = P2_P3_PHYADDRPOINTER_REG_14_ & ~n64122;
  assign n64125 = ~n64123 & ~n64124;
  assign n64126 = n63814 & ~n64125;
  assign n64127 = ~n62502 & n63807;
  assign n64128 = ~n62506 & n63809;
  assign n64129 = P2_P3_PHYADDRPOINTER_REG_14_ & n63805;
  assign n64130 = P2_P3_REIP_REG_14_ & n63823;
  assign n64131 = n63821 & ~n64125;
  assign n64132 = ~n62475 & n63818;
  assign n64133 = ~n64129 & ~n64130;
  assign n64134 = ~n64131 & n64133;
  assign n64135 = ~n64132 & n64134;
  assign n64136 = ~n64121 & ~n64126;
  assign n64137 = ~n64127 & n64136;
  assign n64138 = ~n64128 & n64137;
  assign n11271 = ~n64135 | ~n64138;
  assign n64140 = P2_P3_PHYADDRPOINTER_REG_14_ & n64117;
  assign n64141 = ~P2_P3_PHYADDRPOINTER_REG_15_ & n64140;
  assign n64142 = P2_P3_PHYADDRPOINTER_REG_15_ & ~n64140;
  assign n64143 = ~n64141 & ~n64142;
  assign n64144 = n63812 & ~n64143;
  assign n64145 = P2_P3_PHYADDRPOINTER_REG_14_ & n64122;
  assign n64146 = ~P2_P3_PHYADDRPOINTER_REG_15_ & n64145;
  assign n64147 = P2_P3_PHYADDRPOINTER_REG_15_ & ~n64145;
  assign n64148 = ~n64146 & ~n64147;
  assign n64149 = n63814 & ~n64148;
  assign n64150 = ~n62579 & n63807;
  assign n64151 = n62584 & n63809;
  assign n64152 = P2_P3_PHYADDRPOINTER_REG_15_ & n63805;
  assign n64153 = P2_P3_REIP_REG_15_ & n63823;
  assign n64154 = n63821 & ~n64148;
  assign n64155 = n62551 & n63818;
  assign n64156 = ~n64152 & ~n64153;
  assign n64157 = ~n64154 & n64156;
  assign n64158 = ~n64155 & n64157;
  assign n64159 = ~n64144 & ~n64149;
  assign n64160 = ~n64150 & n64159;
  assign n64161 = ~n64151 & n64160;
  assign n11276 = ~n64158 | ~n64161;
  assign n64163 = P2_P3_PHYADDRPOINTER_REG_15_ & n64140;
  assign n64164 = ~P2_P3_PHYADDRPOINTER_REG_16_ & n64163;
  assign n64165 = P2_P3_PHYADDRPOINTER_REG_16_ & ~n64163;
  assign n64166 = ~n64164 & ~n64165;
  assign n64167 = n63812 & ~n64166;
  assign n64168 = P2_P3_PHYADDRPOINTER_REG_15_ & n64145;
  assign n64169 = ~P2_P3_PHYADDRPOINTER_REG_16_ & n64168;
  assign n64170 = P2_P3_PHYADDRPOINTER_REG_16_ & ~n64168;
  assign n64171 = ~n64169 & ~n64170;
  assign n64172 = n63814 & ~n64171;
  assign n64173 = ~n62643 & n63807;
  assign n64174 = ~n62656 & n63809;
  assign n64175 = P2_P3_PHYADDRPOINTER_REG_16_ & n63805;
  assign n64176 = P2_P3_REIP_REG_16_ & n63823;
  assign n64177 = n63821 & ~n64171;
  assign n64178 = ~n62626 & n63818;
  assign n64179 = ~n64175 & ~n64176;
  assign n64180 = ~n64177 & n64179;
  assign n64181 = ~n64178 & n64180;
  assign n64182 = ~n64167 & ~n64172;
  assign n64183 = ~n64173 & n64182;
  assign n64184 = ~n64174 & n64183;
  assign n11281 = ~n64181 | ~n64184;
  assign n64186 = P2_P3_PHYADDRPOINTER_REG_16_ & n64163;
  assign n64187 = ~P2_P3_PHYADDRPOINTER_REG_17_ & n64186;
  assign n64188 = P2_P3_PHYADDRPOINTER_REG_17_ & ~n64186;
  assign n64189 = ~n64187 & ~n64188;
  assign n64190 = n63812 & ~n64189;
  assign n64191 = P2_P3_PHYADDRPOINTER_REG_16_ & n64168;
  assign n64192 = ~P2_P3_PHYADDRPOINTER_REG_17_ & n64191;
  assign n64193 = P2_P3_PHYADDRPOINTER_REG_17_ & ~n64191;
  assign n64194 = ~n64192 & ~n64193;
  assign n64195 = n63814 & ~n64194;
  assign n64196 = n62699 & n63807;
  assign n64197 = n62707 & n63809;
  assign n64198 = P2_P3_PHYADDRPOINTER_REG_17_ & n63805;
  assign n64199 = P2_P3_REIP_REG_17_ & n63823;
  assign n64200 = n63821 & ~n64194;
  assign n64201 = n62733 & n63818;
  assign n64202 = ~n64198 & ~n64199;
  assign n64203 = ~n64200 & n64202;
  assign n64204 = ~n64201 & n64203;
  assign n64205 = ~n64190 & ~n64195;
  assign n64206 = ~n64196 & n64205;
  assign n64207 = ~n64197 & n64206;
  assign n11286 = ~n64204 | ~n64207;
  assign n64209 = P2_P3_PHYADDRPOINTER_REG_17_ & n64186;
  assign n64210 = ~P2_P3_PHYADDRPOINTER_REG_18_ & n64209;
  assign n64211 = P2_P3_PHYADDRPOINTER_REG_18_ & ~n64209;
  assign n64212 = ~n64210 & ~n64211;
  assign n64213 = n63812 & ~n64212;
  assign n64214 = P2_P3_PHYADDRPOINTER_REG_17_ & n64191;
  assign n64215 = ~P2_P3_PHYADDRPOINTER_REG_18_ & n64214;
  assign n64216 = P2_P3_PHYADDRPOINTER_REG_18_ & ~n64214;
  assign n64217 = ~n64215 & ~n64216;
  assign n64218 = n63814 & ~n64217;
  assign n64219 = ~n62793 & n63807;
  assign n64220 = ~n62806 & n63809;
  assign n64221 = P2_P3_PHYADDRPOINTER_REG_18_ & n63805;
  assign n64222 = P2_P3_REIP_REG_18_ & n63823;
  assign n64223 = n63821 & ~n64217;
  assign n64224 = ~n62777 & n63818;
  assign n64225 = ~n64221 & ~n64222;
  assign n64226 = ~n64223 & n64225;
  assign n64227 = ~n64224 & n64226;
  assign n64228 = ~n64213 & ~n64218;
  assign n64229 = ~n64219 & n64228;
  assign n64230 = ~n64220 & n64229;
  assign n11291 = ~n64227 | ~n64230;
  assign n64232 = P2_P3_PHYADDRPOINTER_REG_18_ & n64209;
  assign n64233 = ~P2_P3_PHYADDRPOINTER_REG_19_ & n64232;
  assign n64234 = P2_P3_PHYADDRPOINTER_REG_19_ & ~n64232;
  assign n64235 = ~n64233 & ~n64234;
  assign n64236 = n63812 & ~n64235;
  assign n64237 = P2_P3_PHYADDRPOINTER_REG_18_ & n64214;
  assign n64238 = ~P2_P3_PHYADDRPOINTER_REG_19_ & n64237;
  assign n64239 = P2_P3_PHYADDRPOINTER_REG_19_ & ~n64237;
  assign n64240 = ~n64238 & ~n64239;
  assign n64241 = n63814 & ~n64240;
  assign n64242 = ~n62847 & n63807;
  assign n64243 = n62856 & n63809;
  assign n64244 = P2_P3_PHYADDRPOINTER_REG_19_ & n63805;
  assign n64245 = P2_P3_REIP_REG_19_ & n63823;
  assign n64246 = n63821 & ~n64240;
  assign n64247 = n62882 & n63818;
  assign n64248 = ~n64244 & ~n64245;
  assign n64249 = ~n64246 & n64248;
  assign n64250 = ~n64247 & n64249;
  assign n64251 = ~n64236 & ~n64241;
  assign n64252 = ~n64242 & n64251;
  assign n64253 = ~n64243 & n64252;
  assign n11296 = ~n64250 | ~n64253;
  assign n64255 = P2_P3_PHYADDRPOINTER_REG_19_ & n64232;
  assign n64256 = ~P2_P3_PHYADDRPOINTER_REG_20_ & n64255;
  assign n64257 = P2_P3_PHYADDRPOINTER_REG_20_ & ~n64255;
  assign n64258 = ~n64256 & ~n64257;
  assign n64259 = n63812 & ~n64258;
  assign n64260 = P2_P3_PHYADDRPOINTER_REG_19_ & n64237;
  assign n64261 = ~P2_P3_PHYADDRPOINTER_REG_20_ & n64260;
  assign n64262 = P2_P3_PHYADDRPOINTER_REG_20_ & ~n64260;
  assign n64263 = ~n64261 & ~n64262;
  assign n64264 = n63814 & ~n64263;
  assign n64265 = n62934 & n63809;
  assign n64266 = P2_P3_PHYADDRPOINTER_REG_20_ & n63805;
  assign n64267 = P2_P3_REIP_REG_20_ & n63823;
  assign n64268 = n63821 & ~n64263;
  assign n64269 = n62958 & n63818;
  assign n64270 = ~n64266 & ~n64267;
  assign n64271 = ~n64268 & n64270;
  assign n64272 = ~n64269 & n64271;
  assign n64273 = n62909 & n63807;
  assign n64274 = ~n64259 & ~n64264;
  assign n64275 = ~n64265 & n64274;
  assign n64276 = n64272 & n64275;
  assign n11301 = n64273 | ~n64276;
  assign n64278 = P2_P3_PHYADDRPOINTER_REG_20_ & n64255;
  assign n64279 = ~P2_P3_PHYADDRPOINTER_REG_21_ & n64278;
  assign n64280 = P2_P3_PHYADDRPOINTER_REG_21_ & ~n64278;
  assign n64281 = ~n64279 & ~n64280;
  assign n64282 = n63812 & ~n64281;
  assign n64283 = P2_P3_PHYADDRPOINTER_REG_20_ & n64260;
  assign n64284 = ~P2_P3_PHYADDRPOINTER_REG_21_ & n64283;
  assign n64285 = P2_P3_PHYADDRPOINTER_REG_21_ & ~n64283;
  assign n64286 = ~n64284 & ~n64285;
  assign n64287 = n63814 & ~n64286;
  assign n64288 = n62991 & n63809;
  assign n64289 = P2_P3_PHYADDRPOINTER_REG_21_ & n63805;
  assign n64290 = P2_P3_REIP_REG_21_ & n63823;
  assign n64291 = n63821 & ~n64286;
  assign n64292 = n63016 & n63818;
  assign n64293 = ~n64289 & ~n64290;
  assign n64294 = ~n64291 & n64293;
  assign n64295 = ~n64292 & n64294;
  assign n64296 = ~n63032 & n63807;
  assign n64297 = ~n64282 & ~n64287;
  assign n64298 = ~n64288 & n64297;
  assign n64299 = n64295 & n64298;
  assign n11306 = n64296 | ~n64299;
  assign n64301 = P2_P3_PHYADDRPOINTER_REG_21_ & n64278;
  assign n64302 = ~P2_P3_PHYADDRPOINTER_REG_22_ & n64301;
  assign n64303 = P2_P3_PHYADDRPOINTER_REG_22_ & ~n64301;
  assign n64304 = ~n64302 & ~n64303;
  assign n64305 = n63812 & ~n64304;
  assign n64306 = ~n63093 & n63807;
  assign n64307 = P2_P3_PHYADDRPOINTER_REG_21_ & n64283;
  assign n64308 = ~P2_P3_PHYADDRPOINTER_REG_22_ & n64307;
  assign n64309 = P2_P3_PHYADDRPOINTER_REG_22_ & ~n64307;
  assign n64310 = ~n64308 & ~n64309;
  assign n64311 = n63814 & ~n64310;
  assign n64312 = ~n63110 & n63809;
  assign n64313 = P2_P3_PHYADDRPOINTER_REG_22_ & n63805;
  assign n64314 = P2_P3_REIP_REG_22_ & n63823;
  assign n64315 = n63821 & ~n64310;
  assign n64316 = ~n63072 & n63818;
  assign n64317 = ~n64313 & ~n64314;
  assign n64318 = ~n64315 & n64317;
  assign n64319 = ~n64316 & n64318;
  assign n64320 = ~n64305 & ~n64306;
  assign n64321 = ~n64311 & n64320;
  assign n64322 = ~n64312 & n64321;
  assign n11311 = ~n64319 | ~n64322;
  assign n64324 = P2_P3_PHYADDRPOINTER_REG_22_ & n64301;
  assign n64325 = ~P2_P3_PHYADDRPOINTER_REG_23_ & n64324;
  assign n64326 = P2_P3_PHYADDRPOINTER_REG_23_ & ~n64324;
  assign n64327 = ~n64325 & ~n64326;
  assign n64328 = n63812 & ~n64327;
  assign n64329 = ~n63169 & n63807;
  assign n64330 = P2_P3_PHYADDRPOINTER_REG_22_ & n64307;
  assign n64331 = ~P2_P3_PHYADDRPOINTER_REG_23_ & n64330;
  assign n64332 = P2_P3_PHYADDRPOINTER_REG_23_ & ~n64330;
  assign n64333 = ~n64331 & ~n64332;
  assign n64334 = n63814 & ~n64333;
  assign n64335 = n63187 & n63809;
  assign n64336 = P2_P3_PHYADDRPOINTER_REG_23_ & n63805;
  assign n64337 = P2_P3_REIP_REG_23_ & n63823;
  assign n64338 = n63821 & ~n64333;
  assign n64339 = n63151 & n63818;
  assign n64340 = ~n64336 & ~n64337;
  assign n64341 = ~n64338 & n64340;
  assign n64342 = ~n64339 & n64341;
  assign n64343 = ~n64328 & ~n64329;
  assign n64344 = ~n64334 & n64343;
  assign n64345 = ~n64335 & n64344;
  assign n11316 = ~n64342 | ~n64345;
  assign n64347 = P2_P3_PHYADDRPOINTER_REG_23_ & n64324;
  assign n64348 = ~P2_P3_PHYADDRPOINTER_REG_24_ & n64347;
  assign n64349 = P2_P3_PHYADDRPOINTER_REG_24_ & ~n64347;
  assign n64350 = ~n64348 & ~n64349;
  assign n64351 = n63812 & ~n64350;
  assign n64352 = ~n63244 & n63807;
  assign n64353 = P2_P3_PHYADDRPOINTER_REG_23_ & n64330;
  assign n64354 = ~P2_P3_PHYADDRPOINTER_REG_24_ & n64353;
  assign n64355 = P2_P3_PHYADDRPOINTER_REG_24_ & ~n64353;
  assign n64356 = ~n64354 & ~n64355;
  assign n64357 = n63814 & ~n64356;
  assign n64358 = ~n63252 & n63809;
  assign n64359 = P2_P3_PHYADDRPOINTER_REG_24_ & n63805;
  assign n64360 = P2_P3_REIP_REG_24_ & n63823;
  assign n64361 = n63821 & ~n64356;
  assign n64362 = ~n63217 & n63818;
  assign n64363 = ~n64359 & ~n64360;
  assign n64364 = ~n64361 & n64363;
  assign n64365 = ~n64362 & n64364;
  assign n64366 = ~n64351 & ~n64352;
  assign n64367 = ~n64357 & n64366;
  assign n64368 = ~n64358 & n64367;
  assign n11321 = ~n64365 | ~n64368;
  assign n64370 = P2_P3_PHYADDRPOINTER_REG_24_ & n64347;
  assign n64371 = ~P2_P3_PHYADDRPOINTER_REG_25_ & n64370;
  assign n64372 = P2_P3_PHYADDRPOINTER_REG_25_ & ~n64370;
  assign n64373 = ~n64371 & ~n64372;
  assign n64374 = n63812 & ~n64373;
  assign n64375 = ~n63321 & n63807;
  assign n64376 = P2_P3_PHYADDRPOINTER_REG_24_ & n64353;
  assign n64377 = ~P2_P3_PHYADDRPOINTER_REG_25_ & n64376;
  assign n64378 = P2_P3_PHYADDRPOINTER_REG_25_ & ~n64376;
  assign n64379 = ~n64377 & ~n64378;
  assign n64380 = n63814 & ~n64379;
  assign n64381 = n63327 & n63809;
  assign n64382 = P2_P3_PHYADDRPOINTER_REG_25_ & n63805;
  assign n64383 = P2_P3_REIP_REG_25_ & n63823;
  assign n64384 = n63821 & ~n64379;
  assign n64385 = n63293 & n63818;
  assign n64386 = ~n64382 & ~n64383;
  assign n64387 = ~n64384 & n64386;
  assign n64388 = ~n64385 & n64387;
  assign n64389 = ~n64374 & ~n64375;
  assign n64390 = ~n64380 & n64389;
  assign n64391 = ~n64381 & n64390;
  assign n11326 = ~n64388 | ~n64391;
  assign n64393 = P2_P3_PHYADDRPOINTER_REG_25_ & n64370;
  assign n64394 = ~P2_P3_PHYADDRPOINTER_REG_26_ & n64393;
  assign n64395 = P2_P3_PHYADDRPOINTER_REG_26_ & ~n64393;
  assign n64396 = ~n64394 & ~n64395;
  assign n64397 = n63812 & ~n64396;
  assign n64398 = n63362 & n63807;
  assign n64399 = P2_P3_PHYADDRPOINTER_REG_25_ & n64376;
  assign n64400 = ~P2_P3_PHYADDRPOINTER_REG_26_ & n64399;
  assign n64401 = P2_P3_PHYADDRPOINTER_REG_26_ & ~n64399;
  assign n64402 = ~n64400 & ~n64401;
  assign n64403 = n63814 & ~n64402;
  assign n64404 = n63366 & n63809;
  assign n64405 = P2_P3_PHYADDRPOINTER_REG_26_ & n63805;
  assign n64406 = n63404 & n63818;
  assign n64407 = n63821 & ~n64402;
  assign n64408 = P2_P3_REIP_REG_26_ & n63823;
  assign n64409 = ~n64405 & ~n64406;
  assign n64410 = ~n64407 & n64409;
  assign n64411 = ~n64408 & n64410;
  assign n64412 = ~n64397 & ~n64398;
  assign n64413 = ~n64403 & n64412;
  assign n64414 = ~n64404 & n64413;
  assign n11331 = ~n64411 | ~n64414;
  assign n64416 = P2_P3_PHYADDRPOINTER_REG_26_ & n64393;
  assign n64417 = ~P2_P3_PHYADDRPOINTER_REG_27_ & n64416;
  assign n64418 = P2_P3_PHYADDRPOINTER_REG_27_ & ~n64416;
  assign n64419 = ~n64417 & ~n64418;
  assign n64420 = n63812 & ~n64419;
  assign n64421 = ~n63433 & n63807;
  assign n64422 = P2_P3_PHYADDRPOINTER_REG_26_ & n64399;
  assign n64423 = ~P2_P3_PHYADDRPOINTER_REG_27_ & n64422;
  assign n64424 = P2_P3_PHYADDRPOINTER_REG_27_ & ~n64422;
  assign n64425 = ~n64423 & ~n64424;
  assign n64426 = n63814 & ~n64425;
  assign n64427 = ~n63437 & n63809;
  assign n64428 = P2_P3_PHYADDRPOINTER_REG_27_ & n63805;
  assign n64429 = ~n63475 & n63818;
  assign n64430 = n63821 & ~n64425;
  assign n64431 = P2_P3_REIP_REG_27_ & n63823;
  assign n64432 = ~n64428 & ~n64429;
  assign n64433 = ~n64430 & n64432;
  assign n64434 = ~n64431 & n64433;
  assign n64435 = ~n64420 & ~n64421;
  assign n64436 = ~n64426 & n64435;
  assign n64437 = ~n64427 & n64436;
  assign n11336 = ~n64434 | ~n64437;
  assign n64439 = n63511 & n63807;
  assign n64440 = n63516 & n63809;
  assign n64441 = P2_P3_PHYADDRPOINTER_REG_27_ & n64416;
  assign n64442 = ~P2_P3_PHYADDRPOINTER_REG_28_ & n64441;
  assign n64443 = P2_P3_PHYADDRPOINTER_REG_28_ & ~n64441;
  assign n64444 = ~n64442 & ~n64443;
  assign n64445 = n63812 & ~n64444;
  assign n64446 = P2_P3_PHYADDRPOINTER_REG_27_ & n64422;
  assign n64447 = ~P2_P3_PHYADDRPOINTER_REG_28_ & n64446;
  assign n64448 = P2_P3_PHYADDRPOINTER_REG_28_ & ~n64446;
  assign n64449 = ~n64447 & ~n64448;
  assign n64450 = n63814 & ~n64449;
  assign n64451 = P2_P3_PHYADDRPOINTER_REG_28_ & n63805;
  assign n64452 = n63555 & n63818;
  assign n64453 = n63821 & ~n64449;
  assign n64454 = P2_P3_REIP_REG_28_ & n63823;
  assign n64455 = ~n64451 & ~n64452;
  assign n64456 = ~n64453 & n64455;
  assign n64457 = ~n64454 & n64456;
  assign n64458 = ~n64439 & ~n64440;
  assign n64459 = ~n64445 & n64458;
  assign n64460 = ~n64450 & n64459;
  assign n11341 = ~n64457 | ~n64460;
  assign n64462 = ~n63584 & n63807;
  assign n64463 = n63588 & n63809;
  assign n64464 = P2_P3_PHYADDRPOINTER_REG_28_ & n64441;
  assign n64465 = ~P2_P3_PHYADDRPOINTER_REG_29_ & n64464;
  assign n64466 = P2_P3_PHYADDRPOINTER_REG_29_ & ~n64464;
  assign n64467 = ~n64465 & ~n64466;
  assign n64468 = n63812 & ~n64467;
  assign n64469 = P2_P3_PHYADDRPOINTER_REG_28_ & n64446;
  assign n64470 = ~P2_P3_PHYADDRPOINTER_REG_29_ & n64469;
  assign n64471 = P2_P3_PHYADDRPOINTER_REG_29_ & ~n64469;
  assign n64472 = ~n64470 & ~n64471;
  assign n64473 = n63814 & ~n64472;
  assign n64474 = P2_P3_PHYADDRPOINTER_REG_29_ & n63805;
  assign n64475 = P2_P3_REIP_REG_29_ & n63823;
  assign n64476 = n63626 & n63818;
  assign n64477 = n63821 & ~n64472;
  assign n64478 = ~n64474 & ~n64475;
  assign n64479 = ~n64476 & n64478;
  assign n64480 = ~n64477 & n64479;
  assign n64481 = ~n64462 & ~n64463;
  assign n64482 = ~n64468 & n64481;
  assign n64483 = ~n64473 & n64482;
  assign n11346 = ~n64480 | ~n64483;
  assign n64485 = ~n63656 & n63807;
  assign n64486 = ~n63660 & n63809;
  assign n64487 = P2_P3_PHYADDRPOINTER_REG_29_ & n64464;
  assign n64488 = ~P2_P3_PHYADDRPOINTER_REG_30_ & n64487;
  assign n64489 = P2_P3_PHYADDRPOINTER_REG_30_ & ~n64487;
  assign n64490 = ~n64488 & ~n64489;
  assign n64491 = n63812 & ~n64490;
  assign n64492 = P2_P3_PHYADDRPOINTER_REG_29_ & n64469;
  assign n64493 = ~P2_P3_PHYADDRPOINTER_REG_30_ & n64492;
  assign n64494 = P2_P3_PHYADDRPOINTER_REG_30_ & ~n64492;
  assign n64495 = ~n64493 & ~n64494;
  assign n64496 = n63814 & ~n64495;
  assign n64497 = P2_P3_PHYADDRPOINTER_REG_30_ & n63805;
  assign n64498 = P2_P3_REIP_REG_30_ & n63823;
  assign n64499 = ~n63698 & n63818;
  assign n64500 = n63821 & ~n64495;
  assign n64501 = ~n64497 & ~n64498;
  assign n64502 = ~n64499 & n64501;
  assign n64503 = ~n64500 & n64502;
  assign n64504 = ~n64485 & ~n64486;
  assign n64505 = ~n64491 & n64504;
  assign n64506 = ~n64496 & n64505;
  assign n11351 = ~n64503 | ~n64506;
  assign n64508 = n63769 & n63807;
  assign n64509 = P2_P3_PHYADDRPOINTER_REG_30_ & n64487;
  assign n64510 = ~P2_P3_PHYADDRPOINTER_REG_31_ & n64509;
  assign n64511 = P2_P3_PHYADDRPOINTER_REG_31_ & ~n64509;
  assign n64512 = ~n64510 & ~n64511;
  assign n64513 = n63812 & ~n64512;
  assign n64514 = ~n63774 & n63809;
  assign n64515 = P2_P3_PHYADDRPOINTER_REG_30_ & n64492;
  assign n64516 = ~P2_P3_PHYADDRPOINTER_REG_31_ & n64515;
  assign n64517 = P2_P3_PHYADDRPOINTER_REG_31_ & ~n64515;
  assign n64518 = ~n64516 & ~n64517;
  assign n64519 = n63814 & ~n64518;
  assign n64520 = P2_P3_PHYADDRPOINTER_REG_31_ & n63805;
  assign n64521 = P2_P3_REIP_REG_31_ & n63823;
  assign n64522 = ~n63722 & n63818;
  assign n64523 = n63821 & ~n64518;
  assign n64524 = ~n64520 & ~n64521;
  assign n64525 = ~n64522 & n64524;
  assign n64526 = ~n64523 & n64525;
  assign n64527 = ~n64508 & ~n64513;
  assign n64528 = ~n64514 & n64527;
  assign n64529 = ~n64519 & n64528;
  assign n11356 = ~n64526 | ~n64529;
  assign n64531 = ~n58594 & n59050;
  assign n64532 = n59019 & n64531;
  assign n64533 = ~n59206 & ~n64532;
  assign n64534 = n59321 & ~n64533;
  assign n64535 = ~n58935 & n64534;
  assign n64536 = P2_BUF2_REG_15_ & n64535;
  assign n64537 = n58935 & n64534;
  assign n64538 = P2_P3_EAX_REG_15_ & n64537;
  assign n64539 = P2_P3_LWORD_REG_15_ & ~n64534;
  assign n64540 = ~n64536 & ~n64538;
  assign n11361 = n64539 | ~n64540;
  assign n64542 = P2_BUF2_REG_14_ & n64535;
  assign n64543 = P2_P3_EAX_REG_14_ & n64537;
  assign n64544 = P2_P3_LWORD_REG_14_ & ~n64534;
  assign n64545 = ~n64542 & ~n64543;
  assign n11366 = n64544 | ~n64545;
  assign n64547 = P2_BUF2_REG_13_ & n64535;
  assign n64548 = P2_P3_EAX_REG_13_ & n64537;
  assign n64549 = P2_P3_LWORD_REG_13_ & ~n64534;
  assign n64550 = ~n64547 & ~n64548;
  assign n11371 = n64549 | ~n64550;
  assign n64552 = P2_BUF2_REG_12_ & n64535;
  assign n64553 = P2_P3_EAX_REG_12_ & n64537;
  assign n64554 = P2_P3_LWORD_REG_12_ & ~n64534;
  assign n64555 = ~n64552 & ~n64553;
  assign n11376 = n64554 | ~n64555;
  assign n64557 = P2_BUF2_REG_11_ & n64535;
  assign n64558 = P2_P3_EAX_REG_11_ & n64537;
  assign n64559 = P2_P3_LWORD_REG_11_ & ~n64534;
  assign n64560 = ~n64557 & ~n64558;
  assign n11381 = n64559 | ~n64560;
  assign n64562 = P2_BUF2_REG_10_ & n64535;
  assign n64563 = P2_P3_EAX_REG_10_ & n64537;
  assign n64564 = P2_P3_LWORD_REG_10_ & ~n64534;
  assign n64565 = ~n64562 & ~n64563;
  assign n11386 = n64564 | ~n64565;
  assign n64567 = P2_BUF2_REG_9_ & n64535;
  assign n64568 = P2_P3_EAX_REG_9_ & n64537;
  assign n64569 = P2_P3_LWORD_REG_9_ & ~n64534;
  assign n64570 = ~n64567 & ~n64568;
  assign n11391 = n64569 | ~n64570;
  assign n64572 = P2_BUF2_REG_8_ & n64535;
  assign n64573 = P2_P3_EAX_REG_8_ & n64537;
  assign n64574 = P2_P3_LWORD_REG_8_ & ~n64534;
  assign n64575 = ~n64572 & ~n64573;
  assign n11396 = n64574 | ~n64575;
  assign n64577 = P2_BUF2_REG_7_ & n64535;
  assign n64578 = P2_P3_EAX_REG_7_ & n64537;
  assign n64579 = P2_P3_LWORD_REG_7_ & ~n64534;
  assign n64580 = ~n64577 & ~n64578;
  assign n11401 = n64579 | ~n64580;
  assign n64582 = P2_BUF2_REG_6_ & n64535;
  assign n64583 = P2_P3_EAX_REG_6_ & n64537;
  assign n64584 = P2_P3_LWORD_REG_6_ & ~n64534;
  assign n64585 = ~n64582 & ~n64583;
  assign n11406 = n64584 | ~n64585;
  assign n64587 = P2_BUF2_REG_5_ & n64535;
  assign n64588 = P2_P3_EAX_REG_5_ & n64537;
  assign n64589 = P2_P3_LWORD_REG_5_ & ~n64534;
  assign n64590 = ~n64587 & ~n64588;
  assign n11411 = n64589 | ~n64590;
  assign n64592 = P2_BUF2_REG_4_ & n64535;
  assign n64593 = P2_P3_EAX_REG_4_ & n64537;
  assign n64594 = P2_P3_LWORD_REG_4_ & ~n64534;
  assign n64595 = ~n64592 & ~n64593;
  assign n11416 = n64594 | ~n64595;
  assign n64597 = P2_BUF2_REG_3_ & n64535;
  assign n64598 = P2_P3_EAX_REG_3_ & n64537;
  assign n64599 = P2_P3_LWORD_REG_3_ & ~n64534;
  assign n64600 = ~n64597 & ~n64598;
  assign n11421 = n64599 | ~n64600;
  assign n64602 = P2_BUF2_REG_2_ & n64535;
  assign n64603 = P2_P3_EAX_REG_2_ & n64537;
  assign n64604 = P2_P3_LWORD_REG_2_ & ~n64534;
  assign n64605 = ~n64602 & ~n64603;
  assign n11426 = n64604 | ~n64605;
  assign n64607 = P2_BUF2_REG_1_ & n64535;
  assign n64608 = P2_P3_EAX_REG_1_ & n64537;
  assign n64609 = P2_P3_LWORD_REG_1_ & ~n64534;
  assign n64610 = ~n64607 & ~n64608;
  assign n11431 = n64609 | ~n64610;
  assign n64612 = P2_BUF2_REG_0_ & n64535;
  assign n64613 = P2_P3_EAX_REG_0_ & n64537;
  assign n64614 = P2_P3_LWORD_REG_0_ & ~n64534;
  assign n64615 = ~n64612 & ~n64613;
  assign n11436 = n64614 | ~n64615;
  assign n64617 = P2_P3_EAX_REG_30_ & n64537;
  assign n64618 = P2_P3_UWORD_REG_14_ & ~n64534;
  assign n64619 = ~n64542 & ~n64617;
  assign n11441 = n64618 | ~n64619;
  assign n64621 = P2_P3_EAX_REG_29_ & n64537;
  assign n64622 = P2_P3_UWORD_REG_13_ & ~n64534;
  assign n64623 = ~n64547 & ~n64621;
  assign n11446 = n64622 | ~n64623;
  assign n64625 = P2_P3_EAX_REG_28_ & n64537;
  assign n64626 = P2_P3_UWORD_REG_12_ & ~n64534;
  assign n64627 = ~n64552 & ~n64625;
  assign n11451 = n64626 | ~n64627;
  assign n64629 = P2_P3_EAX_REG_27_ & n64537;
  assign n64630 = P2_P3_UWORD_REG_11_ & ~n64534;
  assign n64631 = ~n64557 & ~n64629;
  assign n11456 = n64630 | ~n64631;
  assign n64633 = P2_P3_EAX_REG_26_ & n64537;
  assign n64634 = P2_P3_UWORD_REG_10_ & ~n64534;
  assign n64635 = ~n64562 & ~n64633;
  assign n11461 = n64634 | ~n64635;
  assign n64637 = P2_P3_EAX_REG_25_ & n64537;
  assign n64638 = P2_P3_UWORD_REG_9_ & ~n64534;
  assign n64639 = ~n64567 & ~n64637;
  assign n11466 = n64638 | ~n64639;
  assign n64641 = P2_P3_EAX_REG_24_ & n64537;
  assign n64642 = P2_P3_UWORD_REG_8_ & ~n64534;
  assign n64643 = ~n64572 & ~n64641;
  assign n11471 = n64642 | ~n64643;
  assign n64645 = P2_P3_EAX_REG_23_ & n64537;
  assign n64646 = P2_P3_UWORD_REG_7_ & ~n64534;
  assign n64647 = ~n64577 & ~n64645;
  assign n11476 = n64646 | ~n64647;
  assign n64649 = P2_P3_EAX_REG_22_ & n64537;
  assign n64650 = P2_P3_UWORD_REG_6_ & ~n64534;
  assign n64651 = ~n64582 & ~n64649;
  assign n11481 = n64650 | ~n64651;
  assign n64653 = P2_P3_EAX_REG_21_ & n64537;
  assign n64654 = P2_P3_UWORD_REG_5_ & ~n64534;
  assign n64655 = ~n64587 & ~n64653;
  assign n11486 = n64654 | ~n64655;
  assign n64657 = P2_P3_EAX_REG_20_ & n64537;
  assign n64658 = P2_P3_UWORD_REG_4_ & ~n64534;
  assign n64659 = ~n64592 & ~n64657;
  assign n11491 = n64658 | ~n64659;
  assign n64661 = P2_P3_EAX_REG_19_ & n64537;
  assign n64662 = P2_P3_UWORD_REG_3_ & ~n64534;
  assign n64663 = ~n64597 & ~n64661;
  assign n11496 = n64662 | ~n64663;
  assign n64665 = P2_P3_EAX_REG_18_ & n64537;
  assign n64666 = P2_P3_UWORD_REG_2_ & ~n64534;
  assign n64667 = ~n64602 & ~n64665;
  assign n11501 = n64666 | ~n64667;
  assign n64669 = P2_P3_EAX_REG_17_ & n64537;
  assign n64670 = P2_P3_UWORD_REG_1_ & ~n64534;
  assign n64671 = ~n64607 & ~n64669;
  assign n11506 = n64670 | ~n64671;
  assign n64673 = P2_P3_EAX_REG_16_ & n64537;
  assign n64674 = P2_P3_UWORD_REG_0_ & ~n64534;
  assign n64675 = ~n64612 & ~n64673;
  assign n11511 = n64674 | ~n64675;
  assign n64677 = ~P2_P3_STATE2_REG_0_ & n58679;
  assign n64678 = n58685 & n59321;
  assign n64679 = ~n59207 & n64678;
  assign n64680 = ~n64677 & ~n64679;
  assign n64681 = P2_P3_STATE2_REG_0_ & ~n64680;
  assign n64682 = P2_P3_EAX_REG_0_ & n64681;
  assign n64683 = ~P2_P3_STATE2_REG_0_ & ~n64680;
  assign n64684 = P2_P3_LWORD_REG_0_ & n64683;
  assign n64685 = P2_P3_DATAO_REG_0_ & n64680;
  assign n64686 = ~n64682 & ~n64684;
  assign n11516 = n64685 | ~n64686;
  assign n64688 = P2_P3_EAX_REG_1_ & n64681;
  assign n64689 = P2_P3_LWORD_REG_1_ & n64683;
  assign n64690 = P2_P3_DATAO_REG_1_ & n64680;
  assign n64691 = ~n64688 & ~n64689;
  assign n11521 = n64690 | ~n64691;
  assign n64693 = P2_P3_EAX_REG_2_ & n64681;
  assign n64694 = P2_P3_LWORD_REG_2_ & n64683;
  assign n64695 = P2_P3_DATAO_REG_2_ & n64680;
  assign n64696 = ~n64693 & ~n64694;
  assign n11526 = n64695 | ~n64696;
  assign n64698 = P2_P3_EAX_REG_3_ & n64681;
  assign n64699 = P2_P3_LWORD_REG_3_ & n64683;
  assign n64700 = P2_P3_DATAO_REG_3_ & n64680;
  assign n64701 = ~n64698 & ~n64699;
  assign n11531 = n64700 | ~n64701;
  assign n64703 = P2_P3_EAX_REG_4_ & n64681;
  assign n64704 = P2_P3_LWORD_REG_4_ & n64683;
  assign n64705 = P2_P3_DATAO_REG_4_ & n64680;
  assign n64706 = ~n64703 & ~n64704;
  assign n11536 = n64705 | ~n64706;
  assign n64708 = P2_P3_EAX_REG_5_ & n64681;
  assign n64709 = P2_P3_LWORD_REG_5_ & n64683;
  assign n64710 = P2_P3_DATAO_REG_5_ & n64680;
  assign n64711 = ~n64708 & ~n64709;
  assign n11541 = n64710 | ~n64711;
  assign n64713 = P2_P3_EAX_REG_6_ & n64681;
  assign n64714 = P2_P3_LWORD_REG_6_ & n64683;
  assign n64715 = P2_P3_DATAO_REG_6_ & n64680;
  assign n64716 = ~n64713 & ~n64714;
  assign n11546 = n64715 | ~n64716;
  assign n64718 = P2_P3_EAX_REG_7_ & n64681;
  assign n64719 = P2_P3_LWORD_REG_7_ & n64683;
  assign n64720 = P2_P3_DATAO_REG_7_ & n64680;
  assign n64721 = ~n64718 & ~n64719;
  assign n11551 = n64720 | ~n64721;
  assign n64723 = P2_P3_EAX_REG_8_ & n64681;
  assign n64724 = P2_P3_LWORD_REG_8_ & n64683;
  assign n64725 = P2_P3_DATAO_REG_8_ & n64680;
  assign n64726 = ~n64723 & ~n64724;
  assign n11556 = n64725 | ~n64726;
  assign n64728 = P2_P3_EAX_REG_9_ & n64681;
  assign n64729 = P2_P3_LWORD_REG_9_ & n64683;
  assign n64730 = P2_P3_DATAO_REG_9_ & n64680;
  assign n64731 = ~n64728 & ~n64729;
  assign n11561 = n64730 | ~n64731;
  assign n64733 = P2_P3_EAX_REG_10_ & n64681;
  assign n64734 = P2_P3_LWORD_REG_10_ & n64683;
  assign n64735 = P2_P3_DATAO_REG_10_ & n64680;
  assign n64736 = ~n64733 & ~n64734;
  assign n11566 = n64735 | ~n64736;
  assign n64738 = P2_P3_EAX_REG_11_ & n64681;
  assign n64739 = P2_P3_LWORD_REG_11_ & n64683;
  assign n64740 = P2_P3_DATAO_REG_11_ & n64680;
  assign n64741 = ~n64738 & ~n64739;
  assign n11571 = n64740 | ~n64741;
  assign n64743 = P2_P3_EAX_REG_12_ & n64681;
  assign n64744 = P2_P3_LWORD_REG_12_ & n64683;
  assign n64745 = P2_P3_DATAO_REG_12_ & n64680;
  assign n64746 = ~n64743 & ~n64744;
  assign n11576 = n64745 | ~n64746;
  assign n64748 = P2_P3_EAX_REG_13_ & n64681;
  assign n64749 = P2_P3_LWORD_REG_13_ & n64683;
  assign n64750 = P2_P3_DATAO_REG_13_ & n64680;
  assign n64751 = ~n64748 & ~n64749;
  assign n11581 = n64750 | ~n64751;
  assign n64753 = P2_P3_EAX_REG_14_ & n64681;
  assign n64754 = P2_P3_LWORD_REG_14_ & n64683;
  assign n64755 = P2_P3_DATAO_REG_14_ & n64680;
  assign n64756 = ~n64753 & ~n64754;
  assign n11586 = n64755 | ~n64756;
  assign n64758 = P2_P3_EAX_REG_15_ & n64681;
  assign n64759 = P2_P3_LWORD_REG_15_ & n64683;
  assign n64760 = P2_P3_DATAO_REG_15_ & n64680;
  assign n64761 = ~n64758 & ~n64759;
  assign n11591 = n64760 | ~n64761;
  assign n64763 = P2_P3_UWORD_REG_0_ & n64683;
  assign n64764 = P2_P3_DATAO_REG_16_ & n64680;
  assign n64765 = ~n64763 & ~n64764;
  assign n64766 = ~n58966 & n64681;
  assign n64767 = P2_P3_EAX_REG_16_ & n64766;
  assign n11596 = ~n64765 | n64767;
  assign n64769 = P2_P3_UWORD_REG_1_ & n64683;
  assign n64770 = P2_P3_DATAO_REG_17_ & n64680;
  assign n64771 = ~n64769 & ~n64770;
  assign n64772 = P2_P3_EAX_REG_17_ & n64766;
  assign n11601 = ~n64771 | n64772;
  assign n64774 = P2_P3_UWORD_REG_2_ & n64683;
  assign n64775 = P2_P3_DATAO_REG_18_ & n64680;
  assign n64776 = ~n64774 & ~n64775;
  assign n64777 = P2_P3_EAX_REG_18_ & n64766;
  assign n11606 = ~n64776 | n64777;
  assign n64779 = P2_P3_UWORD_REG_3_ & n64683;
  assign n64780 = P2_P3_DATAO_REG_19_ & n64680;
  assign n64781 = ~n64779 & ~n64780;
  assign n64782 = P2_P3_EAX_REG_19_ & n64766;
  assign n11611 = ~n64781 | n64782;
  assign n64784 = P2_P3_UWORD_REG_4_ & n64683;
  assign n64785 = P2_P3_DATAO_REG_20_ & n64680;
  assign n64786 = ~n64784 & ~n64785;
  assign n64787 = P2_P3_EAX_REG_20_ & n64766;
  assign n11616 = ~n64786 | n64787;
  assign n64789 = P2_P3_UWORD_REG_5_ & n64683;
  assign n64790 = P2_P3_DATAO_REG_21_ & n64680;
  assign n64791 = ~n64789 & ~n64790;
  assign n64792 = P2_P3_EAX_REG_21_ & n64766;
  assign n11621 = ~n64791 | n64792;
  assign n64794 = P2_P3_UWORD_REG_6_ & n64683;
  assign n64795 = P2_P3_DATAO_REG_22_ & n64680;
  assign n64796 = ~n64794 & ~n64795;
  assign n64797 = P2_P3_EAX_REG_22_ & n64766;
  assign n11626 = ~n64796 | n64797;
  assign n64799 = P2_P3_UWORD_REG_7_ & n64683;
  assign n64800 = P2_P3_DATAO_REG_23_ & n64680;
  assign n64801 = ~n64799 & ~n64800;
  assign n64802 = P2_P3_EAX_REG_23_ & n64766;
  assign n11631 = ~n64801 | n64802;
  assign n64804 = P2_P3_UWORD_REG_8_ & n64683;
  assign n64805 = P2_P3_DATAO_REG_24_ & n64680;
  assign n64806 = ~n64804 & ~n64805;
  assign n64807 = P2_P3_EAX_REG_24_ & n64766;
  assign n11636 = ~n64806 | n64807;
  assign n64809 = P2_P3_UWORD_REG_9_ & n64683;
  assign n64810 = P2_P3_DATAO_REG_25_ & n64680;
  assign n64811 = ~n64809 & ~n64810;
  assign n64812 = P2_P3_EAX_REG_25_ & n64766;
  assign n11641 = ~n64811 | n64812;
  assign n64814 = P2_P3_UWORD_REG_10_ & n64683;
  assign n64815 = P2_P3_DATAO_REG_26_ & n64680;
  assign n64816 = ~n64814 & ~n64815;
  assign n64817 = P2_P3_EAX_REG_26_ & n64766;
  assign n11646 = ~n64816 | n64817;
  assign n64819 = P2_P3_UWORD_REG_11_ & n64683;
  assign n64820 = P2_P3_DATAO_REG_27_ & n64680;
  assign n64821 = ~n64819 & ~n64820;
  assign n64822 = P2_P3_EAX_REG_27_ & n64766;
  assign n11651 = ~n64821 | n64822;
  assign n64824 = P2_P3_UWORD_REG_12_ & n64683;
  assign n64825 = P2_P3_DATAO_REG_28_ & n64680;
  assign n64826 = ~n64824 & ~n64825;
  assign n64827 = P2_P3_EAX_REG_28_ & n64766;
  assign n11656 = ~n64826 | n64827;
  assign n64829 = P2_P3_UWORD_REG_13_ & n64683;
  assign n64830 = P2_P3_DATAO_REG_29_ & n64680;
  assign n64831 = ~n64829 & ~n64830;
  assign n64832 = P2_P3_EAX_REG_29_ & n64766;
  assign n11661 = ~n64831 | n64832;
  assign n64834 = P2_P3_UWORD_REG_14_ & n64683;
  assign n64835 = P2_P3_DATAO_REG_30_ & n64680;
  assign n64836 = ~n64834 & ~n64835;
  assign n64837 = P2_P3_EAX_REG_30_ & n64766;
  assign n11666 = ~n64836 | n64837;
  assign n11671 = P2_P3_DATAO_REG_31_ & n64680;
  assign n64840 = n59201 & ~n59265;
  assign n64841 = n59321 & ~n64840;
  assign n64842 = n59055 & n64841;
  assign n64843 = ~n61031 & n64842;
  assign n64844 = ~n58838 & n64841;
  assign n64845 = ~n59055 & n64844;
  assign n64846 = P2_BUF2_REG_0_ & n64845;
  assign n64847 = P2_P3_EAX_REG_0_ & ~n64841;
  assign n64848 = n58838 & n64841;
  assign n64849 = ~P2_P3_EAX_REG_0_ & n64848;
  assign n64850 = ~n64847 & ~n64849;
  assign n64851 = ~n64843 & ~n64846;
  assign n11676 = ~n64850 | ~n64851;
  assign n64853 = ~n61149 & n64842;
  assign n64854 = P2_BUF2_REG_1_ & n64845;
  assign n64855 = P2_P3_EAX_REG_1_ & ~n64841;
  assign n64856 = ~P2_P3_EAX_REG_0_ & P2_P3_EAX_REG_1_;
  assign n64857 = P2_P3_EAX_REG_0_ & ~P2_P3_EAX_REG_1_;
  assign n64858 = ~n64856 & ~n64857;
  assign n64859 = n64848 & ~n64858;
  assign n64860 = ~n64855 & ~n64859;
  assign n64861 = ~n64853 & ~n64854;
  assign n11681 = ~n64860 | ~n64861;
  assign n64863 = ~n61269 & n64842;
  assign n64864 = P2_BUF2_REG_2_ & n64845;
  assign n64865 = P2_P3_EAX_REG_2_ & ~n64841;
  assign n64866 = P2_P3_EAX_REG_0_ & P2_P3_EAX_REG_1_;
  assign n64867 = ~P2_P3_EAX_REG_2_ & n64866;
  assign n64868 = P2_P3_EAX_REG_2_ & ~n64866;
  assign n64869 = ~n64867 & ~n64868;
  assign n64870 = n64848 & ~n64869;
  assign n64871 = ~n64865 & ~n64870;
  assign n64872 = ~n64863 & ~n64864;
  assign n11686 = ~n64871 | ~n64872;
  assign n64874 = ~n61393 & n64842;
  assign n64875 = P2_BUF2_REG_3_ & n64845;
  assign n64876 = P2_P3_EAX_REG_3_ & ~n64841;
  assign n64877 = P2_P3_EAX_REG_0_ & P2_P3_EAX_REG_2_;
  assign n64878 = P2_P3_EAX_REG_1_ & n64877;
  assign n64879 = P2_P3_EAX_REG_3_ & ~n64878;
  assign n64880 = ~P2_P3_EAX_REG_3_ & n64878;
  assign n64881 = ~n64879 & ~n64880;
  assign n64882 = n64848 & ~n64881;
  assign n64883 = ~n64876 & ~n64882;
  assign n64884 = ~n64874 & ~n64875;
  assign n11691 = ~n64883 | ~n64884;
  assign n64886 = ~n61520 & n64842;
  assign n64887 = P2_BUF2_REG_4_ & n64845;
  assign n64888 = P2_P3_EAX_REG_4_ & ~n64841;
  assign n64889 = P2_P3_EAX_REG_3_ & n64878;
  assign n64890 = ~P2_P3_EAX_REG_4_ & n64889;
  assign n64891 = P2_P3_EAX_REG_4_ & ~n64889;
  assign n64892 = ~n64890 & ~n64891;
  assign n64893 = n64848 & ~n64892;
  assign n64894 = ~n64888 & ~n64893;
  assign n64895 = ~n64886 & ~n64887;
  assign n11696 = ~n64894 | ~n64895;
  assign n64897 = ~n61661 & n64842;
  assign n64898 = P2_BUF2_REG_5_ & n64845;
  assign n64899 = P2_P3_EAX_REG_5_ & ~n64841;
  assign n64900 = P2_P3_EAX_REG_3_ & P2_P3_EAX_REG_4_;
  assign n64901 = n64878 & n64900;
  assign n64902 = P2_P3_EAX_REG_5_ & ~n64901;
  assign n64903 = ~P2_P3_EAX_REG_5_ & n64901;
  assign n64904 = ~n64902 & ~n64903;
  assign n64905 = n64848 & ~n64904;
  assign n64906 = ~n64899 & ~n64905;
  assign n64907 = ~n64897 & ~n64898;
  assign n11701 = ~n64906 | ~n64907;
  assign n64909 = ~n61793 & n64842;
  assign n64910 = P2_BUF2_REG_6_ & n64845;
  assign n64911 = P2_P3_EAX_REG_6_ & ~n64841;
  assign n64912 = P2_P3_EAX_REG_5_ & n64901;
  assign n64913 = ~P2_P3_EAX_REG_6_ & n64912;
  assign n64914 = P2_P3_EAX_REG_6_ & ~n64912;
  assign n64915 = ~n64913 & ~n64914;
  assign n64916 = n64848 & ~n64915;
  assign n64917 = ~n64911 & ~n64916;
  assign n64918 = ~n64909 & ~n64910;
  assign n11706 = ~n64917 | ~n64918;
  assign n64920 = ~n61065 & n64842;
  assign n64921 = P2_BUF2_REG_7_ & n64845;
  assign n64922 = P2_P3_EAX_REG_7_ & ~n64841;
  assign n64923 = P2_P3_EAX_REG_5_ & P2_P3_EAX_REG_6_;
  assign n64924 = n64901 & n64923;
  assign n64925 = P2_P3_EAX_REG_7_ & ~n64924;
  assign n64926 = ~P2_P3_EAX_REG_7_ & n64924;
  assign n64927 = ~n64925 & ~n64926;
  assign n64928 = n64848 & ~n64927;
  assign n64929 = ~n64922 & ~n64928;
  assign n64930 = ~n64920 & ~n64921;
  assign n11711 = ~n64929 | ~n64930;
  assign n64932 = ~n59215 & ~n59222;
  assign n64933 = ~n59166 & ~n64932;
  assign n64934 = n58696 & n64933;
  assign n64935 = P2_P3_INSTQUEUE_REG_15__0_ & n64934;
  assign n64936 = n58700 & n64933;
  assign n64937 = P2_P3_INSTQUEUE_REG_14__0_ & n64936;
  assign n64938 = n58687 & n64933;
  assign n64939 = P2_P3_INSTQUEUE_REG_13__0_ & n64938;
  assign n64940 = n58691 & n64933;
  assign n64941 = P2_P3_INSTQUEUE_REG_12__0_ & n64940;
  assign n64942 = ~n64935 & ~n64937;
  assign n64943 = ~n64939 & n64942;
  assign n64944 = ~n64941 & n64943;
  assign n64945 = n59166 & ~n64932;
  assign n64946 = n58696 & n64945;
  assign n64947 = P2_P3_INSTQUEUE_REG_11__0_ & n64946;
  assign n64948 = n58700 & n64945;
  assign n64949 = P2_P3_INSTQUEUE_REG_10__0_ & n64948;
  assign n64950 = n58687 & n64945;
  assign n64951 = P2_P3_INSTQUEUE_REG_9__0_ & n64950;
  assign n64952 = n58691 & n64945;
  assign n64953 = P2_P3_INSTQUEUE_REG_8__0_ & n64952;
  assign n64954 = ~n64947 & ~n64949;
  assign n64955 = ~n64951 & n64954;
  assign n64956 = ~n64953 & n64955;
  assign n64957 = ~n59166 & n64932;
  assign n64958 = n58696 & n64957;
  assign n64959 = P2_P3_INSTQUEUE_REG_7__0_ & n64958;
  assign n64960 = n58700 & n64957;
  assign n64961 = P2_P3_INSTQUEUE_REG_6__0_ & n64960;
  assign n64962 = n58687 & n64957;
  assign n64963 = P2_P3_INSTQUEUE_REG_5__0_ & n64962;
  assign n64964 = n58691 & n64957;
  assign n64965 = P2_P3_INSTQUEUE_REG_4__0_ & n64964;
  assign n64966 = ~n64959 & ~n64961;
  assign n64967 = ~n64963 & n64966;
  assign n64968 = ~n64965 & n64967;
  assign n64969 = n59166 & n64932;
  assign n64970 = n58696 & n64969;
  assign n64971 = P2_P3_INSTQUEUE_REG_3__0_ & n64970;
  assign n64972 = n58700 & n64969;
  assign n64973 = P2_P3_INSTQUEUE_REG_2__0_ & n64972;
  assign n64974 = n58687 & n64969;
  assign n64975 = P2_P3_INSTQUEUE_REG_1__0_ & n64974;
  assign n64976 = n58691 & n64969;
  assign n64977 = P2_P3_INSTQUEUE_REG_0__0_ & n64976;
  assign n64978 = ~n64971 & ~n64973;
  assign n64979 = ~n64975 & n64978;
  assign n64980 = ~n64977 & n64979;
  assign n64981 = n64944 & n64956;
  assign n64982 = n64968 & n64981;
  assign n64983 = n64980 & n64982;
  assign n64984 = n64842 & ~n64983;
  assign n64985 = P2_BUF2_REG_8_ & n64845;
  assign n64986 = P2_P3_EAX_REG_8_ & ~n64841;
  assign n64987 = P2_P3_EAX_REG_7_ & n64924;
  assign n64988 = ~P2_P3_EAX_REG_8_ & n64987;
  assign n64989 = P2_P3_EAX_REG_8_ & ~n64987;
  assign n64990 = ~n64988 & ~n64989;
  assign n64991 = n64848 & ~n64990;
  assign n64992 = ~n64986 & ~n64991;
  assign n64993 = ~n64984 & ~n64985;
  assign n11716 = ~n64992 | ~n64993;
  assign n64995 = P2_P3_INSTQUEUE_REG_15__1_ & n64934;
  assign n64996 = P2_P3_INSTQUEUE_REG_14__1_ & n64936;
  assign n64997 = P2_P3_INSTQUEUE_REG_13__1_ & n64938;
  assign n64998 = P2_P3_INSTQUEUE_REG_12__1_ & n64940;
  assign n64999 = ~n64995 & ~n64996;
  assign n65000 = ~n64997 & n64999;
  assign n65001 = ~n64998 & n65000;
  assign n65002 = P2_P3_INSTQUEUE_REG_11__1_ & n64946;
  assign n65003 = P2_P3_INSTQUEUE_REG_10__1_ & n64948;
  assign n65004 = P2_P3_INSTQUEUE_REG_9__1_ & n64950;
  assign n65005 = P2_P3_INSTQUEUE_REG_8__1_ & n64952;
  assign n65006 = ~n65002 & ~n65003;
  assign n65007 = ~n65004 & n65006;
  assign n65008 = ~n65005 & n65007;
  assign n65009 = P2_P3_INSTQUEUE_REG_7__1_ & n64958;
  assign n65010 = P2_P3_INSTQUEUE_REG_6__1_ & n64960;
  assign n65011 = P2_P3_INSTQUEUE_REG_5__1_ & n64962;
  assign n65012 = P2_P3_INSTQUEUE_REG_4__1_ & n64964;
  assign n65013 = ~n65009 & ~n65010;
  assign n65014 = ~n65011 & n65013;
  assign n65015 = ~n65012 & n65014;
  assign n65016 = P2_P3_INSTQUEUE_REG_3__1_ & n64970;
  assign n65017 = P2_P3_INSTQUEUE_REG_2__1_ & n64972;
  assign n65018 = P2_P3_INSTQUEUE_REG_1__1_ & n64974;
  assign n65019 = P2_P3_INSTQUEUE_REG_0__1_ & n64976;
  assign n65020 = ~n65016 & ~n65017;
  assign n65021 = ~n65018 & n65020;
  assign n65022 = ~n65019 & n65021;
  assign n65023 = n65001 & n65008;
  assign n65024 = n65015 & n65023;
  assign n65025 = n65022 & n65024;
  assign n65026 = n64842 & ~n65025;
  assign n65027 = P2_BUF2_REG_9_ & n64845;
  assign n65028 = P2_P3_EAX_REG_9_ & ~n64841;
  assign n65029 = P2_P3_EAX_REG_7_ & P2_P3_EAX_REG_8_;
  assign n65030 = n64924 & n65029;
  assign n65031 = P2_P3_EAX_REG_9_ & ~n65030;
  assign n65032 = ~P2_P3_EAX_REG_9_ & n65030;
  assign n65033 = ~n65031 & ~n65032;
  assign n65034 = n64848 & ~n65033;
  assign n65035 = ~n65028 & ~n65034;
  assign n65036 = ~n65026 & ~n65027;
  assign n11721 = ~n65035 | ~n65036;
  assign n65038 = P2_P3_INSTQUEUE_REG_15__2_ & n64934;
  assign n65039 = P2_P3_INSTQUEUE_REG_14__2_ & n64936;
  assign n65040 = P2_P3_INSTQUEUE_REG_13__2_ & n64938;
  assign n65041 = P2_P3_INSTQUEUE_REG_12__2_ & n64940;
  assign n65042 = ~n65038 & ~n65039;
  assign n65043 = ~n65040 & n65042;
  assign n65044 = ~n65041 & n65043;
  assign n65045 = P2_P3_INSTQUEUE_REG_11__2_ & n64946;
  assign n65046 = P2_P3_INSTQUEUE_REG_10__2_ & n64948;
  assign n65047 = P2_P3_INSTQUEUE_REG_9__2_ & n64950;
  assign n65048 = P2_P3_INSTQUEUE_REG_8__2_ & n64952;
  assign n65049 = ~n65045 & ~n65046;
  assign n65050 = ~n65047 & n65049;
  assign n65051 = ~n65048 & n65050;
  assign n65052 = P2_P3_INSTQUEUE_REG_7__2_ & n64958;
  assign n65053 = P2_P3_INSTQUEUE_REG_6__2_ & n64960;
  assign n65054 = P2_P3_INSTQUEUE_REG_5__2_ & n64962;
  assign n65055 = P2_P3_INSTQUEUE_REG_4__2_ & n64964;
  assign n65056 = ~n65052 & ~n65053;
  assign n65057 = ~n65054 & n65056;
  assign n65058 = ~n65055 & n65057;
  assign n65059 = P2_P3_INSTQUEUE_REG_3__2_ & n64970;
  assign n65060 = P2_P3_INSTQUEUE_REG_2__2_ & n64972;
  assign n65061 = P2_P3_INSTQUEUE_REG_1__2_ & n64974;
  assign n65062 = P2_P3_INSTQUEUE_REG_0__2_ & n64976;
  assign n65063 = ~n65059 & ~n65060;
  assign n65064 = ~n65061 & n65063;
  assign n65065 = ~n65062 & n65064;
  assign n65066 = n65044 & n65051;
  assign n65067 = n65058 & n65066;
  assign n65068 = n65065 & n65067;
  assign n65069 = n64842 & ~n65068;
  assign n65070 = P2_BUF2_REG_10_ & n64845;
  assign n65071 = P2_P3_EAX_REG_10_ & ~n64841;
  assign n65072 = P2_P3_EAX_REG_9_ & n65030;
  assign n65073 = ~P2_P3_EAX_REG_10_ & n65072;
  assign n65074 = P2_P3_EAX_REG_10_ & ~n65072;
  assign n65075 = ~n65073 & ~n65074;
  assign n65076 = n64848 & ~n65075;
  assign n65077 = ~n65071 & ~n65076;
  assign n65078 = ~n65069 & ~n65070;
  assign n11726 = ~n65077 | ~n65078;
  assign n65080 = P2_P3_INSTQUEUE_REG_15__3_ & n64934;
  assign n65081 = P2_P3_INSTQUEUE_REG_14__3_ & n64936;
  assign n65082 = P2_P3_INSTQUEUE_REG_13__3_ & n64938;
  assign n65083 = P2_P3_INSTQUEUE_REG_12__3_ & n64940;
  assign n65084 = ~n65080 & ~n65081;
  assign n65085 = ~n65082 & n65084;
  assign n65086 = ~n65083 & n65085;
  assign n65087 = P2_P3_INSTQUEUE_REG_11__3_ & n64946;
  assign n65088 = P2_P3_INSTQUEUE_REG_10__3_ & n64948;
  assign n65089 = P2_P3_INSTQUEUE_REG_9__3_ & n64950;
  assign n65090 = P2_P3_INSTQUEUE_REG_8__3_ & n64952;
  assign n65091 = ~n65087 & ~n65088;
  assign n65092 = ~n65089 & n65091;
  assign n65093 = ~n65090 & n65092;
  assign n65094 = P2_P3_INSTQUEUE_REG_7__3_ & n64958;
  assign n65095 = P2_P3_INSTQUEUE_REG_6__3_ & n64960;
  assign n65096 = P2_P3_INSTQUEUE_REG_5__3_ & n64962;
  assign n65097 = P2_P3_INSTQUEUE_REG_4__3_ & n64964;
  assign n65098 = ~n65094 & ~n65095;
  assign n65099 = ~n65096 & n65098;
  assign n65100 = ~n65097 & n65099;
  assign n65101 = P2_P3_INSTQUEUE_REG_3__3_ & n64970;
  assign n65102 = P2_P3_INSTQUEUE_REG_2__3_ & n64972;
  assign n65103 = P2_P3_INSTQUEUE_REG_1__3_ & n64974;
  assign n65104 = P2_P3_INSTQUEUE_REG_0__3_ & n64976;
  assign n65105 = ~n65101 & ~n65102;
  assign n65106 = ~n65103 & n65105;
  assign n65107 = ~n65104 & n65106;
  assign n65108 = n65086 & n65093;
  assign n65109 = n65100 & n65108;
  assign n65110 = n65107 & n65109;
  assign n65111 = n64842 & ~n65110;
  assign n65112 = P2_BUF2_REG_11_ & n64845;
  assign n65113 = P2_P3_EAX_REG_11_ & ~n64841;
  assign n65114 = P2_P3_EAX_REG_9_ & P2_P3_EAX_REG_10_;
  assign n65115 = n65030 & n65114;
  assign n65116 = P2_P3_EAX_REG_11_ & ~n65115;
  assign n65117 = ~P2_P3_EAX_REG_11_ & n65115;
  assign n65118 = ~n65116 & ~n65117;
  assign n65119 = n64848 & ~n65118;
  assign n65120 = ~n65113 & ~n65119;
  assign n65121 = ~n65111 & ~n65112;
  assign n11731 = ~n65120 | ~n65121;
  assign n65123 = P2_P3_INSTQUEUE_REG_15__4_ & n64934;
  assign n65124 = P2_P3_INSTQUEUE_REG_14__4_ & n64936;
  assign n65125 = P2_P3_INSTQUEUE_REG_13__4_ & n64938;
  assign n65126 = P2_P3_INSTQUEUE_REG_12__4_ & n64940;
  assign n65127 = ~n65123 & ~n65124;
  assign n65128 = ~n65125 & n65127;
  assign n65129 = ~n65126 & n65128;
  assign n65130 = P2_P3_INSTQUEUE_REG_11__4_ & n64946;
  assign n65131 = P2_P3_INSTQUEUE_REG_10__4_ & n64948;
  assign n65132 = P2_P3_INSTQUEUE_REG_9__4_ & n64950;
  assign n65133 = P2_P3_INSTQUEUE_REG_8__4_ & n64952;
  assign n65134 = ~n65130 & ~n65131;
  assign n65135 = ~n65132 & n65134;
  assign n65136 = ~n65133 & n65135;
  assign n65137 = P2_P3_INSTQUEUE_REG_7__4_ & n64958;
  assign n65138 = P2_P3_INSTQUEUE_REG_6__4_ & n64960;
  assign n65139 = P2_P3_INSTQUEUE_REG_5__4_ & n64962;
  assign n65140 = P2_P3_INSTQUEUE_REG_4__4_ & n64964;
  assign n65141 = ~n65137 & ~n65138;
  assign n65142 = ~n65139 & n65141;
  assign n65143 = ~n65140 & n65142;
  assign n65144 = P2_P3_INSTQUEUE_REG_3__4_ & n64970;
  assign n65145 = P2_P3_INSTQUEUE_REG_2__4_ & n64972;
  assign n65146 = P2_P3_INSTQUEUE_REG_1__4_ & n64974;
  assign n65147 = P2_P3_INSTQUEUE_REG_0__4_ & n64976;
  assign n65148 = ~n65144 & ~n65145;
  assign n65149 = ~n65146 & n65148;
  assign n65150 = ~n65147 & n65149;
  assign n65151 = n65129 & n65136;
  assign n65152 = n65143 & n65151;
  assign n65153 = n65150 & n65152;
  assign n65154 = n64842 & ~n65153;
  assign n65155 = P2_BUF2_REG_12_ & n64845;
  assign n65156 = P2_P3_EAX_REG_12_ & ~n64841;
  assign n65157 = P2_P3_EAX_REG_11_ & n65115;
  assign n65158 = ~P2_P3_EAX_REG_12_ & n65157;
  assign n65159 = P2_P3_EAX_REG_12_ & ~n65157;
  assign n65160 = ~n65158 & ~n65159;
  assign n65161 = n64848 & ~n65160;
  assign n65162 = ~n65156 & ~n65161;
  assign n65163 = ~n65154 & ~n65155;
  assign n11736 = ~n65162 | ~n65163;
  assign n65165 = P2_BUF2_REG_13_ & n64845;
  assign n65166 = P2_P3_INSTQUEUE_REG_15__5_ & n64934;
  assign n65167 = P2_P3_INSTQUEUE_REG_14__5_ & n64936;
  assign n65168 = P2_P3_INSTQUEUE_REG_13__5_ & n64938;
  assign n65169 = P2_P3_INSTQUEUE_REG_12__5_ & n64940;
  assign n65170 = ~n65166 & ~n65167;
  assign n65171 = ~n65168 & n65170;
  assign n65172 = ~n65169 & n65171;
  assign n65173 = P2_P3_INSTQUEUE_REG_11__5_ & n64946;
  assign n65174 = P2_P3_INSTQUEUE_REG_10__5_ & n64948;
  assign n65175 = P2_P3_INSTQUEUE_REG_9__5_ & n64950;
  assign n65176 = P2_P3_INSTQUEUE_REG_8__5_ & n64952;
  assign n65177 = ~n65173 & ~n65174;
  assign n65178 = ~n65175 & n65177;
  assign n65179 = ~n65176 & n65178;
  assign n65180 = P2_P3_INSTQUEUE_REG_7__5_ & n64958;
  assign n65181 = P2_P3_INSTQUEUE_REG_6__5_ & n64960;
  assign n65182 = P2_P3_INSTQUEUE_REG_5__5_ & n64962;
  assign n65183 = P2_P3_INSTQUEUE_REG_4__5_ & n64964;
  assign n65184 = ~n65180 & ~n65181;
  assign n65185 = ~n65182 & n65184;
  assign n65186 = ~n65183 & n65185;
  assign n65187 = P2_P3_INSTQUEUE_REG_3__5_ & n64970;
  assign n65188 = P2_P3_INSTQUEUE_REG_2__5_ & n64972;
  assign n65189 = P2_P3_INSTQUEUE_REG_1__5_ & n64974;
  assign n65190 = P2_P3_INSTQUEUE_REG_0__5_ & n64976;
  assign n65191 = ~n65187 & ~n65188;
  assign n65192 = ~n65189 & n65191;
  assign n65193 = ~n65190 & n65192;
  assign n65194 = n65172 & n65179;
  assign n65195 = n65186 & n65194;
  assign n65196 = n65193 & n65195;
  assign n65197 = n64842 & ~n65196;
  assign n65198 = P2_P3_EAX_REG_13_ & ~n64841;
  assign n65199 = ~n65197 & ~n65198;
  assign n65200 = P2_P3_EAX_REG_11_ & P2_P3_EAX_REG_12_;
  assign n65201 = n65115 & n65200;
  assign n65202 = P2_P3_EAX_REG_13_ & ~n65201;
  assign n65203 = ~P2_P3_EAX_REG_13_ & n65201;
  assign n65204 = ~n65202 & ~n65203;
  assign n65205 = n64848 & ~n65204;
  assign n65206 = ~n65165 & n65199;
  assign n11741 = n65205 | ~n65206;
  assign n65208 = P2_BUF2_REG_14_ & n64845;
  assign n65209 = P2_P3_INSTQUEUE_REG_15__6_ & n64934;
  assign n65210 = P2_P3_INSTQUEUE_REG_14__6_ & n64936;
  assign n65211 = P2_P3_INSTQUEUE_REG_13__6_ & n64938;
  assign n65212 = P2_P3_INSTQUEUE_REG_12__6_ & n64940;
  assign n65213 = ~n65209 & ~n65210;
  assign n65214 = ~n65211 & n65213;
  assign n65215 = ~n65212 & n65214;
  assign n65216 = P2_P3_INSTQUEUE_REG_11__6_ & n64946;
  assign n65217 = P2_P3_INSTQUEUE_REG_10__6_ & n64948;
  assign n65218 = P2_P3_INSTQUEUE_REG_9__6_ & n64950;
  assign n65219 = P2_P3_INSTQUEUE_REG_8__6_ & n64952;
  assign n65220 = ~n65216 & ~n65217;
  assign n65221 = ~n65218 & n65220;
  assign n65222 = ~n65219 & n65221;
  assign n65223 = P2_P3_INSTQUEUE_REG_7__6_ & n64958;
  assign n65224 = P2_P3_INSTQUEUE_REG_6__6_ & n64960;
  assign n65225 = P2_P3_INSTQUEUE_REG_5__6_ & n64962;
  assign n65226 = P2_P3_INSTQUEUE_REG_4__6_ & n64964;
  assign n65227 = ~n65223 & ~n65224;
  assign n65228 = ~n65225 & n65227;
  assign n65229 = ~n65226 & n65228;
  assign n65230 = P2_P3_INSTQUEUE_REG_3__6_ & n64970;
  assign n65231 = P2_P3_INSTQUEUE_REG_2__6_ & n64972;
  assign n65232 = P2_P3_INSTQUEUE_REG_1__6_ & n64974;
  assign n65233 = P2_P3_INSTQUEUE_REG_0__6_ & n64976;
  assign n65234 = ~n65230 & ~n65231;
  assign n65235 = ~n65232 & n65234;
  assign n65236 = ~n65233 & n65235;
  assign n65237 = n65215 & n65222;
  assign n65238 = n65229 & n65237;
  assign n65239 = n65236 & n65238;
  assign n65240 = n64842 & ~n65239;
  assign n65241 = P2_P3_EAX_REG_14_ & ~n64841;
  assign n65242 = ~n65240 & ~n65241;
  assign n65243 = P2_P3_EAX_REG_13_ & n65201;
  assign n65244 = ~P2_P3_EAX_REG_14_ & n65243;
  assign n65245 = P2_P3_EAX_REG_14_ & ~n65243;
  assign n65246 = ~n65244 & ~n65245;
  assign n65247 = n64848 & ~n65246;
  assign n65248 = ~n65208 & n65242;
  assign n11746 = n65247 | ~n65248;
  assign n65250 = P2_BUF2_REG_15_ & n64845;
  assign n65251 = P2_P3_INSTQUEUE_REG_15__7_ & n64934;
  assign n65252 = P2_P3_INSTQUEUE_REG_14__7_ & n64936;
  assign n65253 = P2_P3_INSTQUEUE_REG_13__7_ & n64938;
  assign n65254 = P2_P3_INSTQUEUE_REG_12__7_ & n64940;
  assign n65255 = ~n65251 & ~n65252;
  assign n65256 = ~n65253 & n65255;
  assign n65257 = ~n65254 & n65256;
  assign n65258 = P2_P3_INSTQUEUE_REG_11__7_ & n64946;
  assign n65259 = P2_P3_INSTQUEUE_REG_10__7_ & n64948;
  assign n65260 = P2_P3_INSTQUEUE_REG_9__7_ & n64950;
  assign n65261 = P2_P3_INSTQUEUE_REG_8__7_ & n64952;
  assign n65262 = ~n65258 & ~n65259;
  assign n65263 = ~n65260 & n65262;
  assign n65264 = ~n65261 & n65263;
  assign n65265 = P2_P3_INSTQUEUE_REG_7__7_ & n64958;
  assign n65266 = P2_P3_INSTQUEUE_REG_6__7_ & n64960;
  assign n65267 = P2_P3_INSTQUEUE_REG_5__7_ & n64962;
  assign n65268 = P2_P3_INSTQUEUE_REG_4__7_ & n64964;
  assign n65269 = ~n65265 & ~n65266;
  assign n65270 = ~n65267 & n65269;
  assign n65271 = ~n65268 & n65270;
  assign n65272 = P2_P3_INSTQUEUE_REG_3__7_ & n64970;
  assign n65273 = P2_P3_INSTQUEUE_REG_2__7_ & n64972;
  assign n65274 = P2_P3_INSTQUEUE_REG_1__7_ & n64974;
  assign n65275 = P2_P3_INSTQUEUE_REG_0__7_ & n64976;
  assign n65276 = ~n65272 & ~n65273;
  assign n65277 = ~n65274 & n65276;
  assign n65278 = ~n65275 & n65277;
  assign n65279 = n65257 & n65264;
  assign n65280 = n65271 & n65279;
  assign n65281 = n65278 & n65280;
  assign n65282 = n64842 & ~n65281;
  assign n65283 = P2_P3_EAX_REG_15_ & ~n64841;
  assign n65284 = ~n65282 & ~n65283;
  assign n65285 = P2_P3_EAX_REG_13_ & P2_P3_EAX_REG_14_;
  assign n65286 = n65201 & n65285;
  assign n65287 = P2_P3_EAX_REG_15_ & ~n65286;
  assign n65288 = ~P2_P3_EAX_REG_15_ & n65286;
  assign n65289 = ~n65287 & ~n65288;
  assign n65290 = n64848 & ~n65289;
  assign n65291 = ~n65250 & n65284;
  assign n11751 = n65290 | ~n65291;
  assign n65293 = ~n58775 & n64844;
  assign n65294 = P2_BUF2_REG_16_ & n65293;
  assign n65295 = n58744 & n64844;
  assign n65296 = P2_BUF2_REG_0_ & n65295;
  assign n65297 = P2_P3_EAX_REG_16_ & ~n64841;
  assign n65298 = P2_P3_INSTQUEUERD_ADDR_REG_2_ & ~n58700;
  assign n65299 = ~P2_P3_INSTQUEUERD_ADDR_REG_3_ & n65298;
  assign n65300 = P2_P3_INSTQUEUERD_ADDR_REG_3_ & ~n65298;
  assign n65301 = ~n65299 & ~n65300;
  assign n65302 = ~n58701 & ~n65298;
  assign n65303 = n65301 & n65302;
  assign n65304 = n60981 & n65303;
  assign n65305 = P2_P3_INSTQUEUE_REG_7__0_ & n65304;
  assign n65306 = n60978 & n65303;
  assign n65307 = P2_P3_INSTQUEUE_REG_6__0_ & n65306;
  assign n65308 = n60987 & n65303;
  assign n65309 = P2_P3_INSTQUEUE_REG_5__0_ & n65308;
  assign n65310 = n60984 & n65303;
  assign n65311 = P2_P3_INSTQUEUE_REG_4__0_ & n65310;
  assign n65312 = ~n65305 & ~n65307;
  assign n65313 = ~n65309 & n65312;
  assign n65314 = ~n65311 & n65313;
  assign n65315 = n65301 & ~n65302;
  assign n65316 = n60981 & n65315;
  assign n65317 = P2_P3_INSTQUEUE_REG_3__0_ & n65316;
  assign n65318 = n60978 & n65315;
  assign n65319 = P2_P3_INSTQUEUE_REG_2__0_ & n65318;
  assign n65320 = n60987 & n65315;
  assign n65321 = P2_P3_INSTQUEUE_REG_1__0_ & n65320;
  assign n65322 = n60984 & n65315;
  assign n65323 = P2_P3_INSTQUEUE_REG_0__0_ & n65322;
  assign n65324 = ~n65317 & ~n65319;
  assign n65325 = ~n65321 & n65324;
  assign n65326 = ~n65323 & n65325;
  assign n65327 = ~n65301 & n65302;
  assign n65328 = n60981 & n65327;
  assign n65329 = P2_P3_INSTQUEUE_REG_15__0_ & n65328;
  assign n65330 = n60978 & n65327;
  assign n65331 = P2_P3_INSTQUEUE_REG_14__0_ & n65330;
  assign n65332 = n60987 & n65327;
  assign n65333 = P2_P3_INSTQUEUE_REG_13__0_ & n65332;
  assign n65334 = n60984 & n65327;
  assign n65335 = P2_P3_INSTQUEUE_REG_12__0_ & n65334;
  assign n65336 = ~n65329 & ~n65331;
  assign n65337 = ~n65333 & n65336;
  assign n65338 = ~n65335 & n65337;
  assign n65339 = ~n65301 & ~n65302;
  assign n65340 = n60981 & n65339;
  assign n65341 = P2_P3_INSTQUEUE_REG_11__0_ & n65340;
  assign n65342 = n60978 & n65339;
  assign n65343 = P2_P3_INSTQUEUE_REG_10__0_ & n65342;
  assign n65344 = n60987 & n65339;
  assign n65345 = P2_P3_INSTQUEUE_REG_9__0_ & n65344;
  assign n65346 = n60984 & n65339;
  assign n65347 = P2_P3_INSTQUEUE_REG_8__0_ & n65346;
  assign n65348 = ~n65341 & ~n65343;
  assign n65349 = ~n65345 & n65348;
  assign n65350 = ~n65347 & n65349;
  assign n65351 = n65314 & n65326;
  assign n65352 = n65338 & n65351;
  assign n65353 = n65350 & n65352;
  assign n65354 = n64842 & ~n65353;
  assign n65355 = ~n65297 & ~n65354;
  assign n65356 = P2_P3_EAX_REG_15_ & n65286;
  assign n65357 = ~P2_P3_EAX_REG_16_ & n65356;
  assign n65358 = P2_P3_EAX_REG_16_ & ~n65356;
  assign n65359 = ~n65357 & ~n65358;
  assign n65360 = n64848 & ~n65359;
  assign n65361 = ~n65294 & ~n65296;
  assign n65362 = n65355 & n65361;
  assign n11756 = n65360 | ~n65362;
  assign n65364 = P2_BUF2_REG_17_ & n65293;
  assign n65365 = P2_BUF2_REG_1_ & n65295;
  assign n65366 = P2_P3_EAX_REG_17_ & ~n64841;
  assign n65367 = P2_P3_INSTQUEUE_REG_7__1_ & n65304;
  assign n65368 = P2_P3_INSTQUEUE_REG_6__1_ & n65306;
  assign n65369 = P2_P3_INSTQUEUE_REG_5__1_ & n65308;
  assign n65370 = P2_P3_INSTQUEUE_REG_4__1_ & n65310;
  assign n65371 = ~n65367 & ~n65368;
  assign n65372 = ~n65369 & n65371;
  assign n65373 = ~n65370 & n65372;
  assign n65374 = P2_P3_INSTQUEUE_REG_3__1_ & n65316;
  assign n65375 = P2_P3_INSTQUEUE_REG_2__1_ & n65318;
  assign n65376 = P2_P3_INSTQUEUE_REG_1__1_ & n65320;
  assign n65377 = P2_P3_INSTQUEUE_REG_0__1_ & n65322;
  assign n65378 = ~n65374 & ~n65375;
  assign n65379 = ~n65376 & n65378;
  assign n65380 = ~n65377 & n65379;
  assign n65381 = P2_P3_INSTQUEUE_REG_15__1_ & n65328;
  assign n65382 = P2_P3_INSTQUEUE_REG_14__1_ & n65330;
  assign n65383 = P2_P3_INSTQUEUE_REG_13__1_ & n65332;
  assign n65384 = P2_P3_INSTQUEUE_REG_12__1_ & n65334;
  assign n65385 = ~n65381 & ~n65382;
  assign n65386 = ~n65383 & n65385;
  assign n65387 = ~n65384 & n65386;
  assign n65388 = P2_P3_INSTQUEUE_REG_11__1_ & n65340;
  assign n65389 = P2_P3_INSTQUEUE_REG_10__1_ & n65342;
  assign n65390 = P2_P3_INSTQUEUE_REG_9__1_ & n65344;
  assign n65391 = P2_P3_INSTQUEUE_REG_8__1_ & n65346;
  assign n65392 = ~n65388 & ~n65389;
  assign n65393 = ~n65390 & n65392;
  assign n65394 = ~n65391 & n65393;
  assign n65395 = n65373 & n65380;
  assign n65396 = n65387 & n65395;
  assign n65397 = n65394 & n65396;
  assign n65398 = n64842 & ~n65397;
  assign n65399 = ~n65366 & ~n65398;
  assign n65400 = P2_P3_EAX_REG_15_ & P2_P3_EAX_REG_16_;
  assign n65401 = n65286 & n65400;
  assign n65402 = P2_P3_EAX_REG_17_ & ~n65401;
  assign n65403 = ~P2_P3_EAX_REG_17_ & n65401;
  assign n65404 = ~n65402 & ~n65403;
  assign n65405 = n64848 & ~n65404;
  assign n65406 = ~n65364 & ~n65365;
  assign n65407 = n65399 & n65406;
  assign n11761 = n65405 | ~n65407;
  assign n65409 = P2_BUF2_REG_18_ & n65293;
  assign n65410 = P2_BUF2_REG_2_ & n65295;
  assign n65411 = P2_P3_EAX_REG_18_ & ~n64841;
  assign n65412 = P2_P3_INSTQUEUE_REG_7__2_ & n65304;
  assign n65413 = P2_P3_INSTQUEUE_REG_6__2_ & n65306;
  assign n65414 = P2_P3_INSTQUEUE_REG_5__2_ & n65308;
  assign n65415 = P2_P3_INSTQUEUE_REG_4__2_ & n65310;
  assign n65416 = ~n65412 & ~n65413;
  assign n65417 = ~n65414 & n65416;
  assign n65418 = ~n65415 & n65417;
  assign n65419 = P2_P3_INSTQUEUE_REG_3__2_ & n65316;
  assign n65420 = P2_P3_INSTQUEUE_REG_2__2_ & n65318;
  assign n65421 = P2_P3_INSTQUEUE_REG_1__2_ & n65320;
  assign n65422 = P2_P3_INSTQUEUE_REG_0__2_ & n65322;
  assign n65423 = ~n65419 & ~n65420;
  assign n65424 = ~n65421 & n65423;
  assign n65425 = ~n65422 & n65424;
  assign n65426 = P2_P3_INSTQUEUE_REG_15__2_ & n65328;
  assign n65427 = P2_P3_INSTQUEUE_REG_14__2_ & n65330;
  assign n65428 = P2_P3_INSTQUEUE_REG_13__2_ & n65332;
  assign n65429 = P2_P3_INSTQUEUE_REG_12__2_ & n65334;
  assign n65430 = ~n65426 & ~n65427;
  assign n65431 = ~n65428 & n65430;
  assign n65432 = ~n65429 & n65431;
  assign n65433 = P2_P3_INSTQUEUE_REG_11__2_ & n65340;
  assign n65434 = P2_P3_INSTQUEUE_REG_10__2_ & n65342;
  assign n65435 = P2_P3_INSTQUEUE_REG_9__2_ & n65344;
  assign n65436 = P2_P3_INSTQUEUE_REG_8__2_ & n65346;
  assign n65437 = ~n65433 & ~n65434;
  assign n65438 = ~n65435 & n65437;
  assign n65439 = ~n65436 & n65438;
  assign n65440 = n65418 & n65425;
  assign n65441 = n65432 & n65440;
  assign n65442 = n65439 & n65441;
  assign n65443 = n64842 & ~n65442;
  assign n65444 = ~n65411 & ~n65443;
  assign n65445 = P2_P3_EAX_REG_17_ & n65401;
  assign n65446 = ~P2_P3_EAX_REG_18_ & n65445;
  assign n65447 = P2_P3_EAX_REG_18_ & ~n65445;
  assign n65448 = ~n65446 & ~n65447;
  assign n65449 = n64848 & ~n65448;
  assign n65450 = ~n65409 & ~n65410;
  assign n65451 = n65444 & n65450;
  assign n11766 = n65449 | ~n65451;
  assign n65453 = P2_BUF2_REG_19_ & n65293;
  assign n65454 = P2_BUF2_REG_3_ & n65295;
  assign n65455 = P2_P3_EAX_REG_19_ & ~n64841;
  assign n65456 = P2_P3_INSTQUEUE_REG_7__3_ & n65304;
  assign n65457 = P2_P3_INSTQUEUE_REG_6__3_ & n65306;
  assign n65458 = P2_P3_INSTQUEUE_REG_5__3_ & n65308;
  assign n65459 = P2_P3_INSTQUEUE_REG_4__3_ & n65310;
  assign n65460 = ~n65456 & ~n65457;
  assign n65461 = ~n65458 & n65460;
  assign n65462 = ~n65459 & n65461;
  assign n65463 = P2_P3_INSTQUEUE_REG_3__3_ & n65316;
  assign n65464 = P2_P3_INSTQUEUE_REG_2__3_ & n65318;
  assign n65465 = P2_P3_INSTQUEUE_REG_1__3_ & n65320;
  assign n65466 = P2_P3_INSTQUEUE_REG_0__3_ & n65322;
  assign n65467 = ~n65463 & ~n65464;
  assign n65468 = ~n65465 & n65467;
  assign n65469 = ~n65466 & n65468;
  assign n65470 = P2_P3_INSTQUEUE_REG_15__3_ & n65328;
  assign n65471 = P2_P3_INSTQUEUE_REG_14__3_ & n65330;
  assign n65472 = P2_P3_INSTQUEUE_REG_13__3_ & n65332;
  assign n65473 = P2_P3_INSTQUEUE_REG_12__3_ & n65334;
  assign n65474 = ~n65470 & ~n65471;
  assign n65475 = ~n65472 & n65474;
  assign n65476 = ~n65473 & n65475;
  assign n65477 = P2_P3_INSTQUEUE_REG_11__3_ & n65340;
  assign n65478 = P2_P3_INSTQUEUE_REG_10__3_ & n65342;
  assign n65479 = P2_P3_INSTQUEUE_REG_9__3_ & n65344;
  assign n65480 = P2_P3_INSTQUEUE_REG_8__3_ & n65346;
  assign n65481 = ~n65477 & ~n65478;
  assign n65482 = ~n65479 & n65481;
  assign n65483 = ~n65480 & n65482;
  assign n65484 = n65462 & n65469;
  assign n65485 = n65476 & n65484;
  assign n65486 = n65483 & n65485;
  assign n65487 = n64842 & ~n65486;
  assign n65488 = ~n65455 & ~n65487;
  assign n65489 = P2_P3_EAX_REG_17_ & P2_P3_EAX_REG_18_;
  assign n65490 = n65401 & n65489;
  assign n65491 = P2_P3_EAX_REG_19_ & ~n65490;
  assign n65492 = ~P2_P3_EAX_REG_19_ & n65490;
  assign n65493 = ~n65491 & ~n65492;
  assign n65494 = n64848 & ~n65493;
  assign n65495 = ~n65453 & ~n65454;
  assign n65496 = n65488 & n65495;
  assign n11771 = n65494 | ~n65496;
  assign n65498 = P2_BUF2_REG_20_ & n65293;
  assign n65499 = P2_BUF2_REG_4_ & n65295;
  assign n65500 = P2_P3_EAX_REG_20_ & ~n64841;
  assign n65501 = P2_P3_INSTQUEUE_REG_7__4_ & n65304;
  assign n65502 = P2_P3_INSTQUEUE_REG_6__4_ & n65306;
  assign n65503 = P2_P3_INSTQUEUE_REG_5__4_ & n65308;
  assign n65504 = P2_P3_INSTQUEUE_REG_4__4_ & n65310;
  assign n65505 = ~n65501 & ~n65502;
  assign n65506 = ~n65503 & n65505;
  assign n65507 = ~n65504 & n65506;
  assign n65508 = P2_P3_INSTQUEUE_REG_3__4_ & n65316;
  assign n65509 = P2_P3_INSTQUEUE_REG_2__4_ & n65318;
  assign n65510 = P2_P3_INSTQUEUE_REG_1__4_ & n65320;
  assign n65511 = P2_P3_INSTQUEUE_REG_0__4_ & n65322;
  assign n65512 = ~n65508 & ~n65509;
  assign n65513 = ~n65510 & n65512;
  assign n65514 = ~n65511 & n65513;
  assign n65515 = P2_P3_INSTQUEUE_REG_15__4_ & n65328;
  assign n65516 = P2_P3_INSTQUEUE_REG_14__4_ & n65330;
  assign n65517 = P2_P3_INSTQUEUE_REG_13__4_ & n65332;
  assign n65518 = P2_P3_INSTQUEUE_REG_12__4_ & n65334;
  assign n65519 = ~n65515 & ~n65516;
  assign n65520 = ~n65517 & n65519;
  assign n65521 = ~n65518 & n65520;
  assign n65522 = P2_P3_INSTQUEUE_REG_11__4_ & n65340;
  assign n65523 = P2_P3_INSTQUEUE_REG_10__4_ & n65342;
  assign n65524 = P2_P3_INSTQUEUE_REG_9__4_ & n65344;
  assign n65525 = P2_P3_INSTQUEUE_REG_8__4_ & n65346;
  assign n65526 = ~n65522 & ~n65523;
  assign n65527 = ~n65524 & n65526;
  assign n65528 = ~n65525 & n65527;
  assign n65529 = n65507 & n65514;
  assign n65530 = n65521 & n65529;
  assign n65531 = n65528 & n65530;
  assign n65532 = n64842 & ~n65531;
  assign n65533 = ~n65500 & ~n65532;
  assign n65534 = P2_P3_EAX_REG_19_ & n65490;
  assign n65535 = ~P2_P3_EAX_REG_20_ & n65534;
  assign n65536 = P2_P3_EAX_REG_20_ & ~n65534;
  assign n65537 = ~n65535 & ~n65536;
  assign n65538 = n64848 & ~n65537;
  assign n65539 = ~n65498 & ~n65499;
  assign n65540 = n65533 & n65539;
  assign n11776 = n65538 | ~n65540;
  assign n65542 = P2_BUF2_REG_21_ & n65293;
  assign n65543 = P2_BUF2_REG_5_ & n65295;
  assign n65544 = P2_P3_EAX_REG_21_ & ~n64841;
  assign n65545 = P2_P3_INSTQUEUE_REG_7__5_ & n65304;
  assign n65546 = P2_P3_INSTQUEUE_REG_6__5_ & n65306;
  assign n65547 = P2_P3_INSTQUEUE_REG_5__5_ & n65308;
  assign n65548 = P2_P3_INSTQUEUE_REG_4__5_ & n65310;
  assign n65549 = ~n65545 & ~n65546;
  assign n65550 = ~n65547 & n65549;
  assign n65551 = ~n65548 & n65550;
  assign n65552 = P2_P3_INSTQUEUE_REG_3__5_ & n65316;
  assign n65553 = P2_P3_INSTQUEUE_REG_2__5_ & n65318;
  assign n65554 = P2_P3_INSTQUEUE_REG_1__5_ & n65320;
  assign n65555 = P2_P3_INSTQUEUE_REG_0__5_ & n65322;
  assign n65556 = ~n65552 & ~n65553;
  assign n65557 = ~n65554 & n65556;
  assign n65558 = ~n65555 & n65557;
  assign n65559 = P2_P3_INSTQUEUE_REG_15__5_ & n65328;
  assign n65560 = P2_P3_INSTQUEUE_REG_14__5_ & n65330;
  assign n65561 = P2_P3_INSTQUEUE_REG_13__5_ & n65332;
  assign n65562 = P2_P3_INSTQUEUE_REG_12__5_ & n65334;
  assign n65563 = ~n65559 & ~n65560;
  assign n65564 = ~n65561 & n65563;
  assign n65565 = ~n65562 & n65564;
  assign n65566 = P2_P3_INSTQUEUE_REG_11__5_ & n65340;
  assign n65567 = P2_P3_INSTQUEUE_REG_10__5_ & n65342;
  assign n65568 = P2_P3_INSTQUEUE_REG_9__5_ & n65344;
  assign n65569 = P2_P3_INSTQUEUE_REG_8__5_ & n65346;
  assign n65570 = ~n65566 & ~n65567;
  assign n65571 = ~n65568 & n65570;
  assign n65572 = ~n65569 & n65571;
  assign n65573 = n65551 & n65558;
  assign n65574 = n65565 & n65573;
  assign n65575 = n65572 & n65574;
  assign n65576 = n64842 & ~n65575;
  assign n65577 = ~n65544 & ~n65576;
  assign n65578 = P2_P3_EAX_REG_19_ & P2_P3_EAX_REG_20_;
  assign n65579 = n65490 & n65578;
  assign n65580 = P2_P3_EAX_REG_21_ & ~n65579;
  assign n65581 = ~P2_P3_EAX_REG_21_ & n65579;
  assign n65582 = ~n65580 & ~n65581;
  assign n65583 = n64848 & ~n65582;
  assign n65584 = ~n65542 & ~n65543;
  assign n65585 = n65577 & n65584;
  assign n11781 = n65583 | ~n65585;
  assign n65587 = P2_BUF2_REG_22_ & n65293;
  assign n65588 = P2_BUF2_REG_6_ & n65295;
  assign n65589 = P2_P3_EAX_REG_22_ & ~n64841;
  assign n65590 = P2_P3_INSTQUEUE_REG_7__6_ & n65304;
  assign n65591 = P2_P3_INSTQUEUE_REG_6__6_ & n65306;
  assign n65592 = P2_P3_INSTQUEUE_REG_5__6_ & n65308;
  assign n65593 = P2_P3_INSTQUEUE_REG_4__6_ & n65310;
  assign n65594 = ~n65590 & ~n65591;
  assign n65595 = ~n65592 & n65594;
  assign n65596 = ~n65593 & n65595;
  assign n65597 = P2_P3_INSTQUEUE_REG_3__6_ & n65316;
  assign n65598 = P2_P3_INSTQUEUE_REG_2__6_ & n65318;
  assign n65599 = P2_P3_INSTQUEUE_REG_1__6_ & n65320;
  assign n65600 = P2_P3_INSTQUEUE_REG_0__6_ & n65322;
  assign n65601 = ~n65597 & ~n65598;
  assign n65602 = ~n65599 & n65601;
  assign n65603 = ~n65600 & n65602;
  assign n65604 = P2_P3_INSTQUEUE_REG_15__6_ & n65328;
  assign n65605 = P2_P3_INSTQUEUE_REG_14__6_ & n65330;
  assign n65606 = P2_P3_INSTQUEUE_REG_13__6_ & n65332;
  assign n65607 = P2_P3_INSTQUEUE_REG_12__6_ & n65334;
  assign n65608 = ~n65604 & ~n65605;
  assign n65609 = ~n65606 & n65608;
  assign n65610 = ~n65607 & n65609;
  assign n65611 = P2_P3_INSTQUEUE_REG_11__6_ & n65340;
  assign n65612 = P2_P3_INSTQUEUE_REG_10__6_ & n65342;
  assign n65613 = P2_P3_INSTQUEUE_REG_9__6_ & n65344;
  assign n65614 = P2_P3_INSTQUEUE_REG_8__6_ & n65346;
  assign n65615 = ~n65611 & ~n65612;
  assign n65616 = ~n65613 & n65615;
  assign n65617 = ~n65614 & n65616;
  assign n65618 = n65596 & n65603;
  assign n65619 = n65610 & n65618;
  assign n65620 = n65617 & n65619;
  assign n65621 = n64842 & ~n65620;
  assign n65622 = ~n65589 & ~n65621;
  assign n65623 = P2_P3_EAX_REG_21_ & n65579;
  assign n65624 = ~P2_P3_EAX_REG_22_ & n65623;
  assign n65625 = P2_P3_EAX_REG_22_ & ~n65623;
  assign n65626 = ~n65624 & ~n65625;
  assign n65627 = n64848 & ~n65626;
  assign n65628 = ~n65587 & ~n65588;
  assign n65629 = n65622 & n65628;
  assign n11786 = n65627 | ~n65629;
  assign n65631 = P2_BUF2_REG_23_ & n65293;
  assign n65632 = P2_BUF2_REG_7_ & n65295;
  assign n65633 = P2_P3_EAX_REG_23_ & ~n64841;
  assign n65634 = P2_P3_INSTQUEUERD_ADDR_REG_3_ & ~P2_P3_INSTQUEUERD_ADDR_REG_2_;
  assign n65635 = ~n58717 & ~n65634;
  assign n65636 = n58688 & n65635;
  assign n65637 = P2_P3_INSTQUEUE_REG_7__0_ & n65636;
  assign n65638 = n58692 & n65635;
  assign n65639 = P2_P3_INSTQUEUE_REG_6__0_ & n65638;
  assign n65640 = n58697 & n65635;
  assign n65641 = P2_P3_INSTQUEUE_REG_5__0_ & n65640;
  assign n65642 = n58701 & n65635;
  assign n65643 = P2_P3_INSTQUEUE_REG_4__0_ & n65642;
  assign n65644 = ~n65637 & ~n65639;
  assign n65645 = ~n65641 & n65644;
  assign n65646 = ~n65643 & n65645;
  assign n65647 = P2_P3_INSTQUEUERD_ADDR_REG_2_ & n65635;
  assign n65648 = n58687 & n65647;
  assign n65649 = P2_P3_INSTQUEUE_REG_3__0_ & n65648;
  assign n65650 = n58691 & n65647;
  assign n65651 = P2_P3_INSTQUEUE_REG_2__0_ & n65650;
  assign n65652 = n58696 & n65647;
  assign n65653 = P2_P3_INSTQUEUE_REG_1__0_ & n65652;
  assign n65654 = n58700 & n65647;
  assign n65655 = P2_P3_INSTQUEUE_REG_0__0_ & n65654;
  assign n65656 = ~n65649 & ~n65651;
  assign n65657 = ~n65653 & n65656;
  assign n65658 = ~n65655 & n65657;
  assign n65659 = n58688 & ~n65635;
  assign n65660 = P2_P3_INSTQUEUE_REG_15__0_ & n65659;
  assign n65661 = n58692 & ~n65635;
  assign n65662 = P2_P3_INSTQUEUE_REG_14__0_ & n65661;
  assign n65663 = n58697 & ~n65635;
  assign n65664 = P2_P3_INSTQUEUE_REG_13__0_ & n65663;
  assign n65665 = n58701 & ~n65635;
  assign n65666 = P2_P3_INSTQUEUE_REG_12__0_ & n65665;
  assign n65667 = ~n65660 & ~n65662;
  assign n65668 = ~n65664 & n65667;
  assign n65669 = ~n65666 & n65668;
  assign n65670 = P2_P3_INSTQUEUERD_ADDR_REG_2_ & ~n65635;
  assign n65671 = n58687 & n65670;
  assign n65672 = P2_P3_INSTQUEUE_REG_11__0_ & n65671;
  assign n65673 = n58691 & n65670;
  assign n65674 = P2_P3_INSTQUEUE_REG_10__0_ & n65673;
  assign n65675 = n58696 & n65670;
  assign n65676 = P2_P3_INSTQUEUE_REG_9__0_ & n65675;
  assign n65677 = n58700 & n65670;
  assign n65678 = P2_P3_INSTQUEUE_REG_8__0_ & n65677;
  assign n65679 = ~n65672 & ~n65674;
  assign n65680 = ~n65676 & n65679;
  assign n65681 = ~n65678 & n65680;
  assign n65682 = n65646 & n65658;
  assign n65683 = n65669 & n65682;
  assign n65684 = n65681 & n65683;
  assign n65685 = P2_P3_INSTQUEUE_REG_7__7_ & n65304;
  assign n65686 = P2_P3_INSTQUEUE_REG_6__7_ & n65306;
  assign n65687 = P2_P3_INSTQUEUE_REG_5__7_ & n65308;
  assign n65688 = P2_P3_INSTQUEUE_REG_4__7_ & n65310;
  assign n65689 = ~n65685 & ~n65686;
  assign n65690 = ~n65687 & n65689;
  assign n65691 = ~n65688 & n65690;
  assign n65692 = P2_P3_INSTQUEUE_REG_3__7_ & n65316;
  assign n65693 = P2_P3_INSTQUEUE_REG_2__7_ & n65318;
  assign n65694 = P2_P3_INSTQUEUE_REG_1__7_ & n65320;
  assign n65695 = P2_P3_INSTQUEUE_REG_0__7_ & n65322;
  assign n65696 = ~n65692 & ~n65693;
  assign n65697 = ~n65694 & n65696;
  assign n65698 = ~n65695 & n65697;
  assign n65699 = P2_P3_INSTQUEUE_REG_15__7_ & n65328;
  assign n65700 = P2_P3_INSTQUEUE_REG_14__7_ & n65330;
  assign n65701 = P2_P3_INSTQUEUE_REG_13__7_ & n65332;
  assign n65702 = P2_P3_INSTQUEUE_REG_12__7_ & n65334;
  assign n65703 = ~n65699 & ~n65700;
  assign n65704 = ~n65701 & n65703;
  assign n65705 = ~n65702 & n65704;
  assign n65706 = P2_P3_INSTQUEUE_REG_11__7_ & n65340;
  assign n65707 = P2_P3_INSTQUEUE_REG_10__7_ & n65342;
  assign n65708 = P2_P3_INSTQUEUE_REG_9__7_ & n65344;
  assign n65709 = P2_P3_INSTQUEUE_REG_8__7_ & n65346;
  assign n65710 = ~n65706 & ~n65707;
  assign n65711 = ~n65708 & n65710;
  assign n65712 = ~n65709 & n65711;
  assign n65713 = n65691 & n65698;
  assign n65714 = n65705 & n65713;
  assign n65715 = n65712 & n65714;
  assign n65716 = ~n65684 & n65715;
  assign n65717 = n65684 & ~n65715;
  assign n65718 = ~n65716 & ~n65717;
  assign n65719 = n64842 & ~n65718;
  assign n65720 = ~n65633 & ~n65719;
  assign n65721 = P2_P3_EAX_REG_21_ & P2_P3_EAX_REG_22_;
  assign n65722 = n65579 & n65721;
  assign n65723 = P2_P3_EAX_REG_23_ & ~n65722;
  assign n65724 = ~P2_P3_EAX_REG_23_ & n65722;
  assign n65725 = ~n65723 & ~n65724;
  assign n65726 = n64848 & ~n65725;
  assign n65727 = ~n65631 & ~n65632;
  assign n65728 = n65720 & n65727;
  assign n11791 = n65726 | ~n65728;
  assign n65730 = P2_BUF2_REG_24_ & n65293;
  assign n65731 = P2_BUF2_REG_8_ & n65295;
  assign n65732 = P2_P3_EAX_REG_24_ & ~n64841;
  assign n65733 = ~n65684 & ~n65715;
  assign n65734 = P2_P3_INSTQUEUE_REG_7__1_ & n65636;
  assign n65735 = P2_P3_INSTQUEUE_REG_6__1_ & n65638;
  assign n65736 = P2_P3_INSTQUEUE_REG_5__1_ & n65640;
  assign n65737 = P2_P3_INSTQUEUE_REG_4__1_ & n65642;
  assign n65738 = ~n65734 & ~n65735;
  assign n65739 = ~n65736 & n65738;
  assign n65740 = ~n65737 & n65739;
  assign n65741 = P2_P3_INSTQUEUE_REG_3__1_ & n65648;
  assign n65742 = P2_P3_INSTQUEUE_REG_2__1_ & n65650;
  assign n65743 = P2_P3_INSTQUEUE_REG_1__1_ & n65652;
  assign n65744 = P2_P3_INSTQUEUE_REG_0__1_ & n65654;
  assign n65745 = ~n65741 & ~n65742;
  assign n65746 = ~n65743 & n65745;
  assign n65747 = ~n65744 & n65746;
  assign n65748 = P2_P3_INSTQUEUE_REG_15__1_ & n65659;
  assign n65749 = P2_P3_INSTQUEUE_REG_14__1_ & n65661;
  assign n65750 = P2_P3_INSTQUEUE_REG_13__1_ & n65663;
  assign n65751 = P2_P3_INSTQUEUE_REG_12__1_ & n65665;
  assign n65752 = ~n65748 & ~n65749;
  assign n65753 = ~n65750 & n65752;
  assign n65754 = ~n65751 & n65753;
  assign n65755 = P2_P3_INSTQUEUE_REG_11__1_ & n65671;
  assign n65756 = P2_P3_INSTQUEUE_REG_10__1_ & n65673;
  assign n65757 = P2_P3_INSTQUEUE_REG_9__1_ & n65675;
  assign n65758 = P2_P3_INSTQUEUE_REG_8__1_ & n65677;
  assign n65759 = ~n65755 & ~n65756;
  assign n65760 = ~n65757 & n65759;
  assign n65761 = ~n65758 & n65760;
  assign n65762 = n65740 & n65747;
  assign n65763 = n65754 & n65762;
  assign n65764 = n65761 & n65763;
  assign n65765 = n65733 & n65764;
  assign n65766 = ~n65733 & ~n65764;
  assign n65767 = ~n65765 & ~n65766;
  assign n65768 = n64842 & ~n65767;
  assign n65769 = ~n65732 & ~n65768;
  assign n65770 = P2_P3_EAX_REG_23_ & n65722;
  assign n65771 = ~P2_P3_EAX_REG_24_ & n65770;
  assign n65772 = P2_P3_EAX_REG_24_ & ~n65770;
  assign n65773 = ~n65771 & ~n65772;
  assign n65774 = n64848 & ~n65773;
  assign n65775 = ~n65730 & ~n65731;
  assign n65776 = n65769 & n65775;
  assign n11796 = n65774 | ~n65776;
  assign n65778 = P2_BUF2_REG_25_ & n65293;
  assign n65779 = P2_BUF2_REG_9_ & n65295;
  assign n65780 = P2_P3_EAX_REG_25_ & ~n64841;
  assign n65781 = n65733 & ~n65764;
  assign n65782 = P2_P3_INSTQUEUE_REG_7__2_ & n65636;
  assign n65783 = P2_P3_INSTQUEUE_REG_6__2_ & n65638;
  assign n65784 = P2_P3_INSTQUEUE_REG_5__2_ & n65640;
  assign n65785 = P2_P3_INSTQUEUE_REG_4__2_ & n65642;
  assign n65786 = ~n65782 & ~n65783;
  assign n65787 = ~n65784 & n65786;
  assign n65788 = ~n65785 & n65787;
  assign n65789 = P2_P3_INSTQUEUE_REG_3__2_ & n65648;
  assign n65790 = P2_P3_INSTQUEUE_REG_2__2_ & n65650;
  assign n65791 = P2_P3_INSTQUEUE_REG_1__2_ & n65652;
  assign n65792 = P2_P3_INSTQUEUE_REG_0__2_ & n65654;
  assign n65793 = ~n65789 & ~n65790;
  assign n65794 = ~n65791 & n65793;
  assign n65795 = ~n65792 & n65794;
  assign n65796 = P2_P3_INSTQUEUE_REG_15__2_ & n65659;
  assign n65797 = P2_P3_INSTQUEUE_REG_14__2_ & n65661;
  assign n65798 = P2_P3_INSTQUEUE_REG_13__2_ & n65663;
  assign n65799 = P2_P3_INSTQUEUE_REG_12__2_ & n65665;
  assign n65800 = ~n65796 & ~n65797;
  assign n65801 = ~n65798 & n65800;
  assign n65802 = ~n65799 & n65801;
  assign n65803 = P2_P3_INSTQUEUE_REG_11__2_ & n65671;
  assign n65804 = P2_P3_INSTQUEUE_REG_10__2_ & n65673;
  assign n65805 = P2_P3_INSTQUEUE_REG_9__2_ & n65675;
  assign n65806 = P2_P3_INSTQUEUE_REG_8__2_ & n65677;
  assign n65807 = ~n65803 & ~n65804;
  assign n65808 = ~n65805 & n65807;
  assign n65809 = ~n65806 & n65808;
  assign n65810 = n65788 & n65795;
  assign n65811 = n65802 & n65810;
  assign n65812 = n65809 & n65811;
  assign n65813 = n65781 & n65812;
  assign n65814 = ~n65781 & ~n65812;
  assign n65815 = ~n65813 & ~n65814;
  assign n65816 = n64842 & ~n65815;
  assign n65817 = ~n65780 & ~n65816;
  assign n65818 = P2_P3_EAX_REG_23_ & P2_P3_EAX_REG_24_;
  assign n65819 = n65722 & n65818;
  assign n65820 = P2_P3_EAX_REG_25_ & ~n65819;
  assign n65821 = ~P2_P3_EAX_REG_25_ & n65819;
  assign n65822 = ~n65820 & ~n65821;
  assign n65823 = n64848 & ~n65822;
  assign n65824 = ~n65778 & ~n65779;
  assign n65825 = n65817 & n65824;
  assign n11801 = n65823 | ~n65825;
  assign n65827 = P2_BUF2_REG_26_ & n65293;
  assign n65828 = P2_BUF2_REG_10_ & n65295;
  assign n65829 = P2_P3_EAX_REG_26_ & ~n64841;
  assign n65830 = n65781 & ~n65812;
  assign n65831 = P2_P3_INSTQUEUE_REG_7__3_ & n65636;
  assign n65832 = P2_P3_INSTQUEUE_REG_6__3_ & n65638;
  assign n65833 = P2_P3_INSTQUEUE_REG_5__3_ & n65640;
  assign n65834 = P2_P3_INSTQUEUE_REG_4__3_ & n65642;
  assign n65835 = ~n65831 & ~n65832;
  assign n65836 = ~n65833 & n65835;
  assign n65837 = ~n65834 & n65836;
  assign n65838 = P2_P3_INSTQUEUE_REG_3__3_ & n65648;
  assign n65839 = P2_P3_INSTQUEUE_REG_2__3_ & n65650;
  assign n65840 = P2_P3_INSTQUEUE_REG_1__3_ & n65652;
  assign n65841 = P2_P3_INSTQUEUE_REG_0__3_ & n65654;
  assign n65842 = ~n65838 & ~n65839;
  assign n65843 = ~n65840 & n65842;
  assign n65844 = ~n65841 & n65843;
  assign n65845 = P2_P3_INSTQUEUE_REG_15__3_ & n65659;
  assign n65846 = P2_P3_INSTQUEUE_REG_14__3_ & n65661;
  assign n65847 = P2_P3_INSTQUEUE_REG_13__3_ & n65663;
  assign n65848 = P2_P3_INSTQUEUE_REG_12__3_ & n65665;
  assign n65849 = ~n65845 & ~n65846;
  assign n65850 = ~n65847 & n65849;
  assign n65851 = ~n65848 & n65850;
  assign n65852 = P2_P3_INSTQUEUE_REG_11__3_ & n65671;
  assign n65853 = P2_P3_INSTQUEUE_REG_10__3_ & n65673;
  assign n65854 = P2_P3_INSTQUEUE_REG_9__3_ & n65675;
  assign n65855 = P2_P3_INSTQUEUE_REG_8__3_ & n65677;
  assign n65856 = ~n65852 & ~n65853;
  assign n65857 = ~n65854 & n65856;
  assign n65858 = ~n65855 & n65857;
  assign n65859 = n65837 & n65844;
  assign n65860 = n65851 & n65859;
  assign n65861 = n65858 & n65860;
  assign n65862 = n65830 & n65861;
  assign n65863 = ~n65830 & ~n65861;
  assign n65864 = ~n65862 & ~n65863;
  assign n65865 = n64842 & ~n65864;
  assign n65866 = ~n65829 & ~n65865;
  assign n65867 = P2_P3_EAX_REG_25_ & n65819;
  assign n65868 = ~P2_P3_EAX_REG_26_ & n65867;
  assign n65869 = P2_P3_EAX_REG_26_ & ~n65867;
  assign n65870 = ~n65868 & ~n65869;
  assign n65871 = n64848 & ~n65870;
  assign n65872 = ~n65827 & ~n65828;
  assign n65873 = n65866 & n65872;
  assign n11806 = n65871 | ~n65873;
  assign n65875 = P2_BUF2_REG_27_ & n65293;
  assign n65876 = P2_BUF2_REG_11_ & n65295;
  assign n65877 = P2_P3_EAX_REG_27_ & ~n64841;
  assign n65878 = n65830 & ~n65861;
  assign n65879 = P2_P3_INSTQUEUE_REG_7__4_ & n65636;
  assign n65880 = P2_P3_INSTQUEUE_REG_6__4_ & n65638;
  assign n65881 = P2_P3_INSTQUEUE_REG_5__4_ & n65640;
  assign n65882 = P2_P3_INSTQUEUE_REG_4__4_ & n65642;
  assign n65883 = ~n65879 & ~n65880;
  assign n65884 = ~n65881 & n65883;
  assign n65885 = ~n65882 & n65884;
  assign n65886 = P2_P3_INSTQUEUE_REG_3__4_ & n65648;
  assign n65887 = P2_P3_INSTQUEUE_REG_2__4_ & n65650;
  assign n65888 = P2_P3_INSTQUEUE_REG_1__4_ & n65652;
  assign n65889 = P2_P3_INSTQUEUE_REG_0__4_ & n65654;
  assign n65890 = ~n65886 & ~n65887;
  assign n65891 = ~n65888 & n65890;
  assign n65892 = ~n65889 & n65891;
  assign n65893 = P2_P3_INSTQUEUE_REG_15__4_ & n65659;
  assign n65894 = P2_P3_INSTQUEUE_REG_14__4_ & n65661;
  assign n65895 = P2_P3_INSTQUEUE_REG_13__4_ & n65663;
  assign n65896 = P2_P3_INSTQUEUE_REG_12__4_ & n65665;
  assign n65897 = ~n65893 & ~n65894;
  assign n65898 = ~n65895 & n65897;
  assign n65899 = ~n65896 & n65898;
  assign n65900 = P2_P3_INSTQUEUE_REG_11__4_ & n65671;
  assign n65901 = P2_P3_INSTQUEUE_REG_10__4_ & n65673;
  assign n65902 = P2_P3_INSTQUEUE_REG_9__4_ & n65675;
  assign n65903 = P2_P3_INSTQUEUE_REG_8__4_ & n65677;
  assign n65904 = ~n65900 & ~n65901;
  assign n65905 = ~n65902 & n65904;
  assign n65906 = ~n65903 & n65905;
  assign n65907 = n65885 & n65892;
  assign n65908 = n65899 & n65907;
  assign n65909 = n65906 & n65908;
  assign n65910 = n65878 & n65909;
  assign n65911 = ~n65878 & ~n65909;
  assign n65912 = ~n65910 & ~n65911;
  assign n65913 = n64842 & ~n65912;
  assign n65914 = ~n65877 & ~n65913;
  assign n65915 = P2_P3_EAX_REG_25_ & P2_P3_EAX_REG_26_;
  assign n65916 = n65819 & n65915;
  assign n65917 = P2_P3_EAX_REG_27_ & ~n65916;
  assign n65918 = ~P2_P3_EAX_REG_27_ & n65916;
  assign n65919 = ~n65917 & ~n65918;
  assign n65920 = n64848 & ~n65919;
  assign n65921 = ~n65875 & ~n65876;
  assign n65922 = n65914 & n65921;
  assign n11811 = n65920 | ~n65922;
  assign n65924 = P2_BUF2_REG_28_ & n65293;
  assign n65925 = P2_BUF2_REG_12_ & n65295;
  assign n65926 = P2_P3_EAX_REG_28_ & ~n64841;
  assign n65927 = n65878 & ~n65909;
  assign n65928 = P2_P3_INSTQUEUE_REG_7__5_ & n65636;
  assign n65929 = P2_P3_INSTQUEUE_REG_6__5_ & n65638;
  assign n65930 = P2_P3_INSTQUEUE_REG_5__5_ & n65640;
  assign n65931 = P2_P3_INSTQUEUE_REG_4__5_ & n65642;
  assign n65932 = ~n65928 & ~n65929;
  assign n65933 = ~n65930 & n65932;
  assign n65934 = ~n65931 & n65933;
  assign n65935 = P2_P3_INSTQUEUE_REG_3__5_ & n65648;
  assign n65936 = P2_P3_INSTQUEUE_REG_2__5_ & n65650;
  assign n65937 = P2_P3_INSTQUEUE_REG_1__5_ & n65652;
  assign n65938 = P2_P3_INSTQUEUE_REG_0__5_ & n65654;
  assign n65939 = ~n65935 & ~n65936;
  assign n65940 = ~n65937 & n65939;
  assign n65941 = ~n65938 & n65940;
  assign n65942 = P2_P3_INSTQUEUE_REG_15__5_ & n65659;
  assign n65943 = P2_P3_INSTQUEUE_REG_14__5_ & n65661;
  assign n65944 = P2_P3_INSTQUEUE_REG_13__5_ & n65663;
  assign n65945 = P2_P3_INSTQUEUE_REG_12__5_ & n65665;
  assign n65946 = ~n65942 & ~n65943;
  assign n65947 = ~n65944 & n65946;
  assign n65948 = ~n65945 & n65947;
  assign n65949 = P2_P3_INSTQUEUE_REG_11__5_ & n65671;
  assign n65950 = P2_P3_INSTQUEUE_REG_10__5_ & n65673;
  assign n65951 = P2_P3_INSTQUEUE_REG_9__5_ & n65675;
  assign n65952 = P2_P3_INSTQUEUE_REG_8__5_ & n65677;
  assign n65953 = ~n65949 & ~n65950;
  assign n65954 = ~n65951 & n65953;
  assign n65955 = ~n65952 & n65954;
  assign n65956 = n65934 & n65941;
  assign n65957 = n65948 & n65956;
  assign n65958 = n65955 & n65957;
  assign n65959 = n65927 & n65958;
  assign n65960 = ~n65927 & ~n65958;
  assign n65961 = ~n65959 & ~n65960;
  assign n65962 = n64842 & ~n65961;
  assign n65963 = P2_P3_EAX_REG_27_ & n65916;
  assign n65964 = ~P2_P3_EAX_REG_28_ & n65963;
  assign n65965 = P2_P3_EAX_REG_28_ & ~n65963;
  assign n65966 = ~n65964 & ~n65965;
  assign n65967 = n64848 & ~n65966;
  assign n65968 = ~n65924 & ~n65925;
  assign n65969 = ~n65926 & n65968;
  assign n65970 = ~n65962 & n65969;
  assign n11816 = n65967 | ~n65970;
  assign n65972 = P2_BUF2_REG_29_ & n65293;
  assign n65973 = P2_BUF2_REG_13_ & n65295;
  assign n65974 = P2_P3_EAX_REG_29_ & ~n64841;
  assign n65975 = n65927 & ~n65958;
  assign n65976 = P2_P3_INSTQUEUE_REG_7__6_ & n65636;
  assign n65977 = P2_P3_INSTQUEUE_REG_6__6_ & n65638;
  assign n65978 = P2_P3_INSTQUEUE_REG_5__6_ & n65640;
  assign n65979 = P2_P3_INSTQUEUE_REG_4__6_ & n65642;
  assign n65980 = ~n65976 & ~n65977;
  assign n65981 = ~n65978 & n65980;
  assign n65982 = ~n65979 & n65981;
  assign n65983 = P2_P3_INSTQUEUE_REG_3__6_ & n65648;
  assign n65984 = P2_P3_INSTQUEUE_REG_2__6_ & n65650;
  assign n65985 = P2_P3_INSTQUEUE_REG_1__6_ & n65652;
  assign n65986 = P2_P3_INSTQUEUE_REG_0__6_ & n65654;
  assign n65987 = ~n65983 & ~n65984;
  assign n65988 = ~n65985 & n65987;
  assign n65989 = ~n65986 & n65988;
  assign n65990 = P2_P3_INSTQUEUE_REG_15__6_ & n65659;
  assign n65991 = P2_P3_INSTQUEUE_REG_14__6_ & n65661;
  assign n65992 = P2_P3_INSTQUEUE_REG_13__6_ & n65663;
  assign n65993 = P2_P3_INSTQUEUE_REG_12__6_ & n65665;
  assign n65994 = ~n65990 & ~n65991;
  assign n65995 = ~n65992 & n65994;
  assign n65996 = ~n65993 & n65995;
  assign n65997 = P2_P3_INSTQUEUE_REG_11__6_ & n65671;
  assign n65998 = P2_P3_INSTQUEUE_REG_10__6_ & n65673;
  assign n65999 = P2_P3_INSTQUEUE_REG_9__6_ & n65675;
  assign n66000 = P2_P3_INSTQUEUE_REG_8__6_ & n65677;
  assign n66001 = ~n65997 & ~n65998;
  assign n66002 = ~n65999 & n66001;
  assign n66003 = ~n66000 & n66002;
  assign n66004 = n65982 & n65989;
  assign n66005 = n65996 & n66004;
  assign n66006 = n66003 & n66005;
  assign n66007 = n65975 & n66006;
  assign n66008 = ~n65975 & ~n66006;
  assign n66009 = ~n66007 & ~n66008;
  assign n66010 = n64842 & ~n66009;
  assign n66011 = P2_P3_EAX_REG_27_ & P2_P3_EAX_REG_28_;
  assign n66012 = n65916 & n66011;
  assign n66013 = P2_P3_EAX_REG_29_ & ~n66012;
  assign n66014 = ~P2_P3_EAX_REG_29_ & n66012;
  assign n66015 = ~n66013 & ~n66014;
  assign n66016 = n64848 & ~n66015;
  assign n66017 = ~n65972 & ~n65973;
  assign n66018 = ~n65974 & n66017;
  assign n66019 = ~n66010 & n66018;
  assign n11821 = n66016 | ~n66019;
  assign n66021 = P2_BUF2_REG_30_ & n65293;
  assign n66022 = P2_BUF2_REG_14_ & n65295;
  assign n66023 = P2_P3_EAX_REG_30_ & ~n64841;
  assign n66024 = n65975 & ~n66006;
  assign n66025 = P2_P3_INSTQUEUE_REG_7__7_ & n65636;
  assign n66026 = P2_P3_INSTQUEUE_REG_6__7_ & n65638;
  assign n66027 = P2_P3_INSTQUEUE_REG_5__7_ & n65640;
  assign n66028 = P2_P3_INSTQUEUE_REG_4__7_ & n65642;
  assign n66029 = ~n66025 & ~n66026;
  assign n66030 = ~n66027 & n66029;
  assign n66031 = ~n66028 & n66030;
  assign n66032 = P2_P3_INSTQUEUE_REG_3__7_ & n65648;
  assign n66033 = P2_P3_INSTQUEUE_REG_2__7_ & n65650;
  assign n66034 = P2_P3_INSTQUEUE_REG_1__7_ & n65652;
  assign n66035 = P2_P3_INSTQUEUE_REG_0__7_ & n65654;
  assign n66036 = ~n66032 & ~n66033;
  assign n66037 = ~n66034 & n66036;
  assign n66038 = ~n66035 & n66037;
  assign n66039 = P2_P3_INSTQUEUE_REG_15__7_ & n65659;
  assign n66040 = P2_P3_INSTQUEUE_REG_14__7_ & n65661;
  assign n66041 = P2_P3_INSTQUEUE_REG_13__7_ & n65663;
  assign n66042 = P2_P3_INSTQUEUE_REG_12__7_ & n65665;
  assign n66043 = ~n66039 & ~n66040;
  assign n66044 = ~n66041 & n66043;
  assign n66045 = ~n66042 & n66044;
  assign n66046 = P2_P3_INSTQUEUE_REG_11__7_ & n65671;
  assign n66047 = P2_P3_INSTQUEUE_REG_10__7_ & n65673;
  assign n66048 = P2_P3_INSTQUEUE_REG_9__7_ & n65675;
  assign n66049 = P2_P3_INSTQUEUE_REG_8__7_ & n65677;
  assign n66050 = ~n66046 & ~n66047;
  assign n66051 = ~n66048 & n66050;
  assign n66052 = ~n66049 & n66051;
  assign n66053 = n66031 & n66038;
  assign n66054 = n66045 & n66053;
  assign n66055 = n66052 & n66054;
  assign n66056 = n66024 & n66055;
  assign n66057 = ~n66024 & ~n66055;
  assign n66058 = ~n66056 & ~n66057;
  assign n66059 = n64842 & ~n66058;
  assign n66060 = P2_P3_EAX_REG_29_ & n66012;
  assign n66061 = ~P2_P3_EAX_REG_30_ & n66060;
  assign n66062 = P2_P3_EAX_REG_30_ & ~n66060;
  assign n66063 = ~n66061 & ~n66062;
  assign n66064 = n64848 & ~n66063;
  assign n66065 = ~n66021 & ~n66022;
  assign n66066 = ~n66023 & n66065;
  assign n66067 = ~n66059 & n66066;
  assign n11826 = n66064 | ~n66067;
  assign n66069 = P2_P3_EAX_REG_31_ & ~n64841;
  assign n66070 = P2_BUF2_REG_31_ & n65293;
  assign n66071 = P2_P3_EAX_REG_30_ & n66060;
  assign n66072 = ~P2_P3_EAX_REG_31_ & n66071;
  assign n66073 = P2_P3_EAX_REG_31_ & ~n66071;
  assign n66074 = ~n66072 & ~n66073;
  assign n66075 = n64848 & ~n66074;
  assign n66076 = ~n66069 & ~n66070;
  assign n11831 = n66075 | ~n66076;
  assign n66078 = ~n59108 & ~n59202;
  assign n66079 = n59321 & ~n66078;
  assign n66080 = n58838 & n66079;
  assign n66081 = ~P2_P3_EBX_REG_0_ & n66080;
  assign n66082 = ~n58838 & n66079;
  assign n66083 = P2_P3_INSTQUEUE_REG_0__0_ & n66082;
  assign n66084 = P2_P3_EBX_REG_0_ & ~n66079;
  assign n66085 = ~n66081 & ~n66083;
  assign n11836 = n66084 | ~n66085;
  assign n66087 = ~P2_P3_EBX_REG_0_ & P2_P3_EBX_REG_1_;
  assign n66088 = P2_P3_EBX_REG_0_ & ~P2_P3_EBX_REG_1_;
  assign n66089 = ~n66087 & ~n66088;
  assign n66090 = n66080 & ~n66089;
  assign n66091 = P2_P3_INSTQUEUE_REG_0__1_ & n66082;
  assign n66092 = P2_P3_EBX_REG_1_ & ~n66079;
  assign n66093 = ~n66090 & ~n66091;
  assign n11841 = n66092 | ~n66093;
  assign n66095 = P2_P3_EBX_REG_0_ & P2_P3_EBX_REG_1_;
  assign n66096 = ~P2_P3_EBX_REG_2_ & n66095;
  assign n66097 = P2_P3_EBX_REG_2_ & ~n66095;
  assign n66098 = ~n66096 & ~n66097;
  assign n66099 = n66080 & ~n66098;
  assign n66100 = P2_P3_INSTQUEUE_REG_0__2_ & n66082;
  assign n66101 = P2_P3_EBX_REG_2_ & ~n66079;
  assign n66102 = ~n66099 & ~n66100;
  assign n11846 = n66101 | ~n66102;
  assign n66104 = P2_P3_EBX_REG_0_ & P2_P3_EBX_REG_2_;
  assign n66105 = P2_P3_EBX_REG_1_ & n66104;
  assign n66106 = P2_P3_EBX_REG_3_ & ~n66105;
  assign n66107 = ~P2_P3_EBX_REG_3_ & n66105;
  assign n66108 = ~n66106 & ~n66107;
  assign n66109 = n66080 & ~n66108;
  assign n66110 = P2_P3_INSTQUEUE_REG_0__3_ & n66082;
  assign n66111 = P2_P3_EBX_REG_3_ & ~n66079;
  assign n66112 = ~n66109 & ~n66110;
  assign n11851 = n66111 | ~n66112;
  assign n66114 = P2_P3_EBX_REG_3_ & n66105;
  assign n66115 = ~P2_P3_EBX_REG_4_ & n66114;
  assign n66116 = P2_P3_EBX_REG_4_ & ~n66114;
  assign n66117 = ~n66115 & ~n66116;
  assign n66118 = n66080 & ~n66117;
  assign n66119 = P2_P3_INSTQUEUE_REG_0__4_ & n66082;
  assign n66120 = P2_P3_EBX_REG_4_ & ~n66079;
  assign n66121 = ~n66118 & ~n66119;
  assign n11856 = n66120 | ~n66121;
  assign n66123 = P2_P3_EBX_REG_3_ & P2_P3_EBX_REG_4_;
  assign n66124 = n66105 & n66123;
  assign n66125 = P2_P3_EBX_REG_5_ & ~n66124;
  assign n66126 = ~P2_P3_EBX_REG_5_ & n66124;
  assign n66127 = ~n66125 & ~n66126;
  assign n66128 = n66080 & ~n66127;
  assign n66129 = P2_P3_INSTQUEUE_REG_0__5_ & n66082;
  assign n66130 = P2_P3_EBX_REG_5_ & ~n66079;
  assign n66131 = ~n66128 & ~n66129;
  assign n11861 = n66130 | ~n66131;
  assign n66133 = P2_P3_EBX_REG_5_ & n66124;
  assign n66134 = ~P2_P3_EBX_REG_6_ & n66133;
  assign n66135 = P2_P3_EBX_REG_6_ & ~n66133;
  assign n66136 = ~n66134 & ~n66135;
  assign n66137 = n66080 & ~n66136;
  assign n66138 = P2_P3_INSTQUEUE_REG_0__6_ & n66082;
  assign n66139 = P2_P3_EBX_REG_6_ & ~n66079;
  assign n66140 = ~n66137 & ~n66138;
  assign n11866 = n66139 | ~n66140;
  assign n66142 = P2_P3_EBX_REG_5_ & P2_P3_EBX_REG_6_;
  assign n66143 = n66124 & n66142;
  assign n66144 = P2_P3_EBX_REG_7_ & ~n66143;
  assign n66145 = ~P2_P3_EBX_REG_7_ & n66143;
  assign n66146 = ~n66144 & ~n66145;
  assign n66147 = n66080 & ~n66146;
  assign n66148 = P2_P3_INSTQUEUE_REG_0__7_ & n66082;
  assign n66149 = P2_P3_EBX_REG_7_ & ~n66079;
  assign n66150 = ~n66147 & ~n66148;
  assign n11871 = n66149 | ~n66150;
  assign n66152 = P2_P3_EBX_REG_7_ & n66143;
  assign n66153 = ~P2_P3_EBX_REG_8_ & n66152;
  assign n66154 = P2_P3_EBX_REG_8_ & ~n66152;
  assign n66155 = ~n66153 & ~n66154;
  assign n66156 = n66080 & ~n66155;
  assign n66157 = ~n64983 & n66082;
  assign n66158 = P2_P3_EBX_REG_8_ & ~n66079;
  assign n66159 = ~n66156 & ~n66157;
  assign n11876 = n66158 | ~n66159;
  assign n66161 = P2_P3_EBX_REG_7_ & P2_P3_EBX_REG_8_;
  assign n66162 = n66143 & n66161;
  assign n66163 = P2_P3_EBX_REG_9_ & ~n66162;
  assign n66164 = ~P2_P3_EBX_REG_9_ & n66162;
  assign n66165 = ~n66163 & ~n66164;
  assign n66166 = n66080 & ~n66165;
  assign n66167 = ~n65025 & n66082;
  assign n66168 = P2_P3_EBX_REG_9_ & ~n66079;
  assign n66169 = ~n66166 & ~n66167;
  assign n11881 = n66168 | ~n66169;
  assign n66171 = P2_P3_EBX_REG_10_ & ~n66079;
  assign n66172 = ~n65068 & n66082;
  assign n66173 = P2_P3_EBX_REG_9_ & n66162;
  assign n66174 = ~P2_P3_EBX_REG_10_ & n66173;
  assign n66175 = P2_P3_EBX_REG_10_ & ~n66173;
  assign n66176 = ~n66174 & ~n66175;
  assign n66177 = n66080 & ~n66176;
  assign n66178 = ~n66171 & ~n66172;
  assign n11886 = n66177 | ~n66178;
  assign n66180 = P2_P3_EBX_REG_11_ & ~n66079;
  assign n66181 = ~n65110 & n66082;
  assign n66182 = P2_P3_EBX_REG_9_ & P2_P3_EBX_REG_10_;
  assign n66183 = n66162 & n66182;
  assign n66184 = P2_P3_EBX_REG_11_ & ~n66183;
  assign n66185 = ~P2_P3_EBX_REG_11_ & n66183;
  assign n66186 = ~n66184 & ~n66185;
  assign n66187 = n66080 & ~n66186;
  assign n66188 = ~n66180 & ~n66181;
  assign n11891 = n66187 | ~n66188;
  assign n66190 = P2_P3_EBX_REG_12_ & ~n66079;
  assign n66191 = ~n65153 & n66082;
  assign n66192 = P2_P3_EBX_REG_11_ & n66183;
  assign n66193 = ~P2_P3_EBX_REG_12_ & n66192;
  assign n66194 = P2_P3_EBX_REG_12_ & ~n66192;
  assign n66195 = ~n66193 & ~n66194;
  assign n66196 = n66080 & ~n66195;
  assign n66197 = ~n66190 & ~n66191;
  assign n11896 = n66196 | ~n66197;
  assign n66199 = P2_P3_EBX_REG_13_ & ~n66079;
  assign n66200 = ~n65196 & n66082;
  assign n66201 = P2_P3_EBX_REG_11_ & P2_P3_EBX_REG_12_;
  assign n66202 = n66183 & n66201;
  assign n66203 = P2_P3_EBX_REG_13_ & ~n66202;
  assign n66204 = ~P2_P3_EBX_REG_13_ & n66202;
  assign n66205 = ~n66203 & ~n66204;
  assign n66206 = n66080 & ~n66205;
  assign n66207 = ~n66199 & ~n66200;
  assign n11901 = n66206 | ~n66207;
  assign n66209 = P2_P3_EBX_REG_14_ & ~n66079;
  assign n66210 = ~n65239 & n66082;
  assign n66211 = P2_P3_EBX_REG_13_ & n66202;
  assign n66212 = ~P2_P3_EBX_REG_14_ & n66211;
  assign n66213 = P2_P3_EBX_REG_14_ & ~n66211;
  assign n66214 = ~n66212 & ~n66213;
  assign n66215 = n66080 & ~n66214;
  assign n66216 = ~n66209 & ~n66210;
  assign n11906 = n66215 | ~n66216;
  assign n66218 = P2_P3_EBX_REG_15_ & ~n66079;
  assign n66219 = ~n65281 & n66082;
  assign n66220 = P2_P3_EBX_REG_13_ & P2_P3_EBX_REG_14_;
  assign n66221 = n66202 & n66220;
  assign n66222 = P2_P3_EBX_REG_15_ & ~n66221;
  assign n66223 = ~P2_P3_EBX_REG_15_ & n66221;
  assign n66224 = ~n66222 & ~n66223;
  assign n66225 = n66080 & ~n66224;
  assign n66226 = ~n66218 & ~n66219;
  assign n11911 = n66225 | ~n66226;
  assign n66228 = P2_P3_EBX_REG_16_ & ~n66079;
  assign n66229 = ~n65353 & n66082;
  assign n66230 = P2_P3_EBX_REG_15_ & n66221;
  assign n66231 = ~P2_P3_EBX_REG_16_ & n66230;
  assign n66232 = P2_P3_EBX_REG_16_ & ~n66230;
  assign n66233 = ~n66231 & ~n66232;
  assign n66234 = n66080 & ~n66233;
  assign n66235 = ~n66228 & ~n66229;
  assign n11916 = n66234 | ~n66235;
  assign n66237 = P2_P3_EBX_REG_17_ & ~n66079;
  assign n66238 = ~n65397 & n66082;
  assign n66239 = P2_P3_EBX_REG_15_ & P2_P3_EBX_REG_16_;
  assign n66240 = n66221 & n66239;
  assign n66241 = P2_P3_EBX_REG_17_ & ~n66240;
  assign n66242 = ~P2_P3_EBX_REG_17_ & n66240;
  assign n66243 = ~n66241 & ~n66242;
  assign n66244 = n66080 & ~n66243;
  assign n66245 = ~n66237 & ~n66238;
  assign n11921 = n66244 | ~n66245;
  assign n66247 = P2_P3_EBX_REG_18_ & ~n66079;
  assign n66248 = ~n65442 & n66082;
  assign n66249 = P2_P3_EBX_REG_17_ & n66240;
  assign n66250 = ~P2_P3_EBX_REG_18_ & n66249;
  assign n66251 = P2_P3_EBX_REG_18_ & ~n66249;
  assign n66252 = ~n66250 & ~n66251;
  assign n66253 = n66080 & ~n66252;
  assign n66254 = ~n66247 & ~n66248;
  assign n11926 = n66253 | ~n66254;
  assign n66256 = P2_P3_EBX_REG_19_ & ~n66079;
  assign n66257 = ~n65486 & n66082;
  assign n66258 = P2_P3_EBX_REG_17_ & P2_P3_EBX_REG_18_;
  assign n66259 = n66240 & n66258;
  assign n66260 = P2_P3_EBX_REG_19_ & ~n66259;
  assign n66261 = ~P2_P3_EBX_REG_19_ & n66259;
  assign n66262 = ~n66260 & ~n66261;
  assign n66263 = n66080 & ~n66262;
  assign n66264 = ~n66256 & ~n66257;
  assign n11931 = n66263 | ~n66264;
  assign n66266 = P2_P3_EBX_REG_20_ & ~n66079;
  assign n66267 = ~n65531 & n66082;
  assign n66268 = P2_P3_EBX_REG_19_ & n66259;
  assign n66269 = ~P2_P3_EBX_REG_20_ & n66268;
  assign n66270 = P2_P3_EBX_REG_20_ & ~n66268;
  assign n66271 = ~n66269 & ~n66270;
  assign n66272 = n66080 & ~n66271;
  assign n66273 = ~n66266 & ~n66267;
  assign n11936 = n66272 | ~n66273;
  assign n66275 = P2_P3_EBX_REG_21_ & ~n66079;
  assign n66276 = ~n65575 & n66082;
  assign n66277 = P2_P3_EBX_REG_19_ & P2_P3_EBX_REG_20_;
  assign n66278 = n66259 & n66277;
  assign n66279 = P2_P3_EBX_REG_21_ & ~n66278;
  assign n66280 = ~P2_P3_EBX_REG_21_ & n66278;
  assign n66281 = ~n66279 & ~n66280;
  assign n66282 = n66080 & ~n66281;
  assign n66283 = ~n66275 & ~n66276;
  assign n11941 = n66282 | ~n66283;
  assign n66285 = P2_P3_EBX_REG_22_ & ~n66079;
  assign n66286 = ~n65620 & n66082;
  assign n66287 = P2_P3_EBX_REG_21_ & n66278;
  assign n66288 = ~P2_P3_EBX_REG_22_ & n66287;
  assign n66289 = P2_P3_EBX_REG_22_ & ~n66287;
  assign n66290 = ~n66288 & ~n66289;
  assign n66291 = n66080 & ~n66290;
  assign n66292 = ~n66285 & ~n66286;
  assign n11946 = n66291 | ~n66292;
  assign n66294 = P2_P3_EBX_REG_23_ & ~n66079;
  assign n66295 = ~n65718 & n66082;
  assign n66296 = P2_P3_EBX_REG_21_ & P2_P3_EBX_REG_22_;
  assign n66297 = n66278 & n66296;
  assign n66298 = P2_P3_EBX_REG_23_ & ~n66297;
  assign n66299 = ~P2_P3_EBX_REG_23_ & n66297;
  assign n66300 = ~n66298 & ~n66299;
  assign n66301 = n66080 & ~n66300;
  assign n66302 = ~n66294 & ~n66295;
  assign n11951 = n66301 | ~n66302;
  assign n66304 = P2_P3_EBX_REG_24_ & ~n66079;
  assign n66305 = ~n65767 & n66082;
  assign n66306 = P2_P3_EBX_REG_23_ & n66297;
  assign n66307 = ~P2_P3_EBX_REG_24_ & n66306;
  assign n66308 = P2_P3_EBX_REG_24_ & ~n66306;
  assign n66309 = ~n66307 & ~n66308;
  assign n66310 = n66080 & ~n66309;
  assign n66311 = ~n66304 & ~n66305;
  assign n11956 = n66310 | ~n66311;
  assign n66313 = P2_P3_EBX_REG_25_ & ~n66079;
  assign n66314 = ~n65815 & n66082;
  assign n66315 = P2_P3_EBX_REG_23_ & P2_P3_EBX_REG_24_;
  assign n66316 = n66297 & n66315;
  assign n66317 = P2_P3_EBX_REG_25_ & ~n66316;
  assign n66318 = ~P2_P3_EBX_REG_25_ & n66316;
  assign n66319 = ~n66317 & ~n66318;
  assign n66320 = n66080 & ~n66319;
  assign n66321 = ~n66313 & ~n66314;
  assign n11961 = n66320 | ~n66321;
  assign n66323 = P2_P3_EBX_REG_26_ & ~n66079;
  assign n66324 = ~n65864 & n66082;
  assign n66325 = P2_P3_EBX_REG_25_ & n66316;
  assign n66326 = ~P2_P3_EBX_REG_26_ & n66325;
  assign n66327 = P2_P3_EBX_REG_26_ & ~n66325;
  assign n66328 = ~n66326 & ~n66327;
  assign n66329 = n66080 & ~n66328;
  assign n66330 = ~n66323 & ~n66324;
  assign n11966 = n66329 | ~n66330;
  assign n66332 = P2_P3_EBX_REG_27_ & ~n66079;
  assign n66333 = ~n65912 & n66082;
  assign n66334 = P2_P3_EBX_REG_25_ & P2_P3_EBX_REG_26_;
  assign n66335 = n66316 & n66334;
  assign n66336 = P2_P3_EBX_REG_27_ & ~n66335;
  assign n66337 = ~P2_P3_EBX_REG_27_ & n66335;
  assign n66338 = ~n66336 & ~n66337;
  assign n66339 = n66080 & ~n66338;
  assign n66340 = ~n66332 & ~n66333;
  assign n11971 = n66339 | ~n66340;
  assign n66342 = P2_P3_EBX_REG_28_ & ~n66079;
  assign n66343 = ~n65961 & n66082;
  assign n66344 = P2_P3_EBX_REG_27_ & n66335;
  assign n66345 = ~P2_P3_EBX_REG_28_ & n66344;
  assign n66346 = P2_P3_EBX_REG_28_ & ~n66344;
  assign n66347 = ~n66345 & ~n66346;
  assign n66348 = n66080 & ~n66347;
  assign n66349 = ~n66342 & ~n66343;
  assign n11976 = n66348 | ~n66349;
  assign n66351 = P2_P3_EBX_REG_29_ & ~n66079;
  assign n66352 = ~n66009 & n66082;
  assign n66353 = P2_P3_EBX_REG_27_ & P2_P3_EBX_REG_28_;
  assign n66354 = n66335 & n66353;
  assign n66355 = P2_P3_EBX_REG_29_ & ~n66354;
  assign n66356 = ~P2_P3_EBX_REG_29_ & n66354;
  assign n66357 = ~n66355 & ~n66356;
  assign n66358 = n66080 & ~n66357;
  assign n66359 = ~n66351 & ~n66352;
  assign n11981 = n66358 | ~n66359;
  assign n66361 = P2_P3_EBX_REG_30_ & ~n66079;
  assign n66362 = ~n66058 & n66082;
  assign n66363 = P2_P3_EBX_REG_29_ & n66354;
  assign n66364 = ~P2_P3_EBX_REG_30_ & n66363;
  assign n66365 = P2_P3_EBX_REG_30_ & ~n66363;
  assign n66366 = ~n66364 & ~n66365;
  assign n66367 = n66080 & ~n66366;
  assign n66368 = ~n66361 & ~n66362;
  assign n11986 = n66367 | ~n66368;
  assign n66370 = P2_P3_EBX_REG_31_ & ~n66079;
  assign n66371 = P2_P3_EBX_REG_30_ & n66363;
  assign n66372 = ~P2_P3_EBX_REG_31_ & n66371;
  assign n66373 = P2_P3_EBX_REG_31_ & ~n66371;
  assign n66374 = ~n66372 & ~n66373;
  assign n66375 = n66080 & ~n66374;
  assign n11991 = n66370 | n66375;
  assign n66377 = ~n59332 & ~n59371;
  assign n66378 = ~n60935 & n66377;
  assign n66379 = n59199 & n59207;
  assign n66380 = n59321 & ~n66379;
  assign n66381 = n66378 & ~n66380;
  assign n66382 = P2_P3_STATE2_REG_2_ & ~n66381;
  assign n66383 = n59049 & n66382;
  assign n66384 = ~n58682 & n66383;
  assign n66385 = ~P2_P3_EBX_REG_31_ & n66384;
  assign n66386 = n58967 & n66382;
  assign n66387 = ~n58685 & n66386;
  assign n66388 = n58685 & n66386;
  assign n66389 = ~n58682 & n66388;
  assign n66390 = ~n66385 & ~n66387;
  assign n66391 = ~n66389 & n66390;
  assign n66392 = P2_P3_EBX_REG_0_ & ~n66391;
  assign n66393 = n58682 & n66388;
  assign n66394 = P2_P3_REIP_REG_0_ & n66393;
  assign n66395 = P2_P3_EBX_REG_31_ & n66384;
  assign n66396 = P2_P3_EBX_REG_0_ & n66395;
  assign n66397 = n59044 & n66382;
  assign n66398 = ~P2_P3_INSTQUEUERD_ADDR_REG_0_ & n66397;
  assign n66399 = n59040 & n66382;
  assign n66400 = ~P2_P3_INSTQUEUERD_ADDR_REG_0_ & n66399;
  assign n66401 = ~n66398 & ~n66400;
  assign n66402 = ~n66394 & ~n66396;
  assign n66403 = n66401 & n66402;
  assign n66404 = n58682 & n66383;
  assign n66405 = P2_P3_REIP_REG_0_ & n66404;
  assign n66406 = P2_P3_STATE2_REG_1_ & ~n66381;
  assign n66407 = n64518 & n66406;
  assign n66408 = P2_P3_PHYADDRPOINTER_REG_0_ & n66407;
  assign n66409 = P2_P3_REIP_REG_0_ & n66381;
  assign n66410 = P2_P3_STATE2_REG_3_ & ~n66381;
  assign n66411 = P2_P3_PHYADDRPOINTER_REG_0_ & n66410;
  assign n66412 = ~n66409 & ~n66411;
  assign n66413 = ~n64518 & n66406;
  assign n66414 = P2_P3_PHYADDRPOINTER_REG_0_ & n66413;
  assign n66415 = n66412 & ~n66414;
  assign n66416 = ~n66392 & n66403;
  assign n66417 = ~n66405 & n66416;
  assign n66418 = ~n66408 & n66417;
  assign n11996 = ~n66415 | ~n66418;
  assign n66420 = P2_P3_EBX_REG_1_ & ~n66391;
  assign n66421 = ~P2_P3_REIP_REG_1_ & n66393;
  assign n66422 = ~n66089 & n66395;
  assign n66423 = ~n58691 & ~n58696;
  assign n66424 = n66397 & ~n66423;
  assign n66425 = n66399 & ~n66423;
  assign n66426 = ~n66424 & ~n66425;
  assign n66427 = ~n66421 & ~n66422;
  assign n66428 = n66426 & n66427;
  assign n66429 = ~P2_P3_REIP_REG_1_ & n66404;
  assign n66430 = ~P2_P3_PHYADDRPOINTER_REG_1_ & n66407;
  assign n66431 = P2_P3_REIP_REG_1_ & n66381;
  assign n66432 = P2_P3_PHYADDRPOINTER_REG_1_ & n66410;
  assign n66433 = ~n66431 & ~n66432;
  assign n66434 = P2_P3_PHYADDRPOINTER_REG_0_ & P2_P3_PHYADDRPOINTER_REG_1_;
  assign n66435 = ~P2_P3_PHYADDRPOINTER_REG_0_ & ~P2_P3_PHYADDRPOINTER_REG_1_;
  assign n66436 = ~n66434 & ~n66435;
  assign n66437 = n66413 & ~n66436;
  assign n66438 = n66433 & ~n66437;
  assign n66439 = ~n66420 & n66428;
  assign n66440 = ~n66429 & n66439;
  assign n66441 = ~n66430 & n66440;
  assign n12001 = ~n66438 | ~n66441;
  assign n66443 = P2_P3_EBX_REG_2_ & ~n66391;
  assign n66444 = P2_P3_REIP_REG_1_ & ~P2_P3_REIP_REG_2_;
  assign n66445 = ~P2_P3_REIP_REG_1_ & P2_P3_REIP_REG_2_;
  assign n66446 = ~n66444 & ~n66445;
  assign n66447 = n66393 & ~n66446;
  assign n66448 = ~P2_P3_EBX_REG_0_ & ~P2_P3_EBX_REG_1_;
  assign n66449 = P2_P3_EBX_REG_2_ & ~n66448;
  assign n66450 = ~P2_P3_EBX_REG_2_ & n66448;
  assign n66451 = ~n66449 & ~n66450;
  assign n66452 = n66395 & n66451;
  assign n66453 = ~n59169 & n66397;
  assign n66454 = ~n59169 & n66399;
  assign n66455 = ~n66453 & ~n66454;
  assign n66456 = ~n66447 & ~n66452;
  assign n66457 = n66455 & n66456;
  assign n66458 = n66404 & ~n66446;
  assign n66459 = ~n63852 & n66407;
  assign n66460 = P2_P3_REIP_REG_2_ & n66381;
  assign n66461 = P2_P3_PHYADDRPOINTER_REG_2_ & n66410;
  assign n66462 = ~n66460 & ~n66461;
  assign n66463 = ~P2_P3_PHYADDRPOINTER_REG_0_ & P2_P3_PHYADDRPOINTER_REG_1_;
  assign n66464 = ~n63852 & ~n66463;
  assign n66465 = n63852 & n66463;
  assign n66466 = ~n66464 & ~n66465;
  assign n66467 = n66413 & n66466;
  assign n66468 = n66462 & ~n66467;
  assign n66469 = ~n66443 & n66457;
  assign n66470 = ~n66458 & n66469;
  assign n66471 = ~n66459 & n66470;
  assign n12006 = ~n66468 | ~n66471;
  assign n66473 = P2_P3_EBX_REG_3_ & ~n66391;
  assign n66474 = P2_P3_REIP_REG_1_ & P2_P3_REIP_REG_2_;
  assign n66475 = ~P2_P3_REIP_REG_3_ & n66474;
  assign n66476 = P2_P3_REIP_REG_3_ & ~n66474;
  assign n66477 = ~n66475 & ~n66476;
  assign n66478 = n66393 & ~n66477;
  assign n66479 = ~P2_P3_EBX_REG_3_ & n66450;
  assign n66480 = P2_P3_EBX_REG_3_ & ~n66450;
  assign n66481 = ~n66479 & ~n66480;
  assign n66482 = n66395 & n66481;
  assign n66483 = ~P2_P3_INSTQUEUERD_ADDR_REG_3_ & n59217;
  assign n66484 = ~n59218 & ~n66483;
  assign n66485 = n66397 & ~n66484;
  assign n66486 = n66399 & ~n66484;
  assign n66487 = ~n66485 & ~n66486;
  assign n66488 = ~n66478 & ~n66482;
  assign n66489 = n66487 & n66488;
  assign n66490 = n66404 & ~n66477;
  assign n66491 = ~n63874 & n66407;
  assign n66492 = P2_P3_REIP_REG_3_ & n66381;
  assign n66493 = P2_P3_PHYADDRPOINTER_REG_3_ & n66410;
  assign n66494 = ~n66492 & ~n66493;
  assign n66495 = n63874 & n66465;
  assign n66496 = ~n63874 & ~n66465;
  assign n66497 = ~n66495 & ~n66496;
  assign n66498 = n66413 & n66497;
  assign n66499 = n66494 & ~n66498;
  assign n66500 = ~n66473 & n66489;
  assign n66501 = ~n66490 & n66500;
  assign n66502 = ~n66491 & n66501;
  assign n12011 = ~n66499 | ~n66502;
  assign n66504 = P2_P3_INSTQUEUERD_ADDR_REG_3_ & n59217;
  assign n66505 = ~P2_P3_INSTQUEUERD_ADDR_REG_4_ & n66504;
  assign n66506 = P2_P3_INSTQUEUERD_ADDR_REG_4_ & ~n66504;
  assign n66507 = ~n66505 & ~n66506;
  assign n66508 = n66399 & ~n66507;
  assign n66509 = n66397 & ~n66507;
  assign n66510 = ~n66508 & ~n66509;
  assign n66511 = P2_P3_EBX_REG_4_ & ~n66391;
  assign n66512 = P2_P3_EBX_REG_4_ & ~n66479;
  assign n66513 = ~P2_P3_EBX_REG_3_ & ~P2_P3_EBX_REG_4_;
  assign n66514 = n66450 & n66513;
  assign n66515 = ~n66512 & ~n66514;
  assign n66516 = n66395 & n66515;
  assign n66517 = n60934 & ~n66381;
  assign n66518 = P2_P3_REIP_REG_3_ & n66474;
  assign n66519 = ~P2_P3_REIP_REG_4_ & n66518;
  assign n66520 = P2_P3_REIP_REG_4_ & ~n66518;
  assign n66521 = ~n66519 & ~n66520;
  assign n66522 = n66393 & ~n66521;
  assign n66523 = ~n66516 & ~n66517;
  assign n66524 = ~n66522 & n66523;
  assign n66525 = n66404 & ~n66521;
  assign n66526 = ~n63895 & n66407;
  assign n66527 = n66510 & ~n66511;
  assign n66528 = n66524 & n66527;
  assign n66529 = ~n66525 & n66528;
  assign n66530 = ~n66526 & n66529;
  assign n66531 = P2_P3_REIP_REG_4_ & n66381;
  assign n66532 = P2_P3_PHYADDRPOINTER_REG_4_ & n66410;
  assign n66533 = ~n66531 & ~n66532;
  assign n66534 = ~n63895 & ~n66495;
  assign n66535 = n63874 & n63895;
  assign n66536 = n66465 & n66535;
  assign n66537 = ~n66534 & ~n66536;
  assign n66538 = n66413 & n66537;
  assign n66539 = n66533 & ~n66538;
  assign n12016 = ~n66530 | ~n66539;
  assign n66541 = P2_P3_INSTQUEUERD_ADDR_REG_4_ & n66504;
  assign n66542 = n66399 & n66541;
  assign n66543 = n66397 & n66541;
  assign n66544 = ~n66542 & ~n66543;
  assign n66545 = P2_P3_EBX_REG_5_ & ~n66391;
  assign n66546 = ~P2_P3_EBX_REG_5_ & n66514;
  assign n66547 = P2_P3_EBX_REG_5_ & ~n66514;
  assign n66548 = ~n66546 & ~n66547;
  assign n66549 = n66395 & n66548;
  assign n66550 = P2_P3_REIP_REG_4_ & n66518;
  assign n66551 = ~P2_P3_REIP_REG_5_ & n66550;
  assign n66552 = P2_P3_REIP_REG_5_ & ~n66550;
  assign n66553 = ~n66551 & ~n66552;
  assign n66554 = n66393 & ~n66553;
  assign n66555 = ~n66517 & ~n66549;
  assign n66556 = ~n66554 & n66555;
  assign n66557 = n66404 & ~n66553;
  assign n66558 = ~n63918 & n66407;
  assign n66559 = n66544 & ~n66545;
  assign n66560 = n66556 & n66559;
  assign n66561 = ~n66557 & n66560;
  assign n66562 = ~n66558 & n66561;
  assign n66563 = P2_P3_REIP_REG_5_ & n66381;
  assign n66564 = P2_P3_PHYADDRPOINTER_REG_5_ & n66410;
  assign n66565 = ~n66563 & ~n66564;
  assign n66566 = n63918 & n66536;
  assign n66567 = ~n63918 & ~n66536;
  assign n66568 = ~n66566 & ~n66567;
  assign n66569 = n66413 & n66568;
  assign n66570 = n66565 & ~n66569;
  assign n12021 = ~n66562 | ~n66570;
  assign n66572 = P2_P3_REIP_REG_5_ & n66550;
  assign n66573 = ~P2_P3_REIP_REG_6_ & n66572;
  assign n66574 = P2_P3_REIP_REG_6_ & ~n66572;
  assign n66575 = ~n66573 & ~n66574;
  assign n66576 = n66404 & ~n66575;
  assign n66577 = P2_P3_EBX_REG_6_ & ~n66391;
  assign n66578 = P2_P3_EBX_REG_6_ & ~n66546;
  assign n66579 = ~P2_P3_EBX_REG_5_ & ~P2_P3_EBX_REG_6_;
  assign n66580 = n66514 & n66579;
  assign n66581 = ~n66578 & ~n66580;
  assign n66582 = n66395 & n66581;
  assign n66583 = n66393 & ~n66575;
  assign n66584 = ~n66517 & ~n66582;
  assign n66585 = ~n66583 & n66584;
  assign n66586 = ~n63941 & ~n66566;
  assign n66587 = n63918 & n63941;
  assign n66588 = n66536 & n66587;
  assign n66589 = ~n66586 & ~n66588;
  assign n66590 = n66413 & n66589;
  assign n66591 = P2_P3_REIP_REG_6_ & n66381;
  assign n66592 = P2_P3_PHYADDRPOINTER_REG_6_ & n66410;
  assign n66593 = ~n66591 & ~n66592;
  assign n66594 = ~n63941 & n66407;
  assign n66595 = n66593 & ~n66594;
  assign n66596 = ~n66576 & ~n66577;
  assign n66597 = n66585 & n66596;
  assign n66598 = ~n66590 & n66597;
  assign n12026 = ~n66595 | ~n66598;
  assign n66600 = P2_P3_REIP_REG_6_ & n66572;
  assign n66601 = ~P2_P3_REIP_REG_7_ & n66600;
  assign n66602 = P2_P3_REIP_REG_7_ & ~n66600;
  assign n66603 = ~n66601 & ~n66602;
  assign n66604 = n66404 & ~n66603;
  assign n66605 = P2_P3_EBX_REG_7_ & ~n66391;
  assign n66606 = ~P2_P3_EBX_REG_7_ & n66580;
  assign n66607 = P2_P3_EBX_REG_7_ & ~n66580;
  assign n66608 = ~n66606 & ~n66607;
  assign n66609 = n66395 & n66608;
  assign n66610 = n66393 & ~n66603;
  assign n66611 = ~n66517 & ~n66609;
  assign n66612 = ~n66610 & n66611;
  assign n66613 = n63964 & n66588;
  assign n66614 = ~n63964 & ~n66588;
  assign n66615 = ~n66613 & ~n66614;
  assign n66616 = n66413 & n66615;
  assign n66617 = P2_P3_REIP_REG_7_ & n66381;
  assign n66618 = P2_P3_PHYADDRPOINTER_REG_7_ & n66410;
  assign n66619 = ~n66617 & ~n66618;
  assign n66620 = ~n63964 & n66407;
  assign n66621 = n66619 & ~n66620;
  assign n66622 = ~n66604 & ~n66605;
  assign n66623 = n66612 & n66622;
  assign n66624 = ~n66616 & n66623;
  assign n12031 = ~n66621 | ~n66624;
  assign n66626 = P2_P3_REIP_REG_7_ & n66600;
  assign n66627 = ~P2_P3_REIP_REG_8_ & n66626;
  assign n66628 = P2_P3_REIP_REG_8_ & ~n66626;
  assign n66629 = ~n66627 & ~n66628;
  assign n66630 = n66404 & ~n66629;
  assign n66631 = P2_P3_EBX_REG_8_ & ~n66391;
  assign n66632 = P2_P3_EBX_REG_8_ & ~n66606;
  assign n66633 = ~P2_P3_EBX_REG_7_ & ~P2_P3_EBX_REG_8_;
  assign n66634 = n66580 & n66633;
  assign n66635 = ~n66632 & ~n66634;
  assign n66636 = n66395 & n66635;
  assign n66637 = n66393 & ~n66629;
  assign n66638 = ~n66517 & ~n66636;
  assign n66639 = ~n66637 & n66638;
  assign n66640 = ~n63987 & ~n66613;
  assign n66641 = n63964 & n63987;
  assign n66642 = n66588 & n66641;
  assign n66643 = ~n66640 & ~n66642;
  assign n66644 = n66413 & n66643;
  assign n66645 = P2_P3_REIP_REG_8_ & n66381;
  assign n66646 = P2_P3_PHYADDRPOINTER_REG_8_ & n66410;
  assign n66647 = ~n66645 & ~n66646;
  assign n66648 = ~n63987 & n66407;
  assign n66649 = n66647 & ~n66648;
  assign n66650 = ~n66630 & ~n66631;
  assign n66651 = n66639 & n66650;
  assign n66652 = ~n66644 & n66651;
  assign n12036 = ~n66649 | ~n66652;
  assign n66654 = P2_P3_REIP_REG_8_ & n66626;
  assign n66655 = ~P2_P3_REIP_REG_9_ & n66654;
  assign n66656 = P2_P3_REIP_REG_9_ & ~n66654;
  assign n66657 = ~n66655 & ~n66656;
  assign n66658 = n66404 & ~n66657;
  assign n66659 = P2_P3_EBX_REG_9_ & ~n66391;
  assign n66660 = ~P2_P3_EBX_REG_9_ & n66634;
  assign n66661 = P2_P3_EBX_REG_9_ & ~n66634;
  assign n66662 = ~n66660 & ~n66661;
  assign n66663 = n66395 & n66662;
  assign n66664 = n66393 & ~n66657;
  assign n66665 = ~n66517 & ~n66663;
  assign n66666 = ~n66664 & n66665;
  assign n66667 = n64010 & n66642;
  assign n66668 = ~n64010 & ~n66642;
  assign n66669 = ~n66667 & ~n66668;
  assign n66670 = n66413 & n66669;
  assign n66671 = P2_P3_REIP_REG_9_ & n66381;
  assign n66672 = P2_P3_PHYADDRPOINTER_REG_9_ & n66410;
  assign n66673 = ~n66671 & ~n66672;
  assign n66674 = ~n64010 & n66407;
  assign n66675 = n66673 & ~n66674;
  assign n66676 = ~n66658 & ~n66659;
  assign n66677 = n66666 & n66676;
  assign n66678 = ~n66670 & n66677;
  assign n12041 = ~n66675 | ~n66678;
  assign n66680 = P2_P3_REIP_REG_9_ & n66654;
  assign n66681 = ~P2_P3_REIP_REG_10_ & n66680;
  assign n66682 = P2_P3_REIP_REG_10_ & ~n66680;
  assign n66683 = ~n66681 & ~n66682;
  assign n66684 = n66404 & ~n66683;
  assign n66685 = P2_P3_EBX_REG_10_ & ~n66391;
  assign n66686 = P2_P3_EBX_REG_10_ & ~n66660;
  assign n66687 = ~P2_P3_EBX_REG_9_ & ~P2_P3_EBX_REG_10_;
  assign n66688 = n66634 & n66687;
  assign n66689 = ~n66686 & ~n66688;
  assign n66690 = n66395 & n66689;
  assign n66691 = n66393 & ~n66683;
  assign n66692 = ~n66517 & ~n66690;
  assign n66693 = ~n66691 & n66692;
  assign n66694 = ~n64033 & ~n66667;
  assign n66695 = n64010 & n64033;
  assign n66696 = n66642 & n66695;
  assign n66697 = ~n66694 & ~n66696;
  assign n66698 = n66413 & n66697;
  assign n66699 = P2_P3_REIP_REG_10_ & n66381;
  assign n66700 = P2_P3_PHYADDRPOINTER_REG_10_ & n66410;
  assign n66701 = ~n66699 & ~n66700;
  assign n66702 = ~n64033 & n66407;
  assign n66703 = n66701 & ~n66702;
  assign n66704 = ~n66684 & ~n66685;
  assign n66705 = n66693 & n66704;
  assign n66706 = ~n66698 & n66705;
  assign n12046 = ~n66703 | ~n66706;
  assign n66708 = P2_P3_REIP_REG_10_ & n66680;
  assign n66709 = ~P2_P3_REIP_REG_11_ & n66708;
  assign n66710 = P2_P3_REIP_REG_11_ & ~n66708;
  assign n66711 = ~n66709 & ~n66710;
  assign n66712 = n66404 & ~n66711;
  assign n66713 = P2_P3_EBX_REG_11_ & ~n66391;
  assign n66714 = ~P2_P3_EBX_REG_11_ & n66688;
  assign n66715 = P2_P3_EBX_REG_11_ & ~n66688;
  assign n66716 = ~n66714 & ~n66715;
  assign n66717 = n66395 & n66716;
  assign n66718 = n66393 & ~n66711;
  assign n66719 = ~n66517 & ~n66717;
  assign n66720 = ~n66718 & n66719;
  assign n66721 = n64056 & n66696;
  assign n66722 = ~n64056 & ~n66696;
  assign n66723 = ~n66721 & ~n66722;
  assign n66724 = n66413 & n66723;
  assign n66725 = P2_P3_REIP_REG_11_ & n66381;
  assign n66726 = P2_P3_PHYADDRPOINTER_REG_11_ & n66410;
  assign n66727 = ~n66725 & ~n66726;
  assign n66728 = ~n64056 & n66407;
  assign n66729 = n66727 & ~n66728;
  assign n66730 = ~n66712 & ~n66713;
  assign n66731 = n66720 & n66730;
  assign n66732 = ~n66724 & n66731;
  assign n12051 = ~n66729 | ~n66732;
  assign n66734 = P2_P3_REIP_REG_11_ & n66708;
  assign n66735 = ~P2_P3_REIP_REG_12_ & n66734;
  assign n66736 = P2_P3_REIP_REG_12_ & ~n66734;
  assign n66737 = ~n66735 & ~n66736;
  assign n66738 = n66404 & ~n66737;
  assign n66739 = P2_P3_EBX_REG_12_ & ~n66391;
  assign n66740 = P2_P3_EBX_REG_12_ & ~n66714;
  assign n66741 = ~P2_P3_EBX_REG_11_ & ~P2_P3_EBX_REG_12_;
  assign n66742 = n66688 & n66741;
  assign n66743 = ~n66740 & ~n66742;
  assign n66744 = n66395 & n66743;
  assign n66745 = n66393 & ~n66737;
  assign n66746 = ~n66517 & ~n66744;
  assign n66747 = ~n66745 & n66746;
  assign n66748 = ~n64079 & ~n66721;
  assign n66749 = n64056 & n64079;
  assign n66750 = n66696 & n66749;
  assign n66751 = ~n66748 & ~n66750;
  assign n66752 = n66413 & n66751;
  assign n66753 = P2_P3_REIP_REG_12_ & n66381;
  assign n66754 = P2_P3_PHYADDRPOINTER_REG_12_ & n66410;
  assign n66755 = ~n66753 & ~n66754;
  assign n66756 = ~n64079 & n66407;
  assign n66757 = n66755 & ~n66756;
  assign n66758 = ~n66738 & ~n66739;
  assign n66759 = n66747 & n66758;
  assign n66760 = ~n66752 & n66759;
  assign n12056 = ~n66757 | ~n66760;
  assign n66762 = P2_P3_REIP_REG_12_ & n66734;
  assign n66763 = ~P2_P3_REIP_REG_13_ & n66762;
  assign n66764 = P2_P3_REIP_REG_13_ & ~n66762;
  assign n66765 = ~n66763 & ~n66764;
  assign n66766 = n66404 & ~n66765;
  assign n66767 = P2_P3_EBX_REG_13_ & ~n66391;
  assign n66768 = ~P2_P3_EBX_REG_13_ & n66742;
  assign n66769 = P2_P3_EBX_REG_13_ & ~n66742;
  assign n66770 = ~n66768 & ~n66769;
  assign n66771 = n66395 & n66770;
  assign n66772 = n66393 & ~n66765;
  assign n66773 = ~n66517 & ~n66771;
  assign n66774 = ~n66772 & n66773;
  assign n66775 = n64102 & n66750;
  assign n66776 = ~n64102 & ~n66750;
  assign n66777 = ~n66775 & ~n66776;
  assign n66778 = n66413 & n66777;
  assign n66779 = P2_P3_REIP_REG_13_ & n66381;
  assign n66780 = P2_P3_PHYADDRPOINTER_REG_13_ & n66410;
  assign n66781 = ~n66779 & ~n66780;
  assign n66782 = ~n64102 & n66407;
  assign n66783 = n66781 & ~n66782;
  assign n66784 = ~n66766 & ~n66767;
  assign n66785 = n66774 & n66784;
  assign n66786 = ~n66778 & n66785;
  assign n12061 = ~n66783 | ~n66786;
  assign n66788 = P2_P3_REIP_REG_13_ & n66762;
  assign n66789 = ~P2_P3_REIP_REG_14_ & n66788;
  assign n66790 = P2_P3_REIP_REG_14_ & ~n66788;
  assign n66791 = ~n66789 & ~n66790;
  assign n66792 = n66404 & ~n66791;
  assign n66793 = P2_P3_EBX_REG_14_ & ~n66391;
  assign n66794 = P2_P3_EBX_REG_14_ & ~n66768;
  assign n66795 = ~P2_P3_EBX_REG_13_ & ~P2_P3_EBX_REG_14_;
  assign n66796 = n66742 & n66795;
  assign n66797 = ~n66794 & ~n66796;
  assign n66798 = n66395 & n66797;
  assign n66799 = n66393 & ~n66791;
  assign n66800 = ~n66517 & ~n66798;
  assign n66801 = ~n66799 & n66800;
  assign n66802 = ~n64125 & ~n66775;
  assign n66803 = n64102 & n64125;
  assign n66804 = n66750 & n66803;
  assign n66805 = ~n66802 & ~n66804;
  assign n66806 = n66413 & n66805;
  assign n66807 = P2_P3_REIP_REG_14_ & n66381;
  assign n66808 = P2_P3_PHYADDRPOINTER_REG_14_ & n66410;
  assign n66809 = ~n66807 & ~n66808;
  assign n66810 = ~n64125 & n66407;
  assign n66811 = n66809 & ~n66810;
  assign n66812 = ~n66792 & ~n66793;
  assign n66813 = n66801 & n66812;
  assign n66814 = ~n66806 & n66813;
  assign n12066 = ~n66811 | ~n66814;
  assign n66816 = P2_P3_REIP_REG_14_ & n66788;
  assign n66817 = ~P2_P3_REIP_REG_15_ & n66816;
  assign n66818 = P2_P3_REIP_REG_15_ & ~n66816;
  assign n66819 = ~n66817 & ~n66818;
  assign n66820 = n66404 & ~n66819;
  assign n66821 = P2_P3_EBX_REG_15_ & ~n66391;
  assign n66822 = ~P2_P3_EBX_REG_15_ & n66796;
  assign n66823 = P2_P3_EBX_REG_15_ & ~n66796;
  assign n66824 = ~n66822 & ~n66823;
  assign n66825 = n66395 & n66824;
  assign n66826 = n66393 & ~n66819;
  assign n66827 = ~n66517 & ~n66825;
  assign n66828 = ~n66826 & n66827;
  assign n66829 = n64148 & n66804;
  assign n66830 = ~n64148 & ~n66804;
  assign n66831 = ~n66829 & ~n66830;
  assign n66832 = n66413 & n66831;
  assign n66833 = P2_P3_REIP_REG_15_ & n66381;
  assign n66834 = P2_P3_PHYADDRPOINTER_REG_15_ & n66410;
  assign n66835 = ~n66833 & ~n66834;
  assign n66836 = ~n64148 & n66407;
  assign n66837 = n66835 & ~n66836;
  assign n66838 = ~n66820 & ~n66821;
  assign n66839 = n66828 & n66838;
  assign n66840 = ~n66832 & n66839;
  assign n12071 = ~n66837 | ~n66840;
  assign n66842 = P2_P3_REIP_REG_15_ & n66816;
  assign n66843 = ~P2_P3_REIP_REG_16_ & n66842;
  assign n66844 = P2_P3_REIP_REG_16_ & ~n66842;
  assign n66845 = ~n66843 & ~n66844;
  assign n66846 = n66404 & ~n66845;
  assign n66847 = P2_P3_EBX_REG_16_ & ~n66391;
  assign n66848 = P2_P3_EBX_REG_16_ & ~n66822;
  assign n66849 = ~P2_P3_EBX_REG_15_ & ~P2_P3_EBX_REG_16_;
  assign n66850 = n66796 & n66849;
  assign n66851 = ~n66848 & ~n66850;
  assign n66852 = n66395 & n66851;
  assign n66853 = n66393 & ~n66845;
  assign n66854 = ~n66517 & ~n66852;
  assign n66855 = ~n66853 & n66854;
  assign n66856 = ~n64171 & ~n66829;
  assign n66857 = n64148 & n64171;
  assign n66858 = n66804 & n66857;
  assign n66859 = ~n66856 & ~n66858;
  assign n66860 = n66413 & n66859;
  assign n66861 = P2_P3_REIP_REG_16_ & n66381;
  assign n66862 = P2_P3_PHYADDRPOINTER_REG_16_ & n66410;
  assign n66863 = ~n66861 & ~n66862;
  assign n66864 = ~n64171 & n66407;
  assign n66865 = n66863 & ~n66864;
  assign n66866 = ~n66846 & ~n66847;
  assign n66867 = n66855 & n66866;
  assign n66868 = ~n66860 & n66867;
  assign n12076 = ~n66865 | ~n66868;
  assign n66870 = P2_P3_REIP_REG_16_ & n66842;
  assign n66871 = ~P2_P3_REIP_REG_17_ & n66870;
  assign n66872 = P2_P3_REIP_REG_17_ & ~n66870;
  assign n66873 = ~n66871 & ~n66872;
  assign n66874 = n66404 & ~n66873;
  assign n66875 = P2_P3_EBX_REG_17_ & ~n66391;
  assign n66876 = ~P2_P3_EBX_REG_17_ & n66850;
  assign n66877 = P2_P3_EBX_REG_17_ & ~n66850;
  assign n66878 = ~n66876 & ~n66877;
  assign n66879 = n66395 & n66878;
  assign n66880 = n66393 & ~n66873;
  assign n66881 = ~n66517 & ~n66879;
  assign n66882 = ~n66880 & n66881;
  assign n66883 = n64194 & n66858;
  assign n66884 = ~n64194 & ~n66858;
  assign n66885 = ~n66883 & ~n66884;
  assign n66886 = n66413 & n66885;
  assign n66887 = P2_P3_REIP_REG_17_ & n66381;
  assign n66888 = P2_P3_PHYADDRPOINTER_REG_17_ & n66410;
  assign n66889 = ~n66887 & ~n66888;
  assign n66890 = ~n64194 & n66407;
  assign n66891 = n66889 & ~n66890;
  assign n66892 = ~n66874 & ~n66875;
  assign n66893 = n66882 & n66892;
  assign n66894 = ~n66886 & n66893;
  assign n12081 = ~n66891 | ~n66894;
  assign n66896 = P2_P3_REIP_REG_17_ & n66870;
  assign n66897 = ~P2_P3_REIP_REG_18_ & n66896;
  assign n66898 = P2_P3_REIP_REG_18_ & ~n66896;
  assign n66899 = ~n66897 & ~n66898;
  assign n66900 = n66404 & ~n66899;
  assign n66901 = P2_P3_EBX_REG_18_ & ~n66391;
  assign n66902 = P2_P3_EBX_REG_18_ & ~n66876;
  assign n66903 = ~P2_P3_EBX_REG_17_ & ~P2_P3_EBX_REG_18_;
  assign n66904 = n66850 & n66903;
  assign n66905 = ~n66902 & ~n66904;
  assign n66906 = n66395 & n66905;
  assign n66907 = n66393 & ~n66899;
  assign n66908 = ~n66517 & ~n66906;
  assign n66909 = ~n66907 & n66908;
  assign n66910 = ~n64217 & ~n66883;
  assign n66911 = n64194 & n64217;
  assign n66912 = n66858 & n66911;
  assign n66913 = ~n66910 & ~n66912;
  assign n66914 = n66413 & n66913;
  assign n66915 = P2_P3_REIP_REG_18_ & n66381;
  assign n66916 = P2_P3_PHYADDRPOINTER_REG_18_ & n66410;
  assign n66917 = ~n66915 & ~n66916;
  assign n66918 = ~n64217 & n66407;
  assign n66919 = n66917 & ~n66918;
  assign n66920 = ~n66900 & ~n66901;
  assign n66921 = n66909 & n66920;
  assign n66922 = ~n66914 & n66921;
  assign n12086 = ~n66919 | ~n66922;
  assign n66924 = P2_P3_REIP_REG_18_ & n66896;
  assign n66925 = ~P2_P3_REIP_REG_19_ & n66924;
  assign n66926 = P2_P3_REIP_REG_19_ & ~n66924;
  assign n66927 = ~n66925 & ~n66926;
  assign n66928 = n66404 & ~n66927;
  assign n66929 = P2_P3_EBX_REG_19_ & ~n66391;
  assign n66930 = ~P2_P3_EBX_REG_19_ & n66904;
  assign n66931 = P2_P3_EBX_REG_19_ & ~n66904;
  assign n66932 = ~n66930 & ~n66931;
  assign n66933 = n66395 & n66932;
  assign n66934 = n66393 & ~n66927;
  assign n66935 = ~n66517 & ~n66933;
  assign n66936 = ~n66934 & n66935;
  assign n66937 = n64240 & n66912;
  assign n66938 = ~n64240 & ~n66912;
  assign n66939 = ~n66937 & ~n66938;
  assign n66940 = n66413 & n66939;
  assign n66941 = P2_P3_REIP_REG_19_ & n66381;
  assign n66942 = P2_P3_PHYADDRPOINTER_REG_19_ & n66410;
  assign n66943 = ~n66941 & ~n66942;
  assign n66944 = ~n64240 & n66407;
  assign n66945 = n66943 & ~n66944;
  assign n66946 = ~n66928 & ~n66929;
  assign n66947 = n66936 & n66946;
  assign n66948 = ~n66940 & n66947;
  assign n12091 = ~n66945 | ~n66948;
  assign n66950 = P2_P3_REIP_REG_19_ & n66924;
  assign n66951 = ~P2_P3_REIP_REG_20_ & n66950;
  assign n66952 = P2_P3_REIP_REG_20_ & ~n66950;
  assign n66953 = ~n66951 & ~n66952;
  assign n66954 = n66404 & ~n66953;
  assign n66955 = P2_P3_EBX_REG_20_ & ~n66391;
  assign n66956 = n66393 & ~n66953;
  assign n66957 = P2_P3_EBX_REG_20_ & ~n66930;
  assign n66958 = ~P2_P3_EBX_REG_19_ & ~P2_P3_EBX_REG_20_;
  assign n66959 = n66904 & n66958;
  assign n66960 = ~n66957 & ~n66959;
  assign n66961 = n66395 & n66960;
  assign n66962 = ~n66956 & ~n66961;
  assign n66963 = ~n64263 & ~n66937;
  assign n66964 = n64240 & n64263;
  assign n66965 = n66912 & n66964;
  assign n66966 = ~n66963 & ~n66965;
  assign n66967 = n66413 & n66966;
  assign n66968 = P2_P3_REIP_REG_20_ & n66381;
  assign n66969 = P2_P3_PHYADDRPOINTER_REG_20_ & n66410;
  assign n66970 = ~n66968 & ~n66969;
  assign n66971 = ~n64263 & n66407;
  assign n66972 = n66970 & ~n66971;
  assign n66973 = ~n66954 & ~n66955;
  assign n66974 = n66962 & n66973;
  assign n66975 = ~n66967 & n66974;
  assign n12096 = ~n66972 | ~n66975;
  assign n66977 = P2_P3_REIP_REG_20_ & n66950;
  assign n66978 = ~P2_P3_REIP_REG_21_ & n66977;
  assign n66979 = P2_P3_REIP_REG_21_ & ~n66977;
  assign n66980 = ~n66978 & ~n66979;
  assign n66981 = n66404 & ~n66980;
  assign n66982 = P2_P3_EBX_REG_21_ & ~n66391;
  assign n66983 = n66393 & ~n66980;
  assign n66984 = ~P2_P3_EBX_REG_21_ & n66959;
  assign n66985 = P2_P3_EBX_REG_21_ & ~n66959;
  assign n66986 = ~n66984 & ~n66985;
  assign n66987 = n66395 & n66986;
  assign n66988 = ~n66983 & ~n66987;
  assign n66989 = n64286 & n66965;
  assign n66990 = ~n64286 & ~n66965;
  assign n66991 = ~n66989 & ~n66990;
  assign n66992 = n66413 & n66991;
  assign n66993 = P2_P3_REIP_REG_21_ & n66381;
  assign n66994 = P2_P3_PHYADDRPOINTER_REG_21_ & n66410;
  assign n66995 = ~n66993 & ~n66994;
  assign n66996 = ~n64286 & n66407;
  assign n66997 = n66995 & ~n66996;
  assign n66998 = ~n66981 & ~n66982;
  assign n66999 = n66988 & n66998;
  assign n67000 = ~n66992 & n66999;
  assign n12101 = ~n66997 | ~n67000;
  assign n67002 = P2_P3_REIP_REG_21_ & n66977;
  assign n67003 = ~P2_P3_REIP_REG_22_ & n67002;
  assign n67004 = P2_P3_REIP_REG_22_ & ~n67002;
  assign n67005 = ~n67003 & ~n67004;
  assign n67006 = n66404 & ~n67005;
  assign n67007 = P2_P3_EBX_REG_22_ & ~n66391;
  assign n67008 = n66393 & ~n67005;
  assign n67009 = P2_P3_EBX_REG_22_ & ~n66984;
  assign n67010 = ~P2_P3_EBX_REG_21_ & ~P2_P3_EBX_REG_22_;
  assign n67011 = n66959 & n67010;
  assign n67012 = ~n67009 & ~n67011;
  assign n67013 = n66395 & n67012;
  assign n67014 = ~n67008 & ~n67013;
  assign n67015 = ~n64310 & ~n66989;
  assign n67016 = n64286 & n64310;
  assign n67017 = n66965 & n67016;
  assign n67018 = ~n67015 & ~n67017;
  assign n67019 = n66413 & n67018;
  assign n67020 = P2_P3_REIP_REG_22_ & n66381;
  assign n67021 = P2_P3_PHYADDRPOINTER_REG_22_ & n66410;
  assign n67022 = ~n67020 & ~n67021;
  assign n67023 = ~n64310 & n66407;
  assign n67024 = n67022 & ~n67023;
  assign n67025 = ~n67006 & ~n67007;
  assign n67026 = n67014 & n67025;
  assign n67027 = ~n67019 & n67026;
  assign n12106 = ~n67024 | ~n67027;
  assign n67029 = P2_P3_REIP_REG_22_ & n67002;
  assign n67030 = ~P2_P3_REIP_REG_23_ & n67029;
  assign n67031 = P2_P3_REIP_REG_23_ & ~n67029;
  assign n67032 = ~n67030 & ~n67031;
  assign n67033 = n66404 & ~n67032;
  assign n67034 = P2_P3_EBX_REG_23_ & ~n66391;
  assign n67035 = n66393 & ~n67032;
  assign n67036 = ~P2_P3_EBX_REG_23_ & n67011;
  assign n67037 = P2_P3_EBX_REG_23_ & ~n67011;
  assign n67038 = ~n67036 & ~n67037;
  assign n67039 = n66395 & n67038;
  assign n67040 = ~n67035 & ~n67039;
  assign n67041 = n64333 & n67017;
  assign n67042 = ~n64333 & ~n67017;
  assign n67043 = ~n67041 & ~n67042;
  assign n67044 = n66413 & n67043;
  assign n67045 = P2_P3_REIP_REG_23_ & n66381;
  assign n67046 = P2_P3_PHYADDRPOINTER_REG_23_ & n66410;
  assign n67047 = ~n67045 & ~n67046;
  assign n67048 = ~n64333 & n66407;
  assign n67049 = n67047 & ~n67048;
  assign n67050 = ~n67033 & ~n67034;
  assign n67051 = n67040 & n67050;
  assign n67052 = ~n67044 & n67051;
  assign n12111 = ~n67049 | ~n67052;
  assign n67054 = P2_P3_REIP_REG_23_ & n67029;
  assign n67055 = ~P2_P3_REIP_REG_24_ & n67054;
  assign n67056 = P2_P3_REIP_REG_24_ & ~n67054;
  assign n67057 = ~n67055 & ~n67056;
  assign n67058 = n66404 & ~n67057;
  assign n67059 = P2_P3_EBX_REG_24_ & ~n66391;
  assign n67060 = n66393 & ~n67057;
  assign n67061 = P2_P3_EBX_REG_24_ & ~n67036;
  assign n67062 = ~P2_P3_EBX_REG_23_ & ~P2_P3_EBX_REG_24_;
  assign n67063 = n67011 & n67062;
  assign n67064 = ~n67061 & ~n67063;
  assign n67065 = n66395 & n67064;
  assign n67066 = ~n67060 & ~n67065;
  assign n67067 = ~n64356 & ~n67041;
  assign n67068 = n64333 & n64356;
  assign n67069 = n67017 & n67068;
  assign n67070 = ~n67067 & ~n67069;
  assign n67071 = n66413 & n67070;
  assign n67072 = P2_P3_REIP_REG_24_ & n66381;
  assign n67073 = P2_P3_PHYADDRPOINTER_REG_24_ & n66410;
  assign n67074 = ~n67072 & ~n67073;
  assign n67075 = ~n64356 & n66407;
  assign n67076 = n67074 & ~n67075;
  assign n67077 = ~n67058 & ~n67059;
  assign n67078 = n67066 & n67077;
  assign n67079 = ~n67071 & n67078;
  assign n12116 = ~n67076 | ~n67079;
  assign n67081 = P2_P3_REIP_REG_24_ & n67054;
  assign n67082 = ~P2_P3_REIP_REG_25_ & n67081;
  assign n67083 = P2_P3_REIP_REG_25_ & ~n67081;
  assign n67084 = ~n67082 & ~n67083;
  assign n67085 = n66404 & ~n67084;
  assign n67086 = P2_P3_EBX_REG_25_ & ~n66391;
  assign n67087 = n66393 & ~n67084;
  assign n67088 = ~P2_P3_EBX_REG_25_ & n67063;
  assign n67089 = P2_P3_EBX_REG_25_ & ~n67063;
  assign n67090 = ~n67088 & ~n67089;
  assign n67091 = n66395 & n67090;
  assign n67092 = ~n67087 & ~n67091;
  assign n67093 = n64379 & n67069;
  assign n67094 = ~n64379 & ~n67069;
  assign n67095 = ~n67093 & ~n67094;
  assign n67096 = n66413 & n67095;
  assign n67097 = P2_P3_REIP_REG_25_ & n66381;
  assign n67098 = P2_P3_PHYADDRPOINTER_REG_25_ & n66410;
  assign n67099 = ~n67097 & ~n67098;
  assign n67100 = ~n64379 & n66407;
  assign n67101 = n67099 & ~n67100;
  assign n67102 = ~n67085 & ~n67086;
  assign n67103 = n67092 & n67102;
  assign n67104 = ~n67096 & n67103;
  assign n12121 = ~n67101 | ~n67104;
  assign n67106 = P2_P3_REIP_REG_25_ & n67081;
  assign n67107 = ~P2_P3_REIP_REG_26_ & n67106;
  assign n67108 = P2_P3_REIP_REG_26_ & ~n67106;
  assign n67109 = ~n67107 & ~n67108;
  assign n67110 = n66404 & ~n67109;
  assign n67111 = P2_P3_EBX_REG_26_ & ~n66391;
  assign n67112 = n66393 & ~n67109;
  assign n67113 = P2_P3_EBX_REG_26_ & ~n67088;
  assign n67114 = ~P2_P3_EBX_REG_25_ & ~P2_P3_EBX_REG_26_;
  assign n67115 = n67063 & n67114;
  assign n67116 = ~n67113 & ~n67115;
  assign n67117 = n66395 & n67116;
  assign n67118 = ~n67112 & ~n67117;
  assign n67119 = ~n64402 & ~n67093;
  assign n67120 = n64379 & n64402;
  assign n67121 = n67069 & n67120;
  assign n67122 = ~n67119 & ~n67121;
  assign n67123 = n66413 & n67122;
  assign n67124 = P2_P3_REIP_REG_26_ & n66381;
  assign n67125 = P2_P3_PHYADDRPOINTER_REG_26_ & n66410;
  assign n67126 = ~n67124 & ~n67125;
  assign n67127 = ~n64402 & n66407;
  assign n67128 = n67126 & ~n67127;
  assign n67129 = ~n67110 & ~n67111;
  assign n67130 = n67118 & n67129;
  assign n67131 = ~n67123 & n67130;
  assign n12126 = ~n67128 | ~n67131;
  assign n67133 = P2_P3_REIP_REG_26_ & n67106;
  assign n67134 = ~P2_P3_REIP_REG_27_ & n67133;
  assign n67135 = P2_P3_REIP_REG_27_ & ~n67133;
  assign n67136 = ~n67134 & ~n67135;
  assign n67137 = n66404 & ~n67136;
  assign n67138 = P2_P3_EBX_REG_27_ & ~n66391;
  assign n67139 = n66393 & ~n67136;
  assign n67140 = ~P2_P3_EBX_REG_27_ & n67115;
  assign n67141 = P2_P3_EBX_REG_27_ & ~n67115;
  assign n67142 = ~n67140 & ~n67141;
  assign n67143 = n66395 & n67142;
  assign n67144 = ~n67139 & ~n67143;
  assign n67145 = n64425 & n67121;
  assign n67146 = ~n64425 & ~n67121;
  assign n67147 = ~n67145 & ~n67146;
  assign n67148 = n66413 & n67147;
  assign n67149 = P2_P3_REIP_REG_27_ & n66381;
  assign n67150 = P2_P3_PHYADDRPOINTER_REG_27_ & n66410;
  assign n67151 = ~n67149 & ~n67150;
  assign n67152 = ~n64425 & n66407;
  assign n67153 = n67151 & ~n67152;
  assign n67154 = ~n67137 & ~n67138;
  assign n67155 = n67144 & n67154;
  assign n67156 = ~n67148 & n67155;
  assign n12131 = ~n67153 | ~n67156;
  assign n67158 = P2_P3_REIP_REG_27_ & n67133;
  assign n67159 = ~P2_P3_REIP_REG_28_ & n67158;
  assign n67160 = P2_P3_REIP_REG_28_ & ~n67158;
  assign n67161 = ~n67159 & ~n67160;
  assign n67162 = n66404 & ~n67161;
  assign n67163 = P2_P3_EBX_REG_28_ & ~n66391;
  assign n67164 = n66393 & ~n67161;
  assign n67165 = P2_P3_EBX_REG_28_ & ~n67140;
  assign n67166 = ~P2_P3_EBX_REG_27_ & ~P2_P3_EBX_REG_28_;
  assign n67167 = n67115 & n67166;
  assign n67168 = ~n67165 & ~n67167;
  assign n67169 = n66395 & n67168;
  assign n67170 = ~n67164 & ~n67169;
  assign n67171 = ~n64449 & ~n67145;
  assign n67172 = n64425 & n64449;
  assign n67173 = n67121 & n67172;
  assign n67174 = ~n67171 & ~n67173;
  assign n67175 = n66413 & n67174;
  assign n67176 = P2_P3_REIP_REG_28_ & n66381;
  assign n67177 = P2_P3_PHYADDRPOINTER_REG_28_ & n66410;
  assign n67178 = ~n67176 & ~n67177;
  assign n67179 = ~n64449 & n66407;
  assign n67180 = n67178 & ~n67179;
  assign n67181 = ~n67162 & ~n67163;
  assign n67182 = n67170 & n67181;
  assign n67183 = ~n67175 & n67182;
  assign n12136 = ~n67180 | ~n67183;
  assign n67185 = P2_P3_REIP_REG_28_ & n67158;
  assign n67186 = ~P2_P3_REIP_REG_29_ & n67185;
  assign n67187 = P2_P3_REIP_REG_29_ & ~n67185;
  assign n67188 = ~n67186 & ~n67187;
  assign n67189 = n66404 & ~n67188;
  assign n67190 = P2_P3_EBX_REG_29_ & ~n66391;
  assign n67191 = n66393 & ~n67188;
  assign n67192 = P2_P3_EBX_REG_29_ & ~n67167;
  assign n67193 = ~P2_P3_EBX_REG_29_ & n67167;
  assign n67194 = ~n67192 & ~n67193;
  assign n67195 = n66395 & n67194;
  assign n67196 = ~n67191 & ~n67195;
  assign n67197 = ~n64472 & ~n67173;
  assign n67198 = n64472 & n67173;
  assign n67199 = ~n67197 & ~n67198;
  assign n67200 = n66413 & n67199;
  assign n67201 = P2_P3_REIP_REG_29_ & n66381;
  assign n67202 = P2_P3_PHYADDRPOINTER_REG_29_ & n66410;
  assign n67203 = ~n67201 & ~n67202;
  assign n67204 = ~n64472 & n66407;
  assign n67205 = n67203 & ~n67204;
  assign n67206 = ~n67189 & ~n67190;
  assign n67207 = n67196 & n67206;
  assign n67208 = ~n67200 & n67207;
  assign n12141 = ~n67205 | ~n67208;
  assign n67210 = P2_P3_REIP_REG_29_ & n67185;
  assign n67211 = ~P2_P3_REIP_REG_30_ & n67210;
  assign n67212 = P2_P3_REIP_REG_30_ & ~n67210;
  assign n67213 = ~n67211 & ~n67212;
  assign n67214 = n66404 & ~n67213;
  assign n67215 = P2_P3_EBX_REG_30_ & ~n66391;
  assign n67216 = n66393 & ~n67213;
  assign n67217 = ~P2_P3_EBX_REG_30_ & n67193;
  assign n67218 = P2_P3_EBX_REG_30_ & ~n67193;
  assign n67219 = ~n67217 & ~n67218;
  assign n67220 = n66395 & n67219;
  assign n67221 = ~n67216 & ~n67220;
  assign n67222 = n64495 & n67198;
  assign n67223 = ~n64495 & ~n67198;
  assign n67224 = ~n67222 & ~n67223;
  assign n67225 = n66413 & n67224;
  assign n67226 = P2_P3_REIP_REG_30_ & n66381;
  assign n67227 = P2_P3_PHYADDRPOINTER_REG_30_ & n66410;
  assign n67228 = ~n67226 & ~n67227;
  assign n67229 = ~n64495 & n66407;
  assign n67230 = n67228 & ~n67229;
  assign n67231 = ~n67214 & ~n67215;
  assign n67232 = n67221 & n67231;
  assign n67233 = ~n67225 & n67232;
  assign n12146 = ~n67230 | ~n67233;
  assign n67235 = ~n64518 & n67222;
  assign n67236 = n64518 & ~n67222;
  assign n67237 = ~n67235 & ~n67236;
  assign n67238 = ~n64518 & n66407;
  assign n67239 = n67237 & ~n67238;
  assign n67240 = P2_P3_EBX_REG_31_ & ~n66391;
  assign n67241 = P2_P3_EBX_REG_31_ & n67217;
  assign n67242 = ~P2_P3_EBX_REG_31_ & ~n67217;
  assign n67243 = ~n67241 & ~n67242;
  assign n67244 = n66395 & ~n67243;
  assign n67245 = P2_P3_REIP_REG_30_ & n67210;
  assign n67246 = ~P2_P3_REIP_REG_31_ & n67245;
  assign n67247 = P2_P3_REIP_REG_31_ & ~n67245;
  assign n67248 = ~n67246 & ~n67247;
  assign n67249 = n66393 & ~n67248;
  assign n67250 = P2_P3_PHYADDRPOINTER_REG_31_ & n66410;
  assign n67251 = P2_P3_REIP_REG_31_ & n66381;
  assign n67252 = ~n67250 & ~n67251;
  assign n67253 = n66404 & ~n67248;
  assign n67254 = n67252 & ~n67253;
  assign n67255 = ~n67240 & ~n67244;
  assign n67256 = ~n67249 & n67255;
  assign n67257 = n67254 & n67256;
  assign n67258 = n67239 & n67257;
  assign n67259 = ~n66413 & ~n67238;
  assign n67260 = n67257 & n67259;
  assign n12151 = ~n67258 & ~n67260;
  assign n67262 = ~P2_P3_DATAWIDTH_REG_1_ & ~P2_P3_REIP_REG_1_;
  assign n67263 = ~P2_P3_DATAWIDTH_REG_30_ & ~P2_P3_DATAWIDTH_REG_31_;
  assign n67264 = P2_P3_DATAWIDTH_REG_0_ & P2_P3_DATAWIDTH_REG_1_;
  assign n67265 = ~P2_P3_DATAWIDTH_REG_28_ & ~P2_P3_DATAWIDTH_REG_29_;
  assign n67266 = ~P2_P3_DATAWIDTH_REG_26_ & ~P2_P3_DATAWIDTH_REG_27_;
  assign n67267 = n67263 & ~n67264;
  assign n67268 = n67265 & n67267;
  assign n67269 = n67266 & n67268;
  assign n67270 = ~P2_P3_DATAWIDTH_REG_22_ & ~P2_P3_DATAWIDTH_REG_23_;
  assign n67271 = ~P2_P3_DATAWIDTH_REG_24_ & n67270;
  assign n67272 = ~P2_P3_DATAWIDTH_REG_25_ & n67271;
  assign n67273 = ~P2_P3_DATAWIDTH_REG_18_ & ~P2_P3_DATAWIDTH_REG_19_;
  assign n67274 = ~P2_P3_DATAWIDTH_REG_20_ & n67273;
  assign n67275 = ~P2_P3_DATAWIDTH_REG_21_ & n67274;
  assign n67276 = n67272 & n67275;
  assign n67277 = ~P2_P3_DATAWIDTH_REG_14_ & ~P2_P3_DATAWIDTH_REG_15_;
  assign n67278 = ~P2_P3_DATAWIDTH_REG_16_ & n67277;
  assign n67279 = ~P2_P3_DATAWIDTH_REG_17_ & n67278;
  assign n67280 = ~P2_P3_DATAWIDTH_REG_10_ & ~P2_P3_DATAWIDTH_REG_11_;
  assign n67281 = ~P2_P3_DATAWIDTH_REG_12_ & n67280;
  assign n67282 = ~P2_P3_DATAWIDTH_REG_13_ & n67281;
  assign n67283 = n67279 & n67282;
  assign n67284 = ~P2_P3_DATAWIDTH_REG_6_ & ~P2_P3_DATAWIDTH_REG_7_;
  assign n67285 = ~P2_P3_DATAWIDTH_REG_8_ & n67284;
  assign n67286 = ~P2_P3_DATAWIDTH_REG_9_ & n67285;
  assign n67287 = ~P2_P3_DATAWIDTH_REG_2_ & ~P2_P3_DATAWIDTH_REG_3_;
  assign n67288 = ~P2_P3_DATAWIDTH_REG_4_ & n67287;
  assign n67289 = ~P2_P3_DATAWIDTH_REG_5_ & n67288;
  assign n67290 = n67286 & n67289;
  assign n67291 = n67269 & n67276;
  assign n67292 = n67283 & n67291;
  assign n67293 = n67290 & n67292;
  assign n67294 = n67262 & n67293;
  assign n67295 = P2_P3_BYTEENABLE_REG_3_ & ~n67293;
  assign n67296 = ~P2_P3_DATAWIDTH_REG_0_ & ~P2_P3_REIP_REG_0_;
  assign n67297 = ~P2_P3_DATAWIDTH_REG_1_ & n67296;
  assign n67298 = n67293 & n67297;
  assign n67299 = ~n67294 & ~n67295;
  assign n12156 = n67298 | ~n67299;
  assign n67301 = P2_P3_REIP_REG_0_ & P2_P3_REIP_REG_1_;
  assign n67302 = P2_P3_DATAWIDTH_REG_0_ & ~P2_P3_REIP_REG_0_;
  assign n67303 = ~P2_P3_DATAWIDTH_REG_0_ & ~P2_P3_DATAWIDTH_REG_1_;
  assign n67304 = ~n67302 & ~n67303;
  assign n67305 = ~P2_P3_REIP_REG_1_ & ~n67304;
  assign n67306 = ~n67301 & ~n67305;
  assign n67307 = n67293 & ~n67306;
  assign n67308 = P2_P3_BYTEENABLE_REG_2_ & ~n67293;
  assign n12161 = n67307 | n67308;
  assign n67310 = P2_P3_REIP_REG_1_ & n67293;
  assign n67311 = P2_P3_BYTEENABLE_REG_1_ & ~n67293;
  assign n67312 = ~n67310 & ~n67311;
  assign n12166 = n67298 | ~n67312;
  assign n67314 = ~P2_P3_REIP_REG_0_ & ~P2_P3_REIP_REG_1_;
  assign n67315 = n67293 & ~n67314;
  assign n67316 = P2_P3_BYTEENABLE_REG_0_ & ~n67293;
  assign n12171 = n67315 | n67316;
  assign n67318 = P2_P3_W_R_N_REG & ~n58421;
  assign n67319 = ~P2_P3_READREQUEST_REG & n58421;
  assign n12176 = n67318 | n67319;
  assign n67321 = n59089 & n59321;
  assign n67322 = ~n59037 & n59321;
  assign n67323 = P2_P3_FLUSH_REG & ~n67322;
  assign n12181 = n67321 | n67323;
  assign n67325 = P2_P3_MORE_REG & ~n67322;
  assign n67326 = ~n59083 & n67322;
  assign n12186 = n67325 | n67326;
  assign n67328 = BS & ~n58642;
  assign n67329 = P2_P3_STATEBS16_REG & n58642;
  assign n67330 = ~P2_P3_STATE_REG_0_ & n58597;
  assign n67331 = ~n67328 & ~n67329;
  assign n12191 = n67330 | ~n67331;
  assign n67333 = ~n58967 & ~n59040;
  assign n67334 = ~n58685 & ~n67333;
  assign n67335 = ~P2_P3_STATEBS16_REG & n58967;
  assign n67336 = ~n58594 & ~n67335;
  assign n67337 = P2_P3_STATE2_REG_2_ & ~n67334;
  assign n67338 = n67336 & n67337;
  assign n67339 = P2_P3_STATE2_REG_0_ & ~n67338;
  assign n67340 = ~n59337 & ~n67339;
  assign n67341 = ~n58594 & n58679;
  assign n67342 = ~n59327 & ~n67341;
  assign n67343 = ~P2_P3_STATE2_REG_0_ & ~n67342;
  assign n67344 = ~n59399 & ~n67343;
  assign n67345 = ~n66380 & n67344;
  assign n67346 = ~n67340 & ~n67345;
  assign n67347 = P2_P3_REQUESTPENDING_REG & n67345;
  assign n12196 = n67346 | n67347;
  assign n67349 = P2_P3_D_C_N_REG & ~n58421;
  assign n67350 = ~P2_P3_CODEFETCH_REG & n58421;
  assign n67351 = ~n67349 & ~n67350;
  assign n12201 = n67330 | ~n67351;
  assign n67353 = P2_P3_MEMORYFETCH_REG & n58421;
  assign n67354 = P2_P3_M_IO_N_REG & ~n58421;
  assign n12206 = n67353 | n67354;
  assign n67356 = P2_P3_STATE2_REG_0_ & n60934;
  assign n67357 = n59036 & n59321;
  assign n67358 = P2_P3_CODEFETCH_REG & ~n67357;
  assign n12211 = n67356 | n67358;
  assign n67360 = P2_P3_STATE_REG_0_ & P2_P3_ADS_N_REG;
  assign n12216 = ~n58642 | n67360;
  assign n67362 = P2_P3_STATE2_REG_2_ & ~n59049;
  assign n67363 = ~n59044 & n67362;
  assign n67364 = ~n60934 & ~n66380;
  assign n67365 = ~n67363 & ~n67364;
  assign n67366 = P2_P3_READREQUEST_REG & n67364;
  assign n12221 = n67365 | n67366;
  assign n67368 = P2_P3_STATE2_REG_2_ & n58966;
  assign n67369 = ~n67364 & ~n67368;
  assign n67370 = P2_P3_MEMORYFETCH_REG & n67364;
  assign n12226 = n67369 | n67370;
  assign n67372 = P2_P2_STATE_REG_1_ & ~P2_P2_STATE_REG_0_;
  assign n67373 = P2_P2_BYTEENABLE_REG_3_ & n67372;
  assign n67374 = P2_P2_BE_N_REG_3_ & ~n67372;
  assign n12231 = n67373 | n67374;
  assign n67376 = P2_P2_BYTEENABLE_REG_2_ & n67372;
  assign n67377 = P2_P2_BE_N_REG_2_ & ~n67372;
  assign n12236 = n67376 | n67377;
  assign n67379 = P2_P2_BYTEENABLE_REG_1_ & n67372;
  assign n67380 = P2_P2_BE_N_REG_1_ & ~n67372;
  assign n12241 = n67379 | n67380;
  assign n67382 = P2_P2_BYTEENABLE_REG_0_ & n67372;
  assign n67383 = P2_P2_BE_N_REG_0_ & ~n67372;
  assign n12246 = n67382 | n67383;
  assign n67385 = P2_P2_STATE_REG_2_ & n67372;
  assign n67386 = P2_P2_REIP_REG_30_ & n67385;
  assign n67387 = ~P2_P2_STATE_REG_2_ & n67372;
  assign n67388 = P2_P2_REIP_REG_31_ & n67387;
  assign n67389 = P2_P2_ADDRESS_REG_29_ & ~n67372;
  assign n67390 = ~n67386 & ~n67388;
  assign n12251 = n67389 | ~n67390;
  assign n67392 = P2_P2_REIP_REG_29_ & n67385;
  assign n67393 = P2_P2_REIP_REG_30_ & n67387;
  assign n67394 = P2_P2_ADDRESS_REG_28_ & ~n67372;
  assign n67395 = ~n67392 & ~n67393;
  assign n12256 = n67394 | ~n67395;
  assign n67397 = P2_P2_REIP_REG_28_ & n67385;
  assign n67398 = P2_P2_REIP_REG_29_ & n67387;
  assign n67399 = P2_P2_ADDRESS_REG_27_ & ~n67372;
  assign n67400 = ~n67397 & ~n67398;
  assign n12261 = n67399 | ~n67400;
  assign n67402 = P2_P2_REIP_REG_27_ & n67385;
  assign n67403 = P2_P2_REIP_REG_28_ & n67387;
  assign n67404 = P2_P2_ADDRESS_REG_26_ & ~n67372;
  assign n67405 = ~n67402 & ~n67403;
  assign n12266 = n67404 | ~n67405;
  assign n67407 = P2_P2_REIP_REG_26_ & n67385;
  assign n67408 = P2_P2_REIP_REG_27_ & n67387;
  assign n67409 = P2_P2_ADDRESS_REG_25_ & ~n67372;
  assign n67410 = ~n67407 & ~n67408;
  assign n12271 = n67409 | ~n67410;
  assign n67412 = P2_P2_REIP_REG_25_ & n67385;
  assign n67413 = P2_P2_REIP_REG_26_ & n67387;
  assign n67414 = P2_P2_ADDRESS_REG_24_ & ~n67372;
  assign n67415 = ~n67412 & ~n67413;
  assign n12276 = n67414 | ~n67415;
  assign n67417 = P2_P2_REIP_REG_24_ & n67385;
  assign n67418 = P2_P2_REIP_REG_25_ & n67387;
  assign n67419 = P2_P2_ADDRESS_REG_23_ & ~n67372;
  assign n67420 = ~n67417 & ~n67418;
  assign n12281 = n67419 | ~n67420;
  assign n67422 = P2_P2_REIP_REG_23_ & n67385;
  assign n67423 = P2_P2_REIP_REG_24_ & n67387;
  assign n67424 = P2_P2_ADDRESS_REG_22_ & ~n67372;
  assign n67425 = ~n67422 & ~n67423;
  assign n12286 = n67424 | ~n67425;
  assign n67427 = P2_P2_REIP_REG_22_ & n67385;
  assign n67428 = P2_P2_REIP_REG_23_ & n67387;
  assign n67429 = P2_P2_ADDRESS_REG_21_ & ~n67372;
  assign n67430 = ~n67427 & ~n67428;
  assign n12291 = n67429 | ~n67430;
  assign n67432 = P2_P2_REIP_REG_21_ & n67385;
  assign n67433 = P2_P2_REIP_REG_22_ & n67387;
  assign n67434 = P2_P2_ADDRESS_REG_20_ & ~n67372;
  assign n67435 = ~n67432 & ~n67433;
  assign n12296 = n67434 | ~n67435;
  assign n67437 = P2_P2_REIP_REG_20_ & n67385;
  assign n67438 = P2_P2_REIP_REG_21_ & n67387;
  assign n67439 = P2_P2_ADDRESS_REG_19_ & ~n67372;
  assign n67440 = ~n67437 & ~n67438;
  assign n12301 = n67439 | ~n67440;
  assign n67442 = P2_P2_REIP_REG_19_ & n67385;
  assign n67443 = P2_P2_REIP_REG_20_ & n67387;
  assign n67444 = P2_P2_ADDRESS_REG_18_ & ~n67372;
  assign n67445 = ~n67442 & ~n67443;
  assign n12306 = n67444 | ~n67445;
  assign n67447 = P2_P2_REIP_REG_18_ & n67385;
  assign n67448 = P2_P2_REIP_REG_19_ & n67387;
  assign n67449 = P2_P2_ADDRESS_REG_17_ & ~n67372;
  assign n67450 = ~n67447 & ~n67448;
  assign n12311 = n67449 | ~n67450;
  assign n67452 = P2_P2_REIP_REG_17_ & n67385;
  assign n67453 = P2_P2_REIP_REG_18_ & n67387;
  assign n67454 = P2_P2_ADDRESS_REG_16_ & ~n67372;
  assign n67455 = ~n67452 & ~n67453;
  assign n12316 = n67454 | ~n67455;
  assign n67457 = P2_P2_REIP_REG_16_ & n67385;
  assign n67458 = P2_P2_REIP_REG_17_ & n67387;
  assign n67459 = P2_P2_ADDRESS_REG_15_ & ~n67372;
  assign n67460 = ~n67457 & ~n67458;
  assign n12321 = n67459 | ~n67460;
  assign n67462 = P2_P2_REIP_REG_15_ & n67385;
  assign n67463 = P2_P2_REIP_REG_16_ & n67387;
  assign n67464 = P2_P2_ADDRESS_REG_14_ & ~n67372;
  assign n67465 = ~n67462 & ~n67463;
  assign n12326 = n67464 | ~n67465;
  assign n67467 = P2_P2_REIP_REG_14_ & n67385;
  assign n67468 = P2_P2_REIP_REG_15_ & n67387;
  assign n67469 = P2_P2_ADDRESS_REG_13_ & ~n67372;
  assign n67470 = ~n67467 & ~n67468;
  assign n12331 = n67469 | ~n67470;
  assign n67472 = P2_P2_REIP_REG_13_ & n67385;
  assign n67473 = P2_P2_REIP_REG_14_ & n67387;
  assign n67474 = P2_P2_ADDRESS_REG_12_ & ~n67372;
  assign n67475 = ~n67472 & ~n67473;
  assign n12336 = n67474 | ~n67475;
  assign n67477 = P2_P2_REIP_REG_12_ & n67385;
  assign n67478 = P2_P2_REIP_REG_13_ & n67387;
  assign n67479 = P2_P2_ADDRESS_REG_11_ & ~n67372;
  assign n67480 = ~n67477 & ~n67478;
  assign n12341 = n67479 | ~n67480;
  assign n67482 = P2_P2_REIP_REG_11_ & n67385;
  assign n67483 = P2_P2_REIP_REG_12_ & n67387;
  assign n67484 = P2_P2_ADDRESS_REG_10_ & ~n67372;
  assign n67485 = ~n67482 & ~n67483;
  assign n12346 = n67484 | ~n67485;
  assign n67487 = P2_P2_REIP_REG_10_ & n67385;
  assign n67488 = P2_P2_REIP_REG_11_ & n67387;
  assign n67489 = P2_P2_ADDRESS_REG_9_ & ~n67372;
  assign n67490 = ~n67487 & ~n67488;
  assign n12351 = n67489 | ~n67490;
  assign n67492 = P2_P2_REIP_REG_9_ & n67385;
  assign n67493 = P2_P2_REIP_REG_10_ & n67387;
  assign n67494 = P2_P2_ADDRESS_REG_8_ & ~n67372;
  assign n67495 = ~n67492 & ~n67493;
  assign n12356 = n67494 | ~n67495;
  assign n67497 = P2_P2_REIP_REG_8_ & n67385;
  assign n67498 = P2_P2_REIP_REG_9_ & n67387;
  assign n67499 = P2_P2_ADDRESS_REG_7_ & ~n67372;
  assign n67500 = ~n67497 & ~n67498;
  assign n12361 = n67499 | ~n67500;
  assign n67502 = P2_P2_REIP_REG_7_ & n67385;
  assign n67503 = P2_P2_REIP_REG_8_ & n67387;
  assign n67504 = P2_P2_ADDRESS_REG_6_ & ~n67372;
  assign n67505 = ~n67502 & ~n67503;
  assign n12366 = n67504 | ~n67505;
  assign n67507 = P2_P2_REIP_REG_6_ & n67385;
  assign n67508 = P2_P2_REIP_REG_7_ & n67387;
  assign n67509 = P2_P2_ADDRESS_REG_5_ & ~n67372;
  assign n67510 = ~n67507 & ~n67508;
  assign n12371 = n67509 | ~n67510;
  assign n67512 = P2_P2_REIP_REG_5_ & n67385;
  assign n67513 = P2_P2_REIP_REG_6_ & n67387;
  assign n67514 = P2_P2_ADDRESS_REG_4_ & ~n67372;
  assign n67515 = ~n67512 & ~n67513;
  assign n12376 = n67514 | ~n67515;
  assign n67517 = P2_P2_REIP_REG_4_ & n67385;
  assign n67518 = P2_P2_REIP_REG_5_ & n67387;
  assign n67519 = P2_P2_ADDRESS_REG_3_ & ~n67372;
  assign n67520 = ~n67517 & ~n67518;
  assign n12381 = n67519 | ~n67520;
  assign n67522 = P2_P2_REIP_REG_3_ & n67385;
  assign n67523 = P2_P2_REIP_REG_4_ & n67387;
  assign n67524 = P2_P2_ADDRESS_REG_2_ & ~n67372;
  assign n67525 = ~n67522 & ~n67523;
  assign n12386 = n67524 | ~n67525;
  assign n67527 = P2_P2_REIP_REG_2_ & n67385;
  assign n67528 = P2_P2_REIP_REG_3_ & n67387;
  assign n67529 = P2_P2_ADDRESS_REG_1_ & ~n67372;
  assign n67530 = ~n67527 & ~n67528;
  assign n12391 = n67529 | ~n67530;
  assign n67532 = P2_P2_REIP_REG_1_ & n67385;
  assign n67533 = P2_P2_REIP_REG_2_ & n67387;
  assign n67534 = P2_P2_ADDRESS_REG_0_ & ~n67372;
  assign n67535 = ~n67532 & ~n67533;
  assign n12396 = n67534 | ~n67535;
  assign n67537 = ~P2_P2_STATE_REG_2_ & P2_P2_STATE_REG_1_;
  assign n67538 = NA & n67537;
  assign n67539 = P2_P2_STATE_REG_0_ & ~n67538;
  assign n67540 = ~HOLD & ~P2_P2_REQUESTPENDING_REG;
  assign n67541 = P2_READY12_REG & P2_READY21_REG;
  assign n67542 = ~n67540 & n67541;
  assign n67543 = n67537 & n67542;
  assign n67544 = ~P2_P2_STATE_REG_2_ & ~P2_P2_STATE_REG_1_;
  assign n67545 = HOLD & ~P2_P2_REQUESTPENDING_REG;
  assign n67546 = n67544 & n67545;
  assign n67547 = ~n67543 & ~n67546;
  assign n67548 = n67539 & ~n67547;
  assign n67549 = ~n67385 & ~n67548;
  assign n67550 = ~HOLD & P2_P2_REQUESTPENDING_REG;
  assign n67551 = P2_P2_STATE_REG_0_ & ~n67550;
  assign n67552 = ~n67540 & n67551;
  assign n67553 = ~NA & ~P2_P2_STATE_REG_0_;
  assign n67554 = n67540 & ~n67541;
  assign n67555 = ~n67541 & n67550;
  assign n67556 = P2_P2_STATE_REG_1_ & ~n67554;
  assign n67557 = ~n67555 & n67556;
  assign n67558 = ~n67552 & ~n67553;
  assign n67559 = ~n67557 & n67558;
  assign n67560 = P2_P2_STATE_REG_2_ & ~n67559;
  assign n12401 = ~n67549 | n67560;
  assign n67562 = P2_P2_STATE_REG_2_ & ~n67551;
  assign n67563 = P2_P2_STATE_REG_0_ & P2_P2_REQUESTPENDING_REG;
  assign n67564 = ~P2_P2_STATE_REG_2_ & n67563;
  assign n67565 = ~n67562 & ~n67564;
  assign n67566 = ~P2_P2_STATE_REG_1_ & ~n67565;
  assign n67567 = HOLD & ~n67541;
  assign n67568 = P2_P2_STATE_REG_0_ & ~n67567;
  assign n67569 = P2_P2_STATE_REG_2_ & ~n67568;
  assign n67570 = ~n67554 & ~n67569;
  assign n67571 = P2_P2_STATE_REG_1_ & n67570;
  assign n67572 = n67372 & n67541;
  assign n67573 = ~n67387 & ~n67572;
  assign n67574 = ~n67566 & ~n67571;
  assign n12406 = ~n67573 | ~n67574;
  assign n67576 = P2_P2_STATE_REG_1_ & ~n67555;
  assign n67577 = n67563 & ~n67576;
  assign n67578 = ~P2_P2_STATE_REG_2_ & ~n67577;
  assign n67579 = P2_P2_STATE_REG_2_ & n67551;
  assign n67580 = NA & ~P2_P2_STATE_REG_0_;
  assign n67581 = P2_P2_STATE_REG_2_ & ~n67550;
  assign n67582 = ~n67580 & ~n67581;
  assign n67583 = ~P2_P2_STATE_REG_1_ & ~n67582;
  assign n67584 = ~n67578 & ~n67579;
  assign n12411 = n67583 | ~n67584;
  assign n67586 = ~BS & ~n67544;
  assign n67587 = P2_P2_STATE_REG_0_ & n67537;
  assign n67588 = ~P2_P2_STATE_REG_1_ & ~P2_P2_STATE_REG_0_;
  assign n67589 = ~n67587 & ~n67588;
  assign n67590 = n67586 & ~n67589;
  assign n67591 = P2_P2_DATAWIDTH_REG_0_ & n67589;
  assign n12416 = n67590 | n67591;
  assign n67593 = P2_P2_DATAWIDTH_REG_1_ & n67589;
  assign n67594 = ~n67586 & ~n67589;
  assign n12421 = n67593 | n67594;
  assign n12426 = P2_P2_DATAWIDTH_REG_2_ & n67589;
  assign n12431 = P2_P2_DATAWIDTH_REG_3_ & n67589;
  assign n12436 = P2_P2_DATAWIDTH_REG_4_ & n67589;
  assign n12441 = P2_P2_DATAWIDTH_REG_5_ & n67589;
  assign n12446 = P2_P2_DATAWIDTH_REG_6_ & n67589;
  assign n12451 = P2_P2_DATAWIDTH_REG_7_ & n67589;
  assign n12456 = P2_P2_DATAWIDTH_REG_8_ & n67589;
  assign n12461 = P2_P2_DATAWIDTH_REG_9_ & n67589;
  assign n12466 = P2_P2_DATAWIDTH_REG_10_ & n67589;
  assign n12471 = P2_P2_DATAWIDTH_REG_11_ & n67589;
  assign n12476 = P2_P2_DATAWIDTH_REG_12_ & n67589;
  assign n12481 = P2_P2_DATAWIDTH_REG_13_ & n67589;
  assign n12486 = P2_P2_DATAWIDTH_REG_14_ & n67589;
  assign n12491 = P2_P2_DATAWIDTH_REG_15_ & n67589;
  assign n12496 = P2_P2_DATAWIDTH_REG_16_ & n67589;
  assign n12501 = P2_P2_DATAWIDTH_REG_17_ & n67589;
  assign n12506 = P2_P2_DATAWIDTH_REG_18_ & n67589;
  assign n12511 = P2_P2_DATAWIDTH_REG_19_ & n67589;
  assign n12516 = P2_P2_DATAWIDTH_REG_20_ & n67589;
  assign n12521 = P2_P2_DATAWIDTH_REG_21_ & n67589;
  assign n12526 = P2_P2_DATAWIDTH_REG_22_ & n67589;
  assign n12531 = P2_P2_DATAWIDTH_REG_23_ & n67589;
  assign n12536 = P2_P2_DATAWIDTH_REG_24_ & n67589;
  assign n12541 = P2_P2_DATAWIDTH_REG_25_ & n67589;
  assign n12546 = P2_P2_DATAWIDTH_REG_26_ & n67589;
  assign n12551 = P2_P2_DATAWIDTH_REG_27_ & n67589;
  assign n12556 = P2_P2_DATAWIDTH_REG_28_ & n67589;
  assign n12561 = P2_P2_DATAWIDTH_REG_29_ & n67589;
  assign n12566 = P2_P2_DATAWIDTH_REG_30_ & n67589;
  assign n12571 = P2_P2_DATAWIDTH_REG_31_ & n67589;
  assign n67626 = P2_P2_STATE2_REG_2_ & P2_P2_STATE2_REG_1_;
  assign n67627 = P2_P2_STATE2_REG_1_ & n67541;
  assign n67628 = ~P2_P2_STATE2_REG_0_ & ~n67627;
  assign n67629 = ~P2_P2_STATEBS16_REG & ~n67541;
  assign n67630 = P2_P2_STATE_REG_2_ & ~P2_P2_STATE_REG_1_;
  assign n67631 = ~n67537 & ~n67630;
  assign n67632 = ~P2_P2_STATE_REG_0_ & ~n67631;
  assign n67633 = n67629 & n67632;
  assign n67634 = P2_P2_INSTQUEUERD_ADDR_REG_1_ & P2_P2_INSTQUEUERD_ADDR_REG_0_;
  assign n67635 = ~P2_P2_INSTQUEUERD_ADDR_REG_2_ & n67634;
  assign n67636 = P2_P2_INSTQUEUERD_ADDR_REG_3_ & n67635;
  assign n67637 = P2_P2_INSTQUEUE_REG_11__5_ & n67636;
  assign n67638 = P2_P2_INSTQUEUERD_ADDR_REG_1_ & ~P2_P2_INSTQUEUERD_ADDR_REG_0_;
  assign n67639 = ~P2_P2_INSTQUEUERD_ADDR_REG_2_ & n67638;
  assign n67640 = P2_P2_INSTQUEUERD_ADDR_REG_3_ & n67639;
  assign n67641 = P2_P2_INSTQUEUE_REG_10__5_ & n67640;
  assign n67642 = ~n67637 & ~n67641;
  assign n67643 = ~P2_P2_INSTQUEUERD_ADDR_REG_1_ & P2_P2_INSTQUEUERD_ADDR_REG_0_;
  assign n67644 = ~P2_P2_INSTQUEUERD_ADDR_REG_2_ & n67643;
  assign n67645 = P2_P2_INSTQUEUERD_ADDR_REG_3_ & n67644;
  assign n67646 = P2_P2_INSTQUEUE_REG_9__5_ & n67645;
  assign n67647 = ~P2_P2_INSTQUEUERD_ADDR_REG_1_ & ~P2_P2_INSTQUEUERD_ADDR_REG_0_;
  assign n67648 = ~P2_P2_INSTQUEUERD_ADDR_REG_2_ & n67647;
  assign n67649 = P2_P2_INSTQUEUERD_ADDR_REG_3_ & n67648;
  assign n67650 = P2_P2_INSTQUEUE_REG_8__5_ & n67649;
  assign n67651 = ~n67646 & ~n67650;
  assign n67652 = P2_P2_INSTQUEUERD_ADDR_REG_3_ & P2_P2_INSTQUEUERD_ADDR_REG_2_;
  assign n67653 = n67634 & n67652;
  assign n67654 = P2_P2_INSTQUEUE_REG_15__5_ & n67653;
  assign n67655 = n67638 & n67652;
  assign n67656 = P2_P2_INSTQUEUE_REG_14__5_ & n67655;
  assign n67657 = n67643 & n67652;
  assign n67658 = P2_P2_INSTQUEUE_REG_13__5_ & n67657;
  assign n67659 = n67647 & n67652;
  assign n67660 = P2_P2_INSTQUEUE_REG_12__5_ & n67659;
  assign n67661 = ~n67654 & ~n67656;
  assign n67662 = ~n67658 & n67661;
  assign n67663 = ~n67660 & n67662;
  assign n67664 = ~P2_P2_INSTQUEUERD_ADDR_REG_3_ & P2_P2_INSTQUEUERD_ADDR_REG_2_;
  assign n67665 = n67634 & n67664;
  assign n67666 = P2_P2_INSTQUEUE_REG_7__5_ & n67665;
  assign n67667 = n67638 & n67664;
  assign n67668 = P2_P2_INSTQUEUE_REG_6__5_ & n67667;
  assign n67669 = n67643 & n67664;
  assign n67670 = P2_P2_INSTQUEUE_REG_5__5_ & n67669;
  assign n67671 = n67647 & n67664;
  assign n67672 = P2_P2_INSTQUEUE_REG_4__5_ & n67671;
  assign n67673 = ~n67666 & ~n67668;
  assign n67674 = ~n67670 & n67673;
  assign n67675 = ~n67672 & n67674;
  assign n67676 = ~P2_P2_INSTQUEUERD_ADDR_REG_3_ & n67635;
  assign n67677 = P2_P2_INSTQUEUE_REG_3__5_ & n67676;
  assign n67678 = ~P2_P2_INSTQUEUERD_ADDR_REG_3_ & ~P2_P2_INSTQUEUERD_ADDR_REG_2_;
  assign n67679 = n67638 & n67678;
  assign n67680 = P2_P2_INSTQUEUE_REG_2__5_ & n67679;
  assign n67681 = n67643 & n67678;
  assign n67682 = P2_P2_INSTQUEUE_REG_1__5_ & n67681;
  assign n67683 = ~P2_P2_INSTQUEUERD_ADDR_REG_3_ & n67648;
  assign n67684 = P2_P2_INSTQUEUE_REG_0__5_ & n67683;
  assign n67685 = ~n67677 & ~n67680;
  assign n67686 = ~n67682 & n67685;
  assign n67687 = ~n67684 & n67686;
  assign n67688 = n67642 & n67651;
  assign n67689 = n67663 & n67688;
  assign n67690 = n67675 & n67689;
  assign n67691 = n67687 & n67690;
  assign n67692 = P2_P2_INSTQUEUE_REG_11__6_ & n67636;
  assign n67693 = P2_P2_INSTQUEUE_REG_10__6_ & n67640;
  assign n67694 = ~n67692 & ~n67693;
  assign n67695 = P2_P2_INSTQUEUE_REG_9__6_ & n67645;
  assign n67696 = P2_P2_INSTQUEUE_REG_8__6_ & n67649;
  assign n67697 = ~n67695 & ~n67696;
  assign n67698 = P2_P2_INSTQUEUE_REG_15__6_ & n67653;
  assign n67699 = P2_P2_INSTQUEUE_REG_14__6_ & n67655;
  assign n67700 = P2_P2_INSTQUEUE_REG_13__6_ & n67657;
  assign n67701 = P2_P2_INSTQUEUE_REG_12__6_ & n67659;
  assign n67702 = ~n67698 & ~n67699;
  assign n67703 = ~n67700 & n67702;
  assign n67704 = ~n67701 & n67703;
  assign n67705 = P2_P2_INSTQUEUE_REG_7__6_ & n67665;
  assign n67706 = P2_P2_INSTQUEUE_REG_6__6_ & n67667;
  assign n67707 = P2_P2_INSTQUEUE_REG_5__6_ & n67669;
  assign n67708 = P2_P2_INSTQUEUE_REG_4__6_ & n67671;
  assign n67709 = ~n67705 & ~n67706;
  assign n67710 = ~n67707 & n67709;
  assign n67711 = ~n67708 & n67710;
  assign n67712 = P2_P2_INSTQUEUE_REG_3__6_ & n67676;
  assign n67713 = P2_P2_INSTQUEUE_REG_2__6_ & n67679;
  assign n67714 = P2_P2_INSTQUEUE_REG_1__6_ & n67681;
  assign n67715 = P2_P2_INSTQUEUE_REG_0__6_ & n67683;
  assign n67716 = ~n67712 & ~n67713;
  assign n67717 = ~n67714 & n67716;
  assign n67718 = ~n67715 & n67717;
  assign n67719 = n67694 & n67697;
  assign n67720 = n67704 & n67719;
  assign n67721 = n67711 & n67720;
  assign n67722 = n67718 & n67721;
  assign n67723 = n67691 & n67722;
  assign n67724 = P2_P2_INSTQUEUE_REG_11__4_ & n67636;
  assign n67725 = P2_P2_INSTQUEUE_REG_10__4_ & n67640;
  assign n67726 = ~n67724 & ~n67725;
  assign n67727 = P2_P2_INSTQUEUE_REG_9__4_ & n67645;
  assign n67728 = P2_P2_INSTQUEUE_REG_8__4_ & n67649;
  assign n67729 = ~n67727 & ~n67728;
  assign n67730 = P2_P2_INSTQUEUE_REG_15__4_ & n67653;
  assign n67731 = P2_P2_INSTQUEUE_REG_14__4_ & n67655;
  assign n67732 = P2_P2_INSTQUEUE_REG_13__4_ & n67657;
  assign n67733 = P2_P2_INSTQUEUE_REG_12__4_ & n67659;
  assign n67734 = ~n67730 & ~n67731;
  assign n67735 = ~n67732 & n67734;
  assign n67736 = ~n67733 & n67735;
  assign n67737 = P2_P2_INSTQUEUE_REG_7__4_ & n67665;
  assign n67738 = P2_P2_INSTQUEUE_REG_6__4_ & n67667;
  assign n67739 = P2_P2_INSTQUEUE_REG_5__4_ & n67669;
  assign n67740 = P2_P2_INSTQUEUE_REG_4__4_ & n67671;
  assign n67741 = ~n67737 & ~n67738;
  assign n67742 = ~n67739 & n67741;
  assign n67743 = ~n67740 & n67742;
  assign n67744 = P2_P2_INSTQUEUE_REG_3__4_ & n67676;
  assign n67745 = P2_P2_INSTQUEUE_REG_2__4_ & n67679;
  assign n67746 = P2_P2_INSTQUEUE_REG_1__4_ & n67681;
  assign n67747 = P2_P2_INSTQUEUE_REG_0__4_ & n67683;
  assign n67748 = ~n67744 & ~n67745;
  assign n67749 = ~n67746 & n67748;
  assign n67750 = ~n67747 & n67749;
  assign n67751 = n67726 & n67729;
  assign n67752 = n67736 & n67751;
  assign n67753 = n67743 & n67752;
  assign n67754 = n67750 & n67753;
  assign n67755 = P2_P2_INSTQUEUE_REG_11__7_ & n67636;
  assign n67756 = P2_P2_INSTQUEUE_REG_10__7_ & n67640;
  assign n67757 = ~n67755 & ~n67756;
  assign n67758 = P2_P2_INSTQUEUE_REG_9__7_ & n67645;
  assign n67759 = P2_P2_INSTQUEUE_REG_8__7_ & n67649;
  assign n67760 = ~n67758 & ~n67759;
  assign n67761 = P2_P2_INSTQUEUE_REG_15__7_ & n67653;
  assign n67762 = P2_P2_INSTQUEUE_REG_14__7_ & n67655;
  assign n67763 = P2_P2_INSTQUEUE_REG_13__7_ & n67657;
  assign n67764 = P2_P2_INSTQUEUE_REG_12__7_ & n67659;
  assign n67765 = ~n67761 & ~n67762;
  assign n67766 = ~n67763 & n67765;
  assign n67767 = ~n67764 & n67766;
  assign n67768 = P2_P2_INSTQUEUE_REG_7__7_ & n67665;
  assign n67769 = P2_P2_INSTQUEUE_REG_6__7_ & n67667;
  assign n67770 = P2_P2_INSTQUEUE_REG_5__7_ & n67669;
  assign n67771 = P2_P2_INSTQUEUE_REG_4__7_ & n67671;
  assign n67772 = ~n67768 & ~n67769;
  assign n67773 = ~n67770 & n67772;
  assign n67774 = ~n67771 & n67773;
  assign n67775 = P2_P2_INSTQUEUE_REG_3__7_ & n67676;
  assign n67776 = P2_P2_INSTQUEUE_REG_2__7_ & n67679;
  assign n67777 = P2_P2_INSTQUEUE_REG_1__7_ & n67681;
  assign n67778 = P2_P2_INSTQUEUE_REG_0__7_ & n67683;
  assign n67779 = ~n67775 & ~n67776;
  assign n67780 = ~n67777 & n67779;
  assign n67781 = ~n67778 & n67780;
  assign n67782 = n67757 & n67760;
  assign n67783 = n67767 & n67782;
  assign n67784 = n67774 & n67783;
  assign n67785 = n67781 & n67784;
  assign n67786 = P2_P2_INSTQUEUE_REG_11__3_ & n67636;
  assign n67787 = P2_P2_INSTQUEUE_REG_10__3_ & n67640;
  assign n67788 = ~n67786 & ~n67787;
  assign n67789 = P2_P2_INSTQUEUE_REG_9__3_ & n67645;
  assign n67790 = P2_P2_INSTQUEUE_REG_8__3_ & n67649;
  assign n67791 = ~n67789 & ~n67790;
  assign n67792 = P2_P2_INSTQUEUE_REG_15__3_ & n67653;
  assign n67793 = P2_P2_INSTQUEUE_REG_14__3_ & n67655;
  assign n67794 = P2_P2_INSTQUEUE_REG_13__3_ & n67657;
  assign n67795 = P2_P2_INSTQUEUE_REG_12__3_ & n67659;
  assign n67796 = ~n67792 & ~n67793;
  assign n67797 = ~n67794 & n67796;
  assign n67798 = ~n67795 & n67797;
  assign n67799 = P2_P2_INSTQUEUE_REG_7__3_ & n67665;
  assign n67800 = P2_P2_INSTQUEUE_REG_6__3_ & n67667;
  assign n67801 = P2_P2_INSTQUEUE_REG_5__3_ & n67669;
  assign n67802 = P2_P2_INSTQUEUE_REG_4__3_ & n67671;
  assign n67803 = ~n67799 & ~n67800;
  assign n67804 = ~n67801 & n67803;
  assign n67805 = ~n67802 & n67804;
  assign n67806 = P2_P2_INSTQUEUE_REG_3__3_ & n67676;
  assign n67807 = P2_P2_INSTQUEUE_REG_2__3_ & n67679;
  assign n67808 = P2_P2_INSTQUEUE_REG_1__3_ & n67681;
  assign n67809 = P2_P2_INSTQUEUE_REG_0__3_ & n67683;
  assign n67810 = ~n67806 & ~n67807;
  assign n67811 = ~n67808 & n67810;
  assign n67812 = ~n67809 & n67811;
  assign n67813 = n67788 & n67791;
  assign n67814 = n67798 & n67813;
  assign n67815 = n67805 & n67814;
  assign n67816 = n67812 & n67815;
  assign n67817 = P2_P2_INSTQUEUE_REG_11__2_ & n67636;
  assign n67818 = P2_P2_INSTQUEUE_REG_10__2_ & n67640;
  assign n67819 = ~n67817 & ~n67818;
  assign n67820 = P2_P2_INSTQUEUE_REG_9__2_ & n67645;
  assign n67821 = P2_P2_INSTQUEUE_REG_8__2_ & n67649;
  assign n67822 = ~n67820 & ~n67821;
  assign n67823 = P2_P2_INSTQUEUE_REG_15__2_ & n67653;
  assign n67824 = P2_P2_INSTQUEUE_REG_14__2_ & n67655;
  assign n67825 = P2_P2_INSTQUEUE_REG_13__2_ & n67657;
  assign n67826 = P2_P2_INSTQUEUE_REG_12__2_ & n67659;
  assign n67827 = ~n67823 & ~n67824;
  assign n67828 = ~n67825 & n67827;
  assign n67829 = ~n67826 & n67828;
  assign n67830 = P2_P2_INSTQUEUE_REG_7__2_ & n67665;
  assign n67831 = P2_P2_INSTQUEUE_REG_6__2_ & n67667;
  assign n67832 = P2_P2_INSTQUEUE_REG_5__2_ & n67669;
  assign n67833 = P2_P2_INSTQUEUE_REG_4__2_ & n67671;
  assign n67834 = ~n67830 & ~n67831;
  assign n67835 = ~n67832 & n67834;
  assign n67836 = ~n67833 & n67835;
  assign n67837 = P2_P2_INSTQUEUE_REG_3__2_ & n67676;
  assign n67838 = P2_P2_INSTQUEUE_REG_2__2_ & n67679;
  assign n67839 = P2_P2_INSTQUEUE_REG_1__2_ & n67681;
  assign n67840 = P2_P2_INSTQUEUE_REG_0__2_ & n67683;
  assign n67841 = ~n67837 & ~n67838;
  assign n67842 = ~n67839 & n67841;
  assign n67843 = ~n67840 & n67842;
  assign n67844 = n67819 & n67822;
  assign n67845 = n67829 & n67844;
  assign n67846 = n67836 & n67845;
  assign n67847 = n67843 & n67846;
  assign n67848 = ~n67785 & ~n67816;
  assign n67849 = n67847 & n67848;
  assign n67850 = n67723 & n67754;
  assign n67851 = n67849 & n67850;
  assign n67852 = P2_P2_INSTQUEUE_REG_11__1_ & n67636;
  assign n67853 = P2_P2_INSTQUEUE_REG_10__1_ & n67640;
  assign n67854 = ~n67852 & ~n67853;
  assign n67855 = P2_P2_INSTQUEUE_REG_9__1_ & n67645;
  assign n67856 = P2_P2_INSTQUEUE_REG_8__1_ & n67649;
  assign n67857 = ~n67855 & ~n67856;
  assign n67858 = P2_P2_INSTQUEUE_REG_15__1_ & n67653;
  assign n67859 = P2_P2_INSTQUEUE_REG_14__1_ & n67655;
  assign n67860 = P2_P2_INSTQUEUE_REG_13__1_ & n67657;
  assign n67861 = P2_P2_INSTQUEUE_REG_12__1_ & n67659;
  assign n67862 = ~n67858 & ~n67859;
  assign n67863 = ~n67860 & n67862;
  assign n67864 = ~n67861 & n67863;
  assign n67865 = P2_P2_INSTQUEUE_REG_7__1_ & n67665;
  assign n67866 = P2_P2_INSTQUEUE_REG_6__1_ & n67667;
  assign n67867 = P2_P2_INSTQUEUE_REG_5__1_ & n67669;
  assign n67868 = P2_P2_INSTQUEUE_REG_4__1_ & n67671;
  assign n67869 = ~n67865 & ~n67866;
  assign n67870 = ~n67867 & n67869;
  assign n67871 = ~n67868 & n67870;
  assign n67872 = P2_P2_INSTQUEUE_REG_3__1_ & n67676;
  assign n67873 = P2_P2_INSTQUEUE_REG_2__1_ & n67679;
  assign n67874 = P2_P2_INSTQUEUE_REG_1__1_ & n67681;
  assign n67875 = P2_P2_INSTQUEUE_REG_0__1_ & n67683;
  assign n67876 = ~n67872 & ~n67873;
  assign n67877 = ~n67874 & n67876;
  assign n67878 = ~n67875 & n67877;
  assign n67879 = n67854 & n67857;
  assign n67880 = n67864 & n67879;
  assign n67881 = n67871 & n67880;
  assign n67882 = n67878 & n67881;
  assign n67883 = P2_P2_INSTQUEUE_REG_11__0_ & n67636;
  assign n67884 = P2_P2_INSTQUEUE_REG_10__0_ & n67640;
  assign n67885 = ~n67883 & ~n67884;
  assign n67886 = P2_P2_INSTQUEUE_REG_9__0_ & n67645;
  assign n67887 = P2_P2_INSTQUEUE_REG_8__0_ & n67649;
  assign n67888 = ~n67886 & ~n67887;
  assign n67889 = P2_P2_INSTQUEUE_REG_15__0_ & n67653;
  assign n67890 = P2_P2_INSTQUEUE_REG_14__0_ & n67655;
  assign n67891 = P2_P2_INSTQUEUE_REG_13__0_ & n67657;
  assign n67892 = P2_P2_INSTQUEUE_REG_12__0_ & n67659;
  assign n67893 = ~n67889 & ~n67890;
  assign n67894 = ~n67891 & n67893;
  assign n67895 = ~n67892 & n67894;
  assign n67896 = P2_P2_INSTQUEUE_REG_7__0_ & n67665;
  assign n67897 = P2_P2_INSTQUEUE_REG_6__0_ & n67667;
  assign n67898 = P2_P2_INSTQUEUE_REG_5__0_ & n67669;
  assign n67899 = P2_P2_INSTQUEUE_REG_4__0_ & n67671;
  assign n67900 = ~n67896 & ~n67897;
  assign n67901 = ~n67898 & n67900;
  assign n67902 = ~n67899 & n67901;
  assign n67903 = P2_P2_INSTQUEUE_REG_3__0_ & n67676;
  assign n67904 = P2_P2_INSTQUEUE_REG_2__0_ & n67679;
  assign n67905 = P2_P2_INSTQUEUE_REG_1__0_ & n67681;
  assign n67906 = P2_P2_INSTQUEUE_REG_0__0_ & n67683;
  assign n67907 = ~n67903 & ~n67904;
  assign n67908 = ~n67905 & n67907;
  assign n67909 = ~n67906 & n67908;
  assign n67910 = n67885 & n67888;
  assign n67911 = n67895 & n67910;
  assign n67912 = n67902 & n67911;
  assign n67913 = n67909 & n67912;
  assign n67914 = n67882 & ~n67913;
  assign n67915 = n67851 & n67914;
  assign n67916 = n67633 & n67915;
  assign n67917 = ~P2_P2_STATE2_REG_1_ & ~n67916;
  assign n67918 = ~n67541 & n67632;
  assign n67919 = ~n67847 & ~n67882;
  assign n67920 = n67918 & n67919;
  assign n67921 = ~n67541 & ~n67847;
  assign n67922 = n67882 & n67921;
  assign n67923 = ~n67541 & n67847;
  assign n67924 = n67882 & ~n67918;
  assign n67925 = n67923 & ~n67924;
  assign n67926 = ~n67920 & ~n67922;
  assign n67927 = ~n67925 & n67926;
  assign n67928 = P2_P2_INSTQUEUERD_ADDR_REG_4_ & ~P2_P2_INSTQUEUEWR_ADDR_REG_4_;
  assign n67929 = ~P2_P2_INSTQUEUERD_ADDR_REG_3_ & P2_P2_INSTQUEUEWR_ADDR_REG_3_;
  assign n67930 = P2_P2_INSTQUEUERD_ADDR_REG_3_ & ~P2_P2_INSTQUEUEWR_ADDR_REG_3_;
  assign n67931 = ~P2_P2_INSTQUEUERD_ADDR_REG_2_ & P2_P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n67932 = P2_P2_INSTQUEUERD_ADDR_REG_2_ & ~P2_P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n67933 = P2_P2_INSTQUEUERD_ADDR_REG_0_ & ~P2_P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n67934 = P2_P2_INSTQUEUEWR_ADDR_REG_1_ & ~n67933;
  assign n67935 = ~P2_P2_INSTQUEUEWR_ADDR_REG_1_ & n67933;
  assign n67936 = ~P2_P2_INSTQUEUERD_ADDR_REG_1_ & ~n67935;
  assign n67937 = ~n67934 & ~n67936;
  assign n67938 = ~n67932 & ~n67937;
  assign n67939 = ~n67931 & ~n67938;
  assign n67940 = ~n67930 & ~n67939;
  assign n67941 = ~n67929 & ~n67940;
  assign n67942 = ~P2_P2_INSTQUEUERD_ADDR_REG_4_ & P2_P2_INSTQUEUEWR_ADDR_REG_4_;
  assign n67943 = n67941 & ~n67942;
  assign n67944 = ~n67928 & ~n67943;
  assign n67945 = ~n67928 & ~n67942;
  assign n67946 = ~n67941 & ~n67945;
  assign n67947 = n67941 & n67945;
  assign n67948 = ~n67946 & ~n67947;
  assign n67949 = ~n67929 & ~n67930;
  assign n67950 = ~n67939 & ~n67949;
  assign n67951 = n67939 & n67949;
  assign n67952 = ~n67950 & ~n67951;
  assign n67953 = ~P2_P2_INSTQUEUERD_ADDR_REG_1_ & P2_P2_INSTQUEUEWR_ADDR_REG_1_;
  assign n67954 = P2_P2_INSTQUEUERD_ADDR_REG_1_ & ~P2_P2_INSTQUEUEWR_ADDR_REG_1_;
  assign n67955 = ~n67953 & ~n67954;
  assign n67956 = ~n67933 & ~n67955;
  assign n67957 = n67933 & n67955;
  assign n67958 = ~n67956 & ~n67957;
  assign n67959 = ~n67931 & ~n67932;
  assign n67960 = ~n67937 & ~n67959;
  assign n67961 = n67937 & n67959;
  assign n67962 = ~n67960 & ~n67961;
  assign n67963 = n67948 & n67952;
  assign n67964 = n67958 & n67963;
  assign n67965 = n67962 & n67964;
  assign n67966 = n67944 & ~n67965;
  assign n67967 = ~n67882 & ~n67966;
  assign n67968 = n67882 & ~n67966;
  assign n67969 = ~n67967 & ~n67968;
  assign n67970 = ~n67785 & n67816;
  assign n67971 = ~n67691 & ~n67722;
  assign n67972 = n67754 & n67971;
  assign n67973 = n67970 & n67972;
  assign n67974 = n67913 & n67973;
  assign n67975 = n67969 & n67974;
  assign n67976 = ~n67847 & ~n67975;
  assign n67977 = ~n67816 & ~n67913;
  assign n67978 = ~n67785 & n67977;
  assign n67979 = n67850 & n67978;
  assign n67980 = ~n67967 & n67979;
  assign n67981 = ~n67968 & n67980;
  assign n67982 = n67847 & ~n67981;
  assign n67983 = ~n67976 & ~n67982;
  assign n67984 = n67927 & n67983;
  assign n67985 = ~P2_P2_FLUSH_REG & ~P2_P2_MORE_REG;
  assign n67986 = n67984 & ~n67985;
  assign n67987 = ~n67882 & n67913;
  assign n67988 = ~n67847 & n67987;
  assign n67989 = n67973 & n67988;
  assign n67990 = ~n67966 & n67989;
  assign n67991 = n67882 & n67913;
  assign n67992 = ~n67847 & n67991;
  assign n67993 = n67973 & n67992;
  assign n67994 = ~n67966 & n67993;
  assign n67995 = n67915 & ~n67966;
  assign n67996 = ~n67882 & ~n67913;
  assign n67997 = n67851 & n67996;
  assign n67998 = ~n67966 & n67997;
  assign n67999 = ~n67990 & ~n67994;
  assign n68000 = ~n67995 & n67999;
  assign n68001 = ~n67998 & n68000;
  assign n68002 = ~n67691 & n67722;
  assign n68003 = ~n67754 & n68002;
  assign n68004 = n67849 & n68003;
  assign n68005 = n67996 & n68004;
  assign n68006 = ~P2_P2_INSTQUEUERD_ADDR_REG_0_ & P2_P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n68007 = ~n67933 & ~n68006;
  assign n68008 = n67958 & n68007;
  assign n68009 = ~n67962 & ~n68008;
  assign n68010 = n67963 & ~n68009;
  assign n68011 = n67944 & ~n68010;
  assign n68012 = n68005 & ~n68011;
  assign n68013 = n67991 & n68004;
  assign n68014 = ~n68011 & n68013;
  assign n68015 = n67849 & n67972;
  assign n68016 = n67914 & n68015;
  assign n68017 = n67948 & ~n68009;
  assign n68018 = n67952 & n68017;
  assign n68019 = n67944 & ~n68018;
  assign n68020 = n68016 & ~n68019;
  assign n68021 = n67996 & n68015;
  assign n68022 = ~n67958 & ~n68007;
  assign n68023 = n67963 & ~n68022;
  assign n68024 = n67962 & n68023;
  assign n68025 = n67944 & ~n68024;
  assign n68026 = n68021 & ~n68025;
  assign n68027 = ~n68012 & ~n68014;
  assign n68028 = ~n68020 & n68027;
  assign n68029 = ~n68026 & n68028;
  assign n68030 = n68001 & n68029;
  assign n68031 = ~n67984 & ~n68030;
  assign n68032 = ~n67882 & ~n68025;
  assign n68033 = n67882 & ~n68019;
  assign n68034 = ~n68032 & ~n68033;
  assign n68035 = ~n67913 & n68015;
  assign n68036 = n68034 & n68035;
  assign n68037 = n67816 & n67847;
  assign n68038 = n67691 & ~n67722;
  assign n68039 = n68037 & n68038;
  assign n68040 = n67991 & n68039;
  assign n68041 = ~n67785 & n68040;
  assign n68042 = n67851 & ~n67913;
  assign n68043 = ~n67989 & ~n68041;
  assign n68044 = ~n68042 & n68043;
  assign n68045 = n67722 & n67816;
  assign n68046 = ~n67754 & n67847;
  assign n68047 = ~n67785 & n67991;
  assign n68048 = n68046 & n68047;
  assign n68049 = n67691 & ~n67847;
  assign n68050 = n67754 & n67785;
  assign n68051 = n68049 & n68050;
  assign n68052 = ~n68048 & ~n68051;
  assign n68053 = n68045 & ~n68052;
  assign n68054 = n67996 & n68050;
  assign n68055 = n68039 & n68054;
  assign n68056 = n67816 & ~n67847;
  assign n68057 = n67785 & n67987;
  assign n68058 = n67972 & n68056;
  assign n68059 = n68057 & n68058;
  assign n68060 = ~n67882 & n68015;
  assign n68061 = ~n68059 & ~n68060;
  assign n68062 = ~n68053 & ~n68055;
  assign n68063 = n68061 & n68062;
  assign n68064 = n67722 & ~n67785;
  assign n68065 = ~n68038 & ~n68064;
  assign n68066 = n67816 & n68065;
  assign n68067 = ~n67847 & ~n68066;
  assign n68068 = ~n67785 & ~n68038;
  assign n68069 = ~n68002 & n68068;
  assign n68070 = ~n67816 & n68069;
  assign n68071 = n67914 & ~n68070;
  assign n68072 = n67971 & n67991;
  assign n68073 = n67691 & n67785;
  assign n68074 = ~n67848 & ~n68073;
  assign n68075 = ~n67882 & n68074;
  assign n68076 = n67722 & n67754;
  assign n68077 = n67913 & n68076;
  assign n68078 = ~n68072 & ~n68075;
  assign n68079 = ~n68077 & n68078;
  assign n68080 = ~n68071 & n68079;
  assign n68081 = n67847 & ~n68080;
  assign n68082 = ~n67816 & ~n68076;
  assign n68083 = n67691 & n68082;
  assign n68084 = n67785 & n67882;
  assign n68085 = n67913 & ~n68084;
  assign n68086 = n67816 & ~n68085;
  assign n68087 = ~n67691 & n68086;
  assign n68088 = ~n67785 & ~n67971;
  assign n68089 = ~n67914 & n68088;
  assign n68090 = ~n67754 & ~n68089;
  assign n68091 = n67722 & ~n67882;
  assign n68092 = n67785 & n68091;
  assign n68093 = n67754 & ~n67882;
  assign n68094 = n68002 & n68093;
  assign n68095 = ~n67971 & n67987;
  assign n68096 = ~n68092 & ~n68094;
  assign n68097 = ~n68095 & n68096;
  assign n68098 = ~n68083 & ~n68087;
  assign n68099 = ~n68090 & n68098;
  assign n68100 = n68097 & n68099;
  assign n68101 = ~n68067 & ~n68081;
  assign n68102 = n68100 & n68101;
  assign n68103 = n68063 & n68102;
  assign n68104 = ~n68040 & n68103;
  assign n68105 = P2_P2_INSTQUEUERD_ADDR_REG_0_ & ~n68104;
  assign n68106 = n68044 & ~n68105;
  assign n68107 = ~P2_P2_INSTQUEUERD_ADDR_REG_2_ & ~n68106;
  assign n68108 = P2_P2_INSTQUEUERD_ADDR_REG_1_ & n68107;
  assign n68109 = P2_P2_INSTQUEUERD_ADDR_REG_2_ & ~n68044;
  assign n68110 = ~P2_P2_INSTQUEUERD_ADDR_REG_1_ & n68109;
  assign n68111 = ~P2_P2_INSTQUEUERD_ADDR_REG_2_ & P2_P2_INSTQUEUERD_ADDR_REG_1_;
  assign n68112 = P2_P2_INSTQUEUERD_ADDR_REG_2_ & ~P2_P2_INSTQUEUERD_ADDR_REG_1_;
  assign n68113 = ~n68111 & ~n68112;
  assign n68114 = n67993 & ~n68113;
  assign n68115 = P2_P2_INSTQUEUERD_ADDR_REG_2_ & ~n67634;
  assign n68116 = ~n67635 & ~n68115;
  assign n68117 = ~n67991 & ~n67996;
  assign n68118 = n68116 & ~n68117;
  assign n68119 = n68004 & n68118;
  assign n68120 = ~n68114 & ~n68119;
  assign n68121 = n67882 & n68045;
  assign n68122 = ~n68046 & ~n68051;
  assign n68123 = n68121 & ~n68122;
  assign n68124 = n68050 & ~n68117;
  assign n68125 = n68039 & n68124;
  assign n68126 = ~n68123 & ~n68125;
  assign n68127 = n68061 & n68126;
  assign n68128 = n68102 & n68127;
  assign n68129 = n68115 & ~n68128;
  assign n68130 = n68120 & ~n68129;
  assign n68131 = ~n68108 & ~n68110;
  assign n68132 = n68130 & n68131;
  assign n68133 = n67754 & n67913;
  assign n68134 = ~n67816 & ~n67987;
  assign n68135 = n68068 & ~n68133;
  assign n68136 = n68134 & n68135;
  assign n68137 = ~n68094 & n68136;
  assign n68138 = n67847 & ~n68137;
  assign n68139 = ~n67847 & ~n67974;
  assign n68140 = n67914 & ~n68069;
  assign n68141 = ~n68138 & ~n68139;
  assign n68142 = ~n68140 & n68141;
  assign n68143 = n68011 & n68013;
  assign n68144 = n67966 & n67993;
  assign n68145 = n67966 & n67997;
  assign n68146 = ~n68144 & ~n68145;
  assign n68147 = ~n67541 & ~n68146;
  assign n68148 = ~n68143 & ~n68147;
  assign n68149 = n68005 & n68011;
  assign n68150 = ~n68002 & n68046;
  assign n68151 = ~n68149 & ~n68150;
  assign n68152 = n67966 & n67989;
  assign n68153 = n67915 & n67966;
  assign n68154 = ~n68152 & ~n68153;
  assign n68155 = n67918 & ~n68154;
  assign n68156 = n68151 & ~n68155;
  assign n68157 = n68142 & n68148;
  assign n68158 = n68156 & n68157;
  assign n68159 = ~n68132 & ~n68158;
  assign n68160 = P2_P2_INSTQUEUERD_ADDR_REG_2_ & n68158;
  assign n68161 = ~n68159 & ~n68160;
  assign n68162 = P2_P2_INSTQUEUERD_ADDR_REG_1_ & n67664;
  assign n68163 = ~n68106 & n68162;
  assign n68164 = P2_P2_INSTQUEUERD_ADDR_REG_2_ & n67634;
  assign n68165 = P2_P2_INSTQUEUERD_ADDR_REG_3_ & ~n68164;
  assign n68166 = ~n68127 & n68165;
  assign n68167 = P2_P2_INSTQUEUERD_ADDR_REG_2_ & P2_P2_INSTQUEUERD_ADDR_REG_1_;
  assign n68168 = ~P2_P2_INSTQUEUERD_ADDR_REG_3_ & n68167;
  assign n68169 = P2_P2_INSTQUEUERD_ADDR_REG_3_ & ~n68167;
  assign n68170 = ~n68168 & ~n68169;
  assign n68171 = n67993 & ~n68170;
  assign n68172 = ~n68166 & ~n68171;
  assign n68173 = ~n67754 & n68041;
  assign n68174 = n67754 & n68041;
  assign n68175 = ~n67915 & ~n67997;
  assign n68176 = ~n67989 & n68175;
  assign n68177 = ~n68173 & ~n68174;
  assign n68178 = n68176 & n68177;
  assign n68179 = n68102 & n68178;
  assign n68180 = n68169 & ~n68179;
  assign n68181 = P2_P2_INSTQUEUERD_ADDR_REG_3_ & ~P2_P2_INSTQUEUERD_ADDR_REG_0_;
  assign n68182 = ~n68102 & n68181;
  assign n68183 = ~n67634 & n67678;
  assign n68184 = ~P2_P2_INSTQUEUERD_ADDR_REG_2_ & ~n67634;
  assign n68185 = P2_P2_INSTQUEUERD_ADDR_REG_3_ & ~n68184;
  assign n68186 = ~n68183 & ~n68185;
  assign n68187 = ~n68117 & n68186;
  assign n68188 = n68004 & n68187;
  assign n68189 = ~n68182 & ~n68188;
  assign n68190 = n68172 & ~n68180;
  assign n68191 = n68189 & n68190;
  assign n68192 = ~n68163 & n68191;
  assign n68193 = ~n68158 & ~n68192;
  assign n68194 = P2_P2_INSTQUEUERD_ADDR_REG_3_ & n68158;
  assign n68195 = ~n68193 & ~n68194;
  assign n68196 = ~n68161 & ~n68195;
  assign n68197 = P2_P2_INSTQUEUERD_ADDR_REG_4_ & n68158;
  assign n68198 = P2_P2_INSTQUEUERD_ADDR_REG_3_ & n68167;
  assign n68199 = ~P2_P2_INSTQUEUERD_ADDR_REG_4_ & n68198;
  assign n68200 = P2_P2_INSTQUEUERD_ADDR_REG_4_ & ~n68198;
  assign n68201 = ~n68199 & ~n68200;
  assign n68202 = n67993 & ~n68201;
  assign n68203 = ~n68158 & n68202;
  assign n68204 = ~n68197 & ~n68203;
  assign n68205 = ~n68196 & n68204;
  assign n68206 = ~P2_P2_INSTQUEUEWR_ADDR_REG_3_ & ~n68195;
  assign n68207 = ~P2_P2_INSTQUEUEWR_ADDR_REG_4_ & ~n68204;
  assign n68208 = P2_P2_INSTQUEUEWR_ADDR_REG_2_ & n68161;
  assign n68209 = P2_P2_INSTQUEUEWR_ADDR_REG_3_ & n68195;
  assign n68210 = n68002 & n68048;
  assign n68211 = ~n68005 & ~n68210;
  assign n68212 = n68040 & n68050;
  assign n68213 = n68103 & ~n68212;
  assign n68214 = n68211 & n68213;
  assign n68215 = ~P2_P2_INSTQUEUERD_ADDR_REG_0_ & ~n68214;
  assign n68216 = P2_P2_INSTQUEUERD_ADDR_REG_0_ & ~n68044;
  assign n68217 = P2_P2_INSTQUEUERD_ADDR_REG_0_ & n67993;
  assign n68218 = ~n68215 & ~n68216;
  assign n68219 = ~n68217 & n68218;
  assign n68220 = ~n68158 & ~n68219;
  assign n68221 = P2_P2_INSTQUEUERD_ADDR_REG_0_ & n68158;
  assign n68222 = ~n68220 & ~n68221;
  assign n68223 = P2_P2_INSTQUEUEWR_ADDR_REG_0_ & n68222;
  assign n68224 = ~P2_P2_INSTQUEUEWR_ADDR_REG_1_ & ~n68223;
  assign n68225 = ~P2_P2_INSTQUEUEWR_ADDR_REG_2_ & ~n68161;
  assign n68226 = ~P2_P2_INSTQUEUERD_ADDR_REG_1_ & ~n68106;
  assign n68227 = ~P2_P2_INSTQUEUERD_ADDR_REG_1_ & n67993;
  assign n68228 = ~n67634 & ~n67647;
  assign n68229 = ~n68211 & n68228;
  assign n68230 = ~n68227 & ~n68229;
  assign n68231 = n67638 & ~n68213;
  assign n68232 = n68230 & ~n68231;
  assign n68233 = ~n68226 & n68232;
  assign n68234 = ~n68158 & ~n68233;
  assign n68235 = P2_P2_INSTQUEUERD_ADDR_REG_1_ & n68158;
  assign n68236 = ~n68234 & ~n68235;
  assign n68237 = P2_P2_INSTQUEUEWR_ADDR_REG_1_ & n68223;
  assign n68238 = ~n68236 & ~n68237;
  assign n68239 = ~n68224 & ~n68225;
  assign n68240 = ~n68238 & n68239;
  assign n68241 = ~n68208 & ~n68209;
  assign n68242 = ~n68240 & n68241;
  assign n68243 = ~n68206 & ~n68207;
  assign n68244 = ~n68242 & n68243;
  assign n68245 = P2_P2_INSTQUEUEWR_ADDR_REG_4_ & n68204;
  assign n68246 = ~n68244 & ~n68245;
  assign n68247 = ~n67986 & ~n68031;
  assign n68248 = ~n68036 & n68247;
  assign n68249 = n68205 & n68248;
  assign n68250 = ~n68246 & n68249;
  assign n68251 = n67917 & n68250;
  assign n68252 = P2_P2_STATE2_REG_0_ & ~n68251;
  assign n68253 = ~n67628 & ~n68252;
  assign n68254 = P2_P2_STATE2_REG_2_ & n68253;
  assign n68255 = P2_P2_STATE2_REG_0_ & ~n68254;
  assign n68256 = n67626 & n68255;
  assign n68257 = P2_P2_STATE2_REG_3_ & ~n68255;
  assign n12576 = n68256 | n68257;
  assign n68259 = ~P2_P2_STATE2_REG_2_ & ~n67541;
  assign n68260 = P2_P2_STATE2_REG_0_ & ~n68259;
  assign n68261 = ~P2_P2_STATE2_REG_0_ & ~P2_P2_STATEBS16_REG;
  assign n68262 = ~n68260 & ~n68261;
  assign n68263 = P2_P2_STATE2_REG_1_ & n68262;
  assign n68264 = P2_P2_STATE2_REG_2_ & ~P2_P2_STATE2_REG_1_;
  assign n68265 = ~n68263 & ~n68264;
  assign n68266 = P2_P2_STATE2_REG_2_ & ~n68255;
  assign n12581 = ~n68265 | n68266;
  assign n68268 = P2_P2_STATE2_REG_0_ & n68264;
  assign n68269 = ~n68254 & n68268;
  assign n68270 = ~P2_P2_STATE2_REG_2_ & P2_P2_STATE2_REG_0_;
  assign n68271 = n67541 & n68270;
  assign n68272 = ~n68254 & ~n68271;
  assign n68273 = P2_P2_STATE2_REG_1_ & ~n68272;
  assign n68274 = ~P2_P2_STATE2_REG_3_ & ~P2_P2_STATE2_REG_1_;
  assign n68275 = ~n67541 & n68274;
  assign n68276 = n68255 & n68275;
  assign n68277 = P2_P2_STATE2_REG_1_ & ~P2_P2_STATE2_REG_0_;
  assign n68278 = ~P2_P2_STATE2_REG_2_ & n68277;
  assign n68279 = ~P2_P2_STATEBS16_REG & n68278;
  assign n68280 = ~n68269 & ~n68273;
  assign n68281 = ~n68276 & n68280;
  assign n12586 = n68279 | ~n68281;
  assign n68283 = P2_P2_STATE2_REG_3_ & ~P2_P2_INSTQUEUERD_ADDR_REG_4_;
  assign n68284 = ~P2_P2_STATE2_REG_2_ & ~P2_P2_STATE2_REG_1_;
  assign n68285 = n68283 & n68284;
  assign n68286 = ~n68254 & ~n68285;
  assign n68287 = ~P2_P2_STATE2_REG_0_ & n68286;
  assign n68288 = P2_P2_INSTADDRPOINTER_REG_0_ & P2_P2_INSTADDRPOINTER_REG_31_;
  assign n68289 = P2_P2_INSTADDRPOINTER_REG_0_ & ~P2_P2_INSTADDRPOINTER_REG_31_;
  assign n68290 = ~n68288 & ~n68289;
  assign n68291 = P2_P2_FLUSH_REG & n68290;
  assign n68292 = P2_P2_INSTQUEUERD_ADDR_REG_0_ & ~P2_P2_FLUSH_REG;
  assign n68293 = ~n68291 & ~n68292;
  assign n68294 = P2_P2_INSTADDRPOINTER_REG_0_ & ~P2_P2_INSTADDRPOINTER_REG_1_;
  assign n68295 = ~P2_P2_INSTADDRPOINTER_REG_0_ & P2_P2_INSTADDRPOINTER_REG_1_;
  assign n68296 = ~n68294 & ~n68295;
  assign n68297 = P2_P2_INSTADDRPOINTER_REG_31_ & ~n68296;
  assign n68298 = P2_P2_INSTADDRPOINTER_REG_1_ & ~P2_P2_INSTADDRPOINTER_REG_31_;
  assign n68299 = ~n68297 & ~n68298;
  assign n68300 = ~n68290 & n68299;
  assign n68301 = P2_P2_FLUSH_REG & n68300;
  assign n68302 = P2_P2_INSTQUEUERD_ADDR_REG_1_ & ~P2_P2_FLUSH_REG;
  assign n68303 = ~n68301 & ~n68302;
  assign n68304 = n68293 & n68303;
  assign n68305 = P2_P2_INSTQUEUERD_ADDR_REG_3_ & ~P2_P2_FLUSH_REG;
  assign n68306 = ~n68290 & ~n68299;
  assign n68307 = P2_P2_FLUSH_REG & n68306;
  assign n68308 = P2_P2_INSTQUEUERD_ADDR_REG_2_ & ~P2_P2_FLUSH_REG;
  assign n68309 = ~n68307 & ~n68308;
  assign n68310 = ~n68304 & n68305;
  assign n68311 = ~n68309 & n68310;
  assign n68312 = P2_P2_INSTQUEUERD_ADDR_REG_4_ & ~P2_P2_FLUSH_REG;
  assign n68313 = ~n68311 & ~n68312;
  assign n68314 = n67626 & n68313;
  assign n68315 = ~n68254 & ~n68314;
  assign n68316 = P2_P2_STATE2_REG_0_ & ~n68315;
  assign n68317 = P2_P2_STATE2_REG_3_ & P2_P2_STATE2_REG_0_;
  assign n68318 = n68284 & n68317;
  assign n68319 = ~n68271 & ~n68318;
  assign n68320 = ~n68250 & n68268;
  assign n68321 = n68319 & ~n68320;
  assign n68322 = ~n68287 & ~n68316;
  assign n12591 = ~n68321 | ~n68322;
  assign n68324 = P2_P2_INSTQUEUEWR_ADDR_REG_1_ & P2_P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n68325 = P2_P2_INSTQUEUEWR_ADDR_REG_2_ & n68324;
  assign n68326 = P2_P2_INSTQUEUEWR_ADDR_REG_3_ & n68325;
  assign n68327 = P2_P2_STATE2_REG_3_ & ~n68326;
  assign n68328 = ~P2_P2_STATE2_REG_2_ & P2_P2_STATE2_REG_1_;
  assign n68329 = ~n68264 & ~n68328;
  assign n68330 = ~n68283 & n68329;
  assign n68331 = ~P2_P2_STATE2_REG_0_ & ~n68330;
  assign n68332 = ~n68327 & n68331;
  assign n68333 = ~P2_P2_INSTQUEUEWR_ADDR_REG_2_ & n68324;
  assign n68334 = P2_P2_INSTQUEUEWR_ADDR_REG_2_ & ~n68324;
  assign n68335 = ~n68333 & ~n68334;
  assign n68336 = ~P2_P2_INSTQUEUEWR_ADDR_REG_3_ & n68325;
  assign n68337 = P2_P2_INSTQUEUEWR_ADDR_REG_3_ & ~n68325;
  assign n68338 = ~n68336 & ~n68337;
  assign n68339 = ~n68335 & ~n68338;
  assign n68340 = ~P2_P2_INSTQUEUEWR_ADDR_REG_1_ & P2_P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n68341 = P2_P2_INSTQUEUEWR_ADDR_REG_1_ & ~P2_P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n68342 = ~n68340 & ~n68341;
  assign n68343 = ~P2_P2_INSTQUEUEWR_ADDR_REG_0_ & ~n68342;
  assign n68344 = n68339 & n68343;
  assign n68345 = ~n68326 & ~n68344;
  assign n68346 = ~P2_P2_STATE2_REG_3_ & ~P2_P2_STATE2_REG_2_;
  assign n68347 = ~P2_P2_STATEBS16_REG & n68346;
  assign n68348 = ~P2_P2_STATE2_REG_2_ & ~n68347;
  assign n68349 = P2_P2_INSTQUEUEWR_ADDR_REG_0_ & ~n68342;
  assign n68350 = ~P2_P2_INSTQUEUEWR_ADDR_REG_0_ & n68342;
  assign n68351 = ~n68349 & ~n68350;
  assign n68352 = ~P2_P2_INSTQUEUEWR_ADDR_REG_0_ & ~n68351;
  assign n68353 = P2_P2_INSTQUEUEWR_ADDR_REG_0_ & n68351;
  assign n68354 = ~n68352 & ~n68353;
  assign n68355 = ~P2_P2_INSTQUEUEWR_ADDR_REG_0_ & ~n68354;
  assign n68356 = ~n68335 & ~n68343;
  assign n68357 = n68335 & n68343;
  assign n68358 = ~n68356 & ~n68357;
  assign n68359 = P2_P2_INSTQUEUEWR_ADDR_REG_0_ & ~n68351;
  assign n68360 = ~n68358 & ~n68359;
  assign n68361 = n68358 & n68359;
  assign n68362 = ~n68360 & ~n68361;
  assign n68363 = ~n68335 & n68338;
  assign n68364 = n68343 & n68363;
  assign n68365 = ~n68335 & n68343;
  assign n68366 = ~n68338 & ~n68365;
  assign n68367 = ~n68364 & ~n68366;
  assign n68368 = n68358 & ~n68367;
  assign n68369 = ~n68359 & ~n68367;
  assign n68370 = ~n68368 & ~n68369;
  assign n68371 = ~n68358 & n68367;
  assign n68372 = n68359 & n68371;
  assign n68373 = n68370 & ~n68372;
  assign n68374 = ~n68362 & ~n68373;
  assign n68375 = n68355 & n68374;
  assign n68376 = ~n68358 & ~n68367;
  assign n68377 = n68359 & n68376;
  assign n68378 = ~n68375 & ~n68377;
  assign n68379 = n68348 & ~n68378;
  assign n68380 = n68345 & ~n68379;
  assign n68381 = n68332 & ~n68380;
  assign n68382 = P2_P2_INSTQUEUE_REG_15__7_ & ~n68381;
  assign n68383 = P2_BUF1_REG_23_ & n12836_1;
  assign n68384 = P2_BUF2_REG_23_ & ~n12836_1;
  assign n68385 = ~n68383 & ~n68384;
  assign n68386 = P2_P2_STATEBS16_REG & n68346;
  assign n68387 = n68331 & n68386;
  assign n68388 = ~n68385 & n68387;
  assign n68389 = n68377 & n68388;
  assign n68390 = P2_P2_STATE2_REG_3_ & n68331;
  assign n68391 = ~n67785 & n68390;
  assign n68392 = n68326 & n68391;
  assign n68393 = ~n68389 & ~n68392;
  assign n68394 = P2_BUF1_REG_31_ & n12836_1;
  assign n68395 = P2_BUF2_REG_31_ & ~n12836_1;
  assign n68396 = ~n68394 & ~n68395;
  assign n68397 = n68387 & ~n68396;
  assign n68398 = n68375 & n68397;
  assign n68399 = n68393 & ~n68398;
  assign n68400 = n68378 & n68386;
  assign n68401 = n68348 & ~n68400;
  assign n68402 = ~n68345 & ~n68401;
  assign n68403 = P2_BUF1_REG_7_ & n12836_1;
  assign n68404 = P2_BUF2_REG_7_ & ~n12836_1;
  assign n68405 = ~n68403 & ~n68404;
  assign n68406 = n68331 & ~n68405;
  assign n68407 = n68402 & n68406;
  assign n68408 = ~n68382 & n68399;
  assign n12596 = n68407 | ~n68408;
  assign n68410 = P2_P2_INSTQUEUE_REG_15__6_ & ~n68381;
  assign n68411 = P2_BUF1_REG_22_ & n12836_1;
  assign n68412 = P2_BUF2_REG_22_ & ~n12836_1;
  assign n68413 = ~n68411 & ~n68412;
  assign n68414 = n68387 & ~n68413;
  assign n68415 = n68377 & n68414;
  assign n68416 = ~n67722 & n68390;
  assign n68417 = n68326 & n68416;
  assign n68418 = ~n68415 & ~n68417;
  assign n68419 = P2_BUF1_REG_30_ & n12836_1;
  assign n68420 = P2_BUF2_REG_30_ & ~n12836_1;
  assign n68421 = ~n68419 & ~n68420;
  assign n68422 = n68387 & ~n68421;
  assign n68423 = n68375 & n68422;
  assign n68424 = n68418 & ~n68423;
  assign n68425 = P2_BUF1_REG_6_ & n12836_1;
  assign n68426 = P2_BUF2_REG_6_ & ~n12836_1;
  assign n68427 = ~n68425 & ~n68426;
  assign n68428 = n68331 & ~n68427;
  assign n68429 = n68402 & n68428;
  assign n68430 = ~n68410 & n68424;
  assign n12601 = n68429 | ~n68430;
  assign n68432 = P2_P2_INSTQUEUE_REG_15__5_ & ~n68381;
  assign n68433 = P2_BUF1_REG_21_ & n12836_1;
  assign n68434 = P2_BUF2_REG_21_ & ~n12836_1;
  assign n68435 = ~n68433 & ~n68434;
  assign n68436 = n68387 & ~n68435;
  assign n68437 = n68377 & n68436;
  assign n68438 = ~n67691 & n68390;
  assign n68439 = n68326 & n68438;
  assign n68440 = ~n68437 & ~n68439;
  assign n68441 = P2_BUF1_REG_29_ & n12836_1;
  assign n68442 = P2_BUF2_REG_29_ & ~n12836_1;
  assign n68443 = ~n68441 & ~n68442;
  assign n68444 = n68387 & ~n68443;
  assign n68445 = n68375 & n68444;
  assign n68446 = n68440 & ~n68445;
  assign n68447 = P2_BUF1_REG_5_ & n12836_1;
  assign n68448 = P2_BUF2_REG_5_ & ~n12836_1;
  assign n68449 = ~n68447 & ~n68448;
  assign n68450 = n68331 & ~n68449;
  assign n68451 = n68402 & n68450;
  assign n68452 = ~n68432 & n68446;
  assign n12606 = n68451 | ~n68452;
  assign n68454 = P2_P2_INSTQUEUE_REG_15__4_ & ~n68381;
  assign n68455 = P2_BUF1_REG_20_ & n12836_1;
  assign n68456 = P2_BUF2_REG_20_ & ~n12836_1;
  assign n68457 = ~n68455 & ~n68456;
  assign n68458 = n68387 & ~n68457;
  assign n68459 = n68377 & n68458;
  assign n68460 = ~n67754 & n68390;
  assign n68461 = n68326 & n68460;
  assign n68462 = ~n68459 & ~n68461;
  assign n68463 = P2_BUF1_REG_28_ & n12836_1;
  assign n68464 = P2_BUF2_REG_28_ & ~n12836_1;
  assign n68465 = ~n68463 & ~n68464;
  assign n68466 = n68387 & ~n68465;
  assign n68467 = n68375 & n68466;
  assign n68468 = n68462 & ~n68467;
  assign n68469 = P2_BUF1_REG_4_ & n12836_1;
  assign n68470 = P2_BUF2_REG_4_ & ~n12836_1;
  assign n68471 = ~n68469 & ~n68470;
  assign n68472 = n68331 & ~n68471;
  assign n68473 = n68402 & n68472;
  assign n68474 = ~n68454 & n68468;
  assign n12611 = n68473 | ~n68474;
  assign n68476 = P2_P2_INSTQUEUE_REG_15__3_ & ~n68381;
  assign n68477 = P2_BUF1_REG_19_ & n12836_1;
  assign n68478 = P2_BUF2_REG_19_ & ~n12836_1;
  assign n68479 = ~n68477 & ~n68478;
  assign n68480 = n68387 & ~n68479;
  assign n68481 = n68377 & n68480;
  assign n68482 = ~n67816 & n68390;
  assign n68483 = n68326 & n68482;
  assign n68484 = ~n68481 & ~n68483;
  assign n68485 = P2_BUF1_REG_27_ & n12836_1;
  assign n68486 = P2_BUF2_REG_27_ & ~n12836_1;
  assign n68487 = ~n68485 & ~n68486;
  assign n68488 = n68387 & ~n68487;
  assign n68489 = n68375 & n68488;
  assign n68490 = n68484 & ~n68489;
  assign n68491 = P2_BUF1_REG_3_ & n12836_1;
  assign n68492 = P2_BUF2_REG_3_ & ~n12836_1;
  assign n68493 = ~n68491 & ~n68492;
  assign n68494 = n68331 & ~n68493;
  assign n68495 = n68402 & n68494;
  assign n68496 = ~n68476 & n68490;
  assign n12616 = n68495 | ~n68496;
  assign n68498 = P2_P2_INSTQUEUE_REG_15__2_ & ~n68381;
  assign n68499 = P2_BUF1_REG_18_ & n12836_1;
  assign n68500 = P2_BUF2_REG_18_ & ~n12836_1;
  assign n68501 = ~n68499 & ~n68500;
  assign n68502 = n68387 & ~n68501;
  assign n68503 = n68377 & n68502;
  assign n68504 = ~n67847 & n68390;
  assign n68505 = n68326 & n68504;
  assign n68506 = ~n68503 & ~n68505;
  assign n68507 = P2_BUF1_REG_26_ & n12836_1;
  assign n68508 = P2_BUF2_REG_26_ & ~n12836_1;
  assign n68509 = ~n68507 & ~n68508;
  assign n68510 = n68387 & ~n68509;
  assign n68511 = n68375 & n68510;
  assign n68512 = n68506 & ~n68511;
  assign n68513 = P2_BUF1_REG_2_ & n12836_1;
  assign n68514 = P2_BUF2_REG_2_ & ~n12836_1;
  assign n68515 = ~n68513 & ~n68514;
  assign n68516 = n68331 & ~n68515;
  assign n68517 = n68402 & n68516;
  assign n68518 = ~n68498 & n68512;
  assign n12621 = n68517 | ~n68518;
  assign n68520 = P2_P2_INSTQUEUE_REG_15__1_ & ~n68381;
  assign n68521 = P2_BUF1_REG_17_ & n12836_1;
  assign n68522 = P2_BUF2_REG_17_ & ~n12836_1;
  assign n68523 = ~n68521 & ~n68522;
  assign n68524 = n68387 & ~n68523;
  assign n68525 = n68377 & n68524;
  assign n68526 = ~n67882 & n68390;
  assign n68527 = n68326 & n68526;
  assign n68528 = ~n68525 & ~n68527;
  assign n68529 = P2_BUF1_REG_25_ & n12836_1;
  assign n68530 = P2_BUF2_REG_25_ & ~n12836_1;
  assign n68531 = ~n68529 & ~n68530;
  assign n68532 = n68387 & ~n68531;
  assign n68533 = n68375 & n68532;
  assign n68534 = n68528 & ~n68533;
  assign n68535 = P2_BUF1_REG_1_ & n12836_1;
  assign n68536 = P2_BUF2_REG_1_ & ~n12836_1;
  assign n68537 = ~n68535 & ~n68536;
  assign n68538 = n68331 & ~n68537;
  assign n68539 = n68402 & n68538;
  assign n68540 = ~n68520 & n68534;
  assign n12626 = n68539 | ~n68540;
  assign n68542 = P2_P2_INSTQUEUE_REG_15__0_ & ~n68381;
  assign n68543 = P2_BUF1_REG_16_ & n12836_1;
  assign n68544 = P2_BUF2_REG_16_ & ~n12836_1;
  assign n68545 = ~n68543 & ~n68544;
  assign n68546 = n68387 & ~n68545;
  assign n68547 = n68377 & n68546;
  assign n68548 = ~n67913 & n68390;
  assign n68549 = n68326 & n68548;
  assign n68550 = ~n68547 & ~n68549;
  assign n68551 = P2_BUF1_REG_24_ & n12836_1;
  assign n68552 = P2_BUF2_REG_24_ & ~n12836_1;
  assign n68553 = ~n68551 & ~n68552;
  assign n68554 = n68387 & ~n68553;
  assign n68555 = n68375 & n68554;
  assign n68556 = n68550 & ~n68555;
  assign n68557 = P2_BUF1_REG_0_ & n12836_1;
  assign n68558 = P2_BUF2_REG_0_ & ~n12836_1;
  assign n68559 = ~n68557 & ~n68558;
  assign n68560 = n68331 & ~n68559;
  assign n68561 = n68402 & n68560;
  assign n68562 = ~n68542 & n68556;
  assign n12631 = n68561 | ~n68562;
  assign n68564 = P2_P2_INSTQUEUEWR_ADDR_REG_3_ & P2_P2_INSTQUEUEWR_ADDR_REG_1_;
  assign n68565 = P2_P2_INSTQUEUEWR_ADDR_REG_2_ & ~P2_P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n68566 = n68564 & n68565;
  assign n68567 = P2_P2_STATE2_REG_3_ & ~n68566;
  assign n68568 = n68331 & ~n68567;
  assign n68569 = n68339 & n68349;
  assign n68570 = ~n68566 & ~n68569;
  assign n68571 = P2_P2_INSTQUEUEWR_ADDR_REG_0_ & ~n68354;
  assign n68572 = n68374 & n68571;
  assign n68573 = n68352 & n68376;
  assign n68574 = ~n68572 & ~n68573;
  assign n68575 = n68348 & ~n68574;
  assign n68576 = n68570 & ~n68575;
  assign n68577 = n68568 & ~n68576;
  assign n68578 = P2_P2_INSTQUEUE_REG_14__7_ & ~n68577;
  assign n68579 = n68388 & n68573;
  assign n68580 = n68391 & n68566;
  assign n68581 = ~n68579 & ~n68580;
  assign n68582 = n68397 & n68572;
  assign n68583 = n68581 & ~n68582;
  assign n68584 = n68386 & n68574;
  assign n68585 = n68348 & ~n68584;
  assign n68586 = ~n68570 & ~n68585;
  assign n68587 = n68406 & n68586;
  assign n68588 = ~n68578 & n68583;
  assign n12636 = n68587 | ~n68588;
  assign n68590 = P2_P2_INSTQUEUE_REG_14__6_ & ~n68577;
  assign n68591 = n68414 & n68573;
  assign n68592 = n68416 & n68566;
  assign n68593 = ~n68591 & ~n68592;
  assign n68594 = n68422 & n68572;
  assign n68595 = n68593 & ~n68594;
  assign n68596 = n68428 & n68586;
  assign n68597 = ~n68590 & n68595;
  assign n12641 = n68596 | ~n68597;
  assign n68599 = P2_P2_INSTQUEUE_REG_14__5_ & ~n68577;
  assign n68600 = n68436 & n68573;
  assign n68601 = n68438 & n68566;
  assign n68602 = ~n68600 & ~n68601;
  assign n68603 = n68444 & n68572;
  assign n68604 = n68602 & ~n68603;
  assign n68605 = n68450 & n68586;
  assign n68606 = ~n68599 & n68604;
  assign n12646 = n68605 | ~n68606;
  assign n68608 = P2_P2_INSTQUEUE_REG_14__4_ & ~n68577;
  assign n68609 = n68458 & n68573;
  assign n68610 = n68460 & n68566;
  assign n68611 = ~n68609 & ~n68610;
  assign n68612 = n68466 & n68572;
  assign n68613 = n68611 & ~n68612;
  assign n68614 = n68472 & n68586;
  assign n68615 = ~n68608 & n68613;
  assign n12651 = n68614 | ~n68615;
  assign n68617 = P2_P2_INSTQUEUE_REG_14__3_ & ~n68577;
  assign n68618 = n68480 & n68573;
  assign n68619 = n68482 & n68566;
  assign n68620 = ~n68618 & ~n68619;
  assign n68621 = n68488 & n68572;
  assign n68622 = n68620 & ~n68621;
  assign n68623 = n68494 & n68586;
  assign n68624 = ~n68617 & n68622;
  assign n12656 = n68623 | ~n68624;
  assign n68626 = P2_P2_INSTQUEUE_REG_14__2_ & ~n68577;
  assign n68627 = n68502 & n68573;
  assign n68628 = n68504 & n68566;
  assign n68629 = ~n68627 & ~n68628;
  assign n68630 = n68510 & n68572;
  assign n68631 = n68629 & ~n68630;
  assign n68632 = n68516 & n68586;
  assign n68633 = ~n68626 & n68631;
  assign n12661 = n68632 | ~n68633;
  assign n68635 = P2_P2_INSTQUEUE_REG_14__1_ & ~n68577;
  assign n68636 = n68524 & n68573;
  assign n68637 = n68526 & n68566;
  assign n68638 = ~n68636 & ~n68637;
  assign n68639 = n68532 & n68572;
  assign n68640 = n68638 & ~n68639;
  assign n68641 = n68538 & n68586;
  assign n68642 = ~n68635 & n68640;
  assign n12666 = n68641 | ~n68642;
  assign n68644 = P2_P2_INSTQUEUE_REG_14__0_ & ~n68577;
  assign n68645 = n68546 & n68573;
  assign n68646 = n68548 & n68566;
  assign n68647 = ~n68645 & ~n68646;
  assign n68648 = n68554 & n68572;
  assign n68649 = n68647 & ~n68648;
  assign n68650 = n68560 & n68586;
  assign n68651 = ~n68644 & n68649;
  assign n12671 = n68650 | ~n68651;
  assign n68653 = P2_P2_INSTQUEUEWR_ADDR_REG_3_ & P2_P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n68654 = n68340 & n68653;
  assign n68655 = P2_P2_STATE2_REG_3_ & ~n68654;
  assign n68656 = n68331 & ~n68655;
  assign n68657 = n68339 & n68350;
  assign n68658 = ~n68654 & ~n68657;
  assign n68659 = ~P2_P2_INSTQUEUEWR_ADDR_REG_0_ & n68354;
  assign n68660 = n68374 & n68659;
  assign n68661 = n68353 & n68376;
  assign n68662 = ~n68660 & ~n68661;
  assign n68663 = n68348 & ~n68662;
  assign n68664 = n68658 & ~n68663;
  assign n68665 = n68656 & ~n68664;
  assign n68666 = P2_P2_INSTQUEUE_REG_13__7_ & ~n68665;
  assign n68667 = n68388 & n68661;
  assign n68668 = n68391 & n68654;
  assign n68669 = ~n68667 & ~n68668;
  assign n68670 = n68397 & n68660;
  assign n68671 = n68669 & ~n68670;
  assign n68672 = n68386 & n68662;
  assign n68673 = n68348 & ~n68672;
  assign n68674 = ~n68658 & ~n68673;
  assign n68675 = n68406 & n68674;
  assign n68676 = ~n68666 & n68671;
  assign n12676 = n68675 | ~n68676;
  assign n68678 = P2_P2_INSTQUEUE_REG_13__6_ & ~n68665;
  assign n68679 = n68414 & n68661;
  assign n68680 = n68416 & n68654;
  assign n68681 = ~n68679 & ~n68680;
  assign n68682 = n68422 & n68660;
  assign n68683 = n68681 & ~n68682;
  assign n68684 = n68428 & n68674;
  assign n68685 = ~n68678 & n68683;
  assign n12681 = n68684 | ~n68685;
  assign n68687 = P2_P2_INSTQUEUE_REG_13__5_ & ~n68665;
  assign n68688 = n68436 & n68661;
  assign n68689 = n68438 & n68654;
  assign n68690 = ~n68688 & ~n68689;
  assign n68691 = n68444 & n68660;
  assign n68692 = n68690 & ~n68691;
  assign n68693 = n68450 & n68674;
  assign n68694 = ~n68687 & n68692;
  assign n12686 = n68693 | ~n68694;
  assign n68696 = P2_P2_INSTQUEUE_REG_13__4_ & ~n68665;
  assign n68697 = n68458 & n68661;
  assign n68698 = n68460 & n68654;
  assign n68699 = ~n68697 & ~n68698;
  assign n68700 = n68466 & n68660;
  assign n68701 = n68699 & ~n68700;
  assign n68702 = n68472 & n68674;
  assign n68703 = ~n68696 & n68701;
  assign n12691 = n68702 | ~n68703;
  assign n68705 = P2_P2_INSTQUEUE_REG_13__3_ & ~n68665;
  assign n68706 = n68480 & n68661;
  assign n68707 = n68482 & n68654;
  assign n68708 = ~n68706 & ~n68707;
  assign n68709 = n68488 & n68660;
  assign n68710 = n68708 & ~n68709;
  assign n68711 = n68494 & n68674;
  assign n68712 = ~n68705 & n68710;
  assign n12696 = n68711 | ~n68712;
  assign n68714 = P2_P2_INSTQUEUE_REG_13__2_ & ~n68665;
  assign n68715 = n68502 & n68661;
  assign n68716 = n68504 & n68654;
  assign n68717 = ~n68715 & ~n68716;
  assign n68718 = n68510 & n68660;
  assign n68719 = n68717 & ~n68718;
  assign n68720 = n68516 & n68674;
  assign n68721 = ~n68714 & n68719;
  assign n12701 = n68720 | ~n68721;
  assign n68723 = P2_P2_INSTQUEUE_REG_13__1_ & ~n68665;
  assign n68724 = n68524 & n68661;
  assign n68725 = n68526 & n68654;
  assign n68726 = ~n68724 & ~n68725;
  assign n68727 = n68532 & n68660;
  assign n68728 = n68726 & ~n68727;
  assign n68729 = n68538 & n68674;
  assign n68730 = ~n68723 & n68728;
  assign n12706 = n68729 | ~n68730;
  assign n68732 = P2_P2_INSTQUEUE_REG_13__0_ & ~n68665;
  assign n68733 = n68546 & n68661;
  assign n68734 = n68548 & n68654;
  assign n68735 = ~n68733 & ~n68734;
  assign n68736 = n68554 & n68660;
  assign n68737 = n68735 & ~n68736;
  assign n68738 = n68560 & n68674;
  assign n68739 = ~n68732 & n68737;
  assign n12711 = n68738 | ~n68739;
  assign n68741 = P2_P2_INSTQUEUEWR_ADDR_REG_3_ & ~P2_P2_INSTQUEUEWR_ADDR_REG_1_;
  assign n68742 = n68565 & n68741;
  assign n68743 = P2_P2_STATE2_REG_3_ & ~n68742;
  assign n68744 = n68331 & ~n68743;
  assign n68745 = P2_P2_INSTQUEUEWR_ADDR_REG_0_ & n68354;
  assign n68746 = n68374 & n68745;
  assign n68747 = ~P2_P2_INSTQUEUEWR_ADDR_REG_0_ & n68351;
  assign n68748 = n68376 & n68747;
  assign n68749 = ~n68746 & ~n68748;
  assign n68750 = n68348 & ~n68749;
  assign n68751 = n68339 & n68342;
  assign n68752 = ~n68750 & ~n68751;
  assign n68753 = n68744 & ~n68752;
  assign n68754 = P2_P2_INSTQUEUE_REG_12__7_ & ~n68753;
  assign n68755 = n68388 & n68748;
  assign n68756 = n68391 & n68742;
  assign n68757 = ~n68755 & ~n68756;
  assign n68758 = n68397 & n68746;
  assign n68759 = n68757 & ~n68758;
  assign n68760 = n68386 & n68749;
  assign n68761 = n68348 & ~n68760;
  assign n68762 = n68751 & ~n68761;
  assign n68763 = n68406 & n68762;
  assign n68764 = ~n68754 & n68759;
  assign n12716 = n68763 | ~n68764;
  assign n68766 = P2_P2_INSTQUEUE_REG_12__6_ & ~n68753;
  assign n68767 = n68414 & n68748;
  assign n68768 = n68416 & n68742;
  assign n68769 = ~n68767 & ~n68768;
  assign n68770 = n68422 & n68746;
  assign n68771 = n68769 & ~n68770;
  assign n68772 = n68428 & n68762;
  assign n68773 = ~n68766 & n68771;
  assign n12721 = n68772 | ~n68773;
  assign n68775 = P2_P2_INSTQUEUE_REG_12__5_ & ~n68753;
  assign n68776 = n68436 & n68748;
  assign n68777 = n68438 & n68742;
  assign n68778 = ~n68776 & ~n68777;
  assign n68779 = n68444 & n68746;
  assign n68780 = n68778 & ~n68779;
  assign n68781 = n68450 & n68762;
  assign n68782 = ~n68775 & n68780;
  assign n12726 = n68781 | ~n68782;
  assign n68784 = P2_P2_INSTQUEUE_REG_12__4_ & ~n68753;
  assign n68785 = n68458 & n68748;
  assign n68786 = n68460 & n68742;
  assign n68787 = ~n68785 & ~n68786;
  assign n68788 = n68466 & n68746;
  assign n68789 = n68787 & ~n68788;
  assign n68790 = n68472 & n68762;
  assign n68791 = ~n68784 & n68789;
  assign n12731 = n68790 | ~n68791;
  assign n68793 = P2_P2_INSTQUEUE_REG_12__3_ & ~n68753;
  assign n68794 = n68480 & n68748;
  assign n68795 = n68482 & n68742;
  assign n68796 = ~n68794 & ~n68795;
  assign n68797 = n68488 & n68746;
  assign n68798 = n68796 & ~n68797;
  assign n68799 = n68494 & n68762;
  assign n68800 = ~n68793 & n68798;
  assign n12736 = n68799 | ~n68800;
  assign n68802 = P2_P2_INSTQUEUE_REG_12__2_ & ~n68753;
  assign n68803 = n68502 & n68748;
  assign n68804 = n68504 & n68742;
  assign n68805 = ~n68803 & ~n68804;
  assign n68806 = n68510 & n68746;
  assign n68807 = n68805 & ~n68806;
  assign n68808 = n68516 & n68762;
  assign n68809 = ~n68802 & n68807;
  assign n12741 = n68808 | ~n68809;
  assign n68811 = P2_P2_INSTQUEUE_REG_12__1_ & ~n68753;
  assign n68812 = n68524 & n68748;
  assign n68813 = n68526 & n68742;
  assign n68814 = ~n68812 & ~n68813;
  assign n68815 = n68532 & n68746;
  assign n68816 = n68814 & ~n68815;
  assign n68817 = n68538 & n68762;
  assign n68818 = ~n68811 & n68816;
  assign n12746 = n68817 | ~n68818;
  assign n68820 = P2_P2_INSTQUEUE_REG_12__0_ & ~n68753;
  assign n68821 = n68546 & n68748;
  assign n68822 = n68548 & n68742;
  assign n68823 = ~n68821 & ~n68822;
  assign n68824 = n68554 & n68746;
  assign n68825 = n68823 & ~n68824;
  assign n68826 = n68560 & n68762;
  assign n68827 = ~n68820 & n68825;
  assign n12751 = n68826 | ~n68827;
  assign n68829 = P2_P2_INSTQUEUEWR_ADDR_REG_3_ & ~P2_P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n68830 = n68324 & n68829;
  assign n68831 = P2_P2_STATE2_REG_3_ & ~n68830;
  assign n68832 = n68331 & ~n68831;
  assign n68833 = n68335 & ~n68338;
  assign n68834 = n68343 & n68833;
  assign n68835 = ~n68830 & ~n68834;
  assign n68836 = n68362 & ~n68373;
  assign n68837 = n68355 & n68836;
  assign n68838 = n68359 & n68368;
  assign n68839 = ~n68837 & ~n68838;
  assign n68840 = n68348 & ~n68839;
  assign n68841 = n68835 & ~n68840;
  assign n68842 = n68832 & ~n68841;
  assign n68843 = P2_P2_INSTQUEUE_REG_11__7_ & ~n68842;
  assign n68844 = n68388 & n68838;
  assign n68845 = n68391 & n68830;
  assign n68846 = ~n68844 & ~n68845;
  assign n68847 = n68397 & n68837;
  assign n68848 = n68846 & ~n68847;
  assign n68849 = n68386 & n68839;
  assign n68850 = n68348 & ~n68849;
  assign n68851 = ~n68835 & ~n68850;
  assign n68852 = n68406 & n68851;
  assign n68853 = ~n68843 & n68848;
  assign n12756 = n68852 | ~n68853;
  assign n68855 = P2_P2_INSTQUEUE_REG_11__6_ & ~n68842;
  assign n68856 = n68414 & n68838;
  assign n68857 = n68416 & n68830;
  assign n68858 = ~n68856 & ~n68857;
  assign n68859 = n68422 & n68837;
  assign n68860 = n68858 & ~n68859;
  assign n68861 = n68428 & n68851;
  assign n68862 = ~n68855 & n68860;
  assign n12761 = n68861 | ~n68862;
  assign n68864 = P2_P2_INSTQUEUE_REG_11__5_ & ~n68842;
  assign n68865 = n68436 & n68838;
  assign n68866 = n68438 & n68830;
  assign n68867 = ~n68865 & ~n68866;
  assign n68868 = n68444 & n68837;
  assign n68869 = n68867 & ~n68868;
  assign n68870 = n68450 & n68851;
  assign n68871 = ~n68864 & n68869;
  assign n12766 = n68870 | ~n68871;
  assign n68873 = P2_P2_INSTQUEUE_REG_11__4_ & ~n68842;
  assign n68874 = n68458 & n68838;
  assign n68875 = n68460 & n68830;
  assign n68876 = ~n68874 & ~n68875;
  assign n68877 = n68466 & n68837;
  assign n68878 = n68876 & ~n68877;
  assign n68879 = n68472 & n68851;
  assign n68880 = ~n68873 & n68878;
  assign n12771 = n68879 | ~n68880;
  assign n68882 = P2_P2_INSTQUEUE_REG_11__3_ & ~n68842;
  assign n68883 = n68480 & n68838;
  assign n68884 = n68482 & n68830;
  assign n68885 = ~n68883 & ~n68884;
  assign n68886 = n68488 & n68837;
  assign n68887 = n68885 & ~n68886;
  assign n68888 = n68494 & n68851;
  assign n68889 = ~n68882 & n68887;
  assign n12776 = n68888 | ~n68889;
  assign n68891 = P2_P2_INSTQUEUE_REG_11__2_ & ~n68842;
  assign n68892 = n68502 & n68838;
  assign n68893 = n68504 & n68830;
  assign n68894 = ~n68892 & ~n68893;
  assign n68895 = n68510 & n68837;
  assign n68896 = n68894 & ~n68895;
  assign n68897 = n68516 & n68851;
  assign n68898 = ~n68891 & n68896;
  assign n12781 = n68897 | ~n68898;
  assign n68900 = P2_P2_INSTQUEUE_REG_11__1_ & ~n68842;
  assign n68901 = n68524 & n68838;
  assign n68902 = n68526 & n68830;
  assign n68903 = ~n68901 & ~n68902;
  assign n68904 = n68532 & n68837;
  assign n68905 = n68903 & ~n68904;
  assign n68906 = n68538 & n68851;
  assign n68907 = ~n68900 & n68905;
  assign n12786 = n68906 | ~n68907;
  assign n68909 = P2_P2_INSTQUEUE_REG_11__0_ & ~n68842;
  assign n68910 = n68546 & n68838;
  assign n68911 = n68548 & n68830;
  assign n68912 = ~n68910 & ~n68911;
  assign n68913 = n68554 & n68837;
  assign n68914 = n68912 & ~n68913;
  assign n68915 = n68560 & n68851;
  assign n68916 = ~n68909 & n68914;
  assign n12791 = n68915 | ~n68916;
  assign n68918 = ~P2_P2_INSTQUEUEWR_ADDR_REG_2_ & ~P2_P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n68919 = n68564 & n68918;
  assign n68920 = P2_P2_STATE2_REG_3_ & ~n68919;
  assign n68921 = n68331 & ~n68920;
  assign n68922 = n68349 & n68833;
  assign n68923 = ~n68919 & ~n68922;
  assign n68924 = n68571 & n68836;
  assign n68925 = n68352 & n68368;
  assign n68926 = ~n68924 & ~n68925;
  assign n68927 = n68348 & ~n68926;
  assign n68928 = n68923 & ~n68927;
  assign n68929 = n68921 & ~n68928;
  assign n68930 = P2_P2_INSTQUEUE_REG_10__7_ & ~n68929;
  assign n68931 = n68388 & n68925;
  assign n68932 = n68391 & n68919;
  assign n68933 = ~n68931 & ~n68932;
  assign n68934 = n68397 & n68924;
  assign n68935 = n68933 & ~n68934;
  assign n68936 = n68386 & n68926;
  assign n68937 = n68348 & ~n68936;
  assign n68938 = ~n68923 & ~n68937;
  assign n68939 = n68406 & n68938;
  assign n68940 = ~n68930 & n68935;
  assign n12796 = n68939 | ~n68940;
  assign n68942 = P2_P2_INSTQUEUE_REG_10__6_ & ~n68929;
  assign n68943 = n68414 & n68925;
  assign n68944 = n68416 & n68919;
  assign n68945 = ~n68943 & ~n68944;
  assign n68946 = n68422 & n68924;
  assign n68947 = n68945 & ~n68946;
  assign n68948 = n68428 & n68938;
  assign n68949 = ~n68942 & n68947;
  assign n12801 = n68948 | ~n68949;
  assign n68951 = P2_P2_INSTQUEUE_REG_10__5_ & ~n68929;
  assign n68952 = n68436 & n68925;
  assign n68953 = n68438 & n68919;
  assign n68954 = ~n68952 & ~n68953;
  assign n68955 = n68444 & n68924;
  assign n68956 = n68954 & ~n68955;
  assign n68957 = n68450 & n68938;
  assign n68958 = ~n68951 & n68956;
  assign n12806 = n68957 | ~n68958;
  assign n68960 = P2_P2_INSTQUEUE_REG_10__4_ & ~n68929;
  assign n68961 = n68458 & n68925;
  assign n68962 = n68460 & n68919;
  assign n68963 = ~n68961 & ~n68962;
  assign n68964 = n68466 & n68924;
  assign n68965 = n68963 & ~n68964;
  assign n68966 = n68472 & n68938;
  assign n68967 = ~n68960 & n68965;
  assign n12811 = n68966 | ~n68967;
  assign n68969 = P2_P2_INSTQUEUE_REG_10__3_ & ~n68929;
  assign n68970 = n68480 & n68925;
  assign n68971 = n68482 & n68919;
  assign n68972 = ~n68970 & ~n68971;
  assign n68973 = n68488 & n68924;
  assign n68974 = n68972 & ~n68973;
  assign n68975 = n68494 & n68938;
  assign n68976 = ~n68969 & n68974;
  assign n12816 = n68975 | ~n68976;
  assign n68978 = P2_P2_INSTQUEUE_REG_10__2_ & ~n68929;
  assign n68979 = n68502 & n68925;
  assign n68980 = n68504 & n68919;
  assign n68981 = ~n68979 & ~n68980;
  assign n68982 = n68510 & n68924;
  assign n68983 = n68981 & ~n68982;
  assign n68984 = n68516 & n68938;
  assign n68985 = ~n68978 & n68983;
  assign n12821 = n68984 | ~n68985;
  assign n68987 = P2_P2_INSTQUEUE_REG_10__1_ & ~n68929;
  assign n68988 = n68524 & n68925;
  assign n68989 = n68526 & n68919;
  assign n68990 = ~n68988 & ~n68989;
  assign n68991 = n68532 & n68924;
  assign n68992 = n68990 & ~n68991;
  assign n68993 = n68538 & n68938;
  assign n68994 = ~n68987 & n68992;
  assign n12826 = n68993 | ~n68994;
  assign n68996 = P2_P2_INSTQUEUE_REG_10__0_ & ~n68929;
  assign n68997 = n68546 & n68925;
  assign n68998 = n68548 & n68919;
  assign n68999 = ~n68997 & ~n68998;
  assign n69000 = n68554 & n68924;
  assign n69001 = n68999 & ~n69000;
  assign n69002 = n68560 & n68938;
  assign n69003 = ~n68996 & n69001;
  assign n12831 = n69002 | ~n69003;
  assign n69005 = n68340 & n68829;
  assign n69006 = P2_P2_STATE2_REG_3_ & ~n69005;
  assign n69007 = n68331 & ~n69006;
  assign n69008 = n68350 & n68833;
  assign n69009 = ~n69005 & ~n69008;
  assign n69010 = n68659 & n68836;
  assign n69011 = n68353 & n68368;
  assign n69012 = ~n69010 & ~n69011;
  assign n69013 = n68348 & ~n69012;
  assign n69014 = n69009 & ~n69013;
  assign n69015 = n69007 & ~n69014;
  assign n69016 = P2_P2_INSTQUEUE_REG_9__7_ & ~n69015;
  assign n69017 = n68388 & n69011;
  assign n69018 = n68391 & n69005;
  assign n69019 = ~n69017 & ~n69018;
  assign n69020 = n68397 & n69010;
  assign n69021 = n69019 & ~n69020;
  assign n69022 = n68386 & n69012;
  assign n69023 = n68348 & ~n69022;
  assign n69024 = ~n69009 & ~n69023;
  assign n69025 = n68406 & n69024;
  assign n69026 = ~n69016 & n69021;
  assign n12836 = n69025 | ~n69026;
  assign n69028 = P2_P2_INSTQUEUE_REG_9__6_ & ~n69015;
  assign n69029 = n68414 & n69011;
  assign n69030 = n68416 & n69005;
  assign n69031 = ~n69029 & ~n69030;
  assign n69032 = n68422 & n69010;
  assign n69033 = n69031 & ~n69032;
  assign n69034 = n68428 & n69024;
  assign n69035 = ~n69028 & n69033;
  assign n12841 = n69034 | ~n69035;
  assign n69037 = P2_P2_INSTQUEUE_REG_9__5_ & ~n69015;
  assign n69038 = n68436 & n69011;
  assign n69039 = n68438 & n69005;
  assign n69040 = ~n69038 & ~n69039;
  assign n69041 = n68444 & n69010;
  assign n69042 = n69040 & ~n69041;
  assign n69043 = n68450 & n69024;
  assign n69044 = ~n69037 & n69042;
  assign n12846 = n69043 | ~n69044;
  assign n69046 = P2_P2_INSTQUEUE_REG_9__4_ & ~n69015;
  assign n69047 = n68458 & n69011;
  assign n69048 = n68460 & n69005;
  assign n69049 = ~n69047 & ~n69048;
  assign n69050 = n68466 & n69010;
  assign n69051 = n69049 & ~n69050;
  assign n69052 = n68472 & n69024;
  assign n69053 = ~n69046 & n69051;
  assign n12851 = n69052 | ~n69053;
  assign n69055 = P2_P2_INSTQUEUE_REG_9__3_ & ~n69015;
  assign n69056 = n68480 & n69011;
  assign n69057 = n68482 & n69005;
  assign n69058 = ~n69056 & ~n69057;
  assign n69059 = n68488 & n69010;
  assign n69060 = n69058 & ~n69059;
  assign n69061 = n68494 & n69024;
  assign n69062 = ~n69055 & n69060;
  assign n12856 = n69061 | ~n69062;
  assign n69064 = P2_P2_INSTQUEUE_REG_9__2_ & ~n69015;
  assign n69065 = n68502 & n69011;
  assign n69066 = n68504 & n69005;
  assign n69067 = ~n69065 & ~n69066;
  assign n69068 = n68510 & n69010;
  assign n69069 = n69067 & ~n69068;
  assign n69070 = n68516 & n69024;
  assign n69071 = ~n69064 & n69069;
  assign n12861 = n69070 | ~n69071;
  assign n69073 = P2_P2_INSTQUEUE_REG_9__1_ & ~n69015;
  assign n69074 = n68524 & n69011;
  assign n69075 = n68526 & n69005;
  assign n69076 = ~n69074 & ~n69075;
  assign n69077 = n68532 & n69010;
  assign n69078 = n69076 & ~n69077;
  assign n69079 = n68538 & n69024;
  assign n69080 = ~n69073 & n69078;
  assign n12866 = n69079 | ~n69080;
  assign n69082 = P2_P2_INSTQUEUE_REG_9__0_ & ~n69015;
  assign n69083 = n68546 & n69011;
  assign n69084 = n68548 & n69005;
  assign n69085 = ~n69083 & ~n69084;
  assign n69086 = n68554 & n69010;
  assign n69087 = n69085 & ~n69086;
  assign n69088 = n68560 & n69024;
  assign n69089 = ~n69082 & n69087;
  assign n12871 = n69088 | ~n69089;
  assign n69091 = n68741 & n68918;
  assign n69092 = P2_P2_STATE2_REG_3_ & ~n69091;
  assign n69093 = n68331 & ~n69092;
  assign n69094 = n68745 & n68836;
  assign n69095 = n68368 & n68747;
  assign n69096 = ~n69094 & ~n69095;
  assign n69097 = n68348 & ~n69096;
  assign n69098 = n68342 & n68833;
  assign n69099 = ~n69097 & ~n69098;
  assign n69100 = n69093 & ~n69099;
  assign n69101 = P2_P2_INSTQUEUE_REG_8__7_ & ~n69100;
  assign n69102 = n68388 & n69095;
  assign n69103 = n68391 & n69091;
  assign n69104 = ~n69102 & ~n69103;
  assign n69105 = n68397 & n69094;
  assign n69106 = n69104 & ~n69105;
  assign n69107 = n68386 & n69096;
  assign n69108 = n68348 & ~n69107;
  assign n69109 = n69098 & ~n69108;
  assign n69110 = n68406 & n69109;
  assign n69111 = ~n69101 & n69106;
  assign n12876 = n69110 | ~n69111;
  assign n69113 = P2_P2_INSTQUEUE_REG_8__6_ & ~n69100;
  assign n69114 = n68414 & n69095;
  assign n69115 = n68416 & n69091;
  assign n69116 = ~n69114 & ~n69115;
  assign n69117 = n68422 & n69094;
  assign n69118 = n69116 & ~n69117;
  assign n69119 = n68428 & n69109;
  assign n69120 = ~n69113 & n69118;
  assign n12881 = n69119 | ~n69120;
  assign n69122 = P2_P2_INSTQUEUE_REG_8__5_ & ~n69100;
  assign n69123 = n68436 & n69095;
  assign n69124 = n68438 & n69091;
  assign n69125 = ~n69123 & ~n69124;
  assign n69126 = n68444 & n69094;
  assign n69127 = n69125 & ~n69126;
  assign n69128 = n68450 & n69109;
  assign n69129 = ~n69122 & n69127;
  assign n12886 = n69128 | ~n69129;
  assign n69131 = P2_P2_INSTQUEUE_REG_8__4_ & ~n69100;
  assign n69132 = n68458 & n69095;
  assign n69133 = n68460 & n69091;
  assign n69134 = ~n69132 & ~n69133;
  assign n69135 = n68466 & n69094;
  assign n69136 = n69134 & ~n69135;
  assign n69137 = n68472 & n69109;
  assign n69138 = ~n69131 & n69136;
  assign n12891 = n69137 | ~n69138;
  assign n69140 = P2_P2_INSTQUEUE_REG_8__3_ & ~n69100;
  assign n69141 = n68480 & n69095;
  assign n69142 = n68482 & n69091;
  assign n69143 = ~n69141 & ~n69142;
  assign n69144 = n68488 & n69094;
  assign n69145 = n69143 & ~n69144;
  assign n69146 = n68494 & n69109;
  assign n69147 = ~n69140 & n69145;
  assign n12896 = n69146 | ~n69147;
  assign n69149 = P2_P2_INSTQUEUE_REG_8__2_ & ~n69100;
  assign n69150 = n68502 & n69095;
  assign n69151 = n68504 & n69091;
  assign n69152 = ~n69150 & ~n69151;
  assign n69153 = n68510 & n69094;
  assign n69154 = n69152 & ~n69153;
  assign n69155 = n68516 & n69109;
  assign n69156 = ~n69149 & n69154;
  assign n12901 = n69155 | ~n69156;
  assign n69158 = P2_P2_INSTQUEUE_REG_8__1_ & ~n69100;
  assign n69159 = n68524 & n69095;
  assign n69160 = n68526 & n69091;
  assign n69161 = ~n69159 & ~n69160;
  assign n69162 = n68532 & n69094;
  assign n69163 = n69161 & ~n69162;
  assign n69164 = n68538 & n69109;
  assign n69165 = ~n69158 & n69163;
  assign n12906 = n69164 | ~n69165;
  assign n69167 = P2_P2_INSTQUEUE_REG_8__0_ & ~n69100;
  assign n69168 = n68546 & n69095;
  assign n69169 = n68548 & n69091;
  assign n69170 = ~n69168 & ~n69169;
  assign n69171 = n68554 & n69094;
  assign n69172 = n69170 & ~n69171;
  assign n69173 = n68560 & n69109;
  assign n69174 = ~n69167 & n69172;
  assign n12911 = n69173 | ~n69174;
  assign n69176 = P2_P2_STATE2_REG_3_ & ~n68336;
  assign n69177 = n68331 & ~n69176;
  assign n69178 = ~n68336 & ~n68364;
  assign n69179 = ~n68362 & n68373;
  assign n69180 = n68355 & n69179;
  assign n69181 = ~n68372 & ~n69180;
  assign n69182 = n68348 & ~n69181;
  assign n69183 = n69178 & ~n69182;
  assign n69184 = n69177 & ~n69183;
  assign n69185 = P2_P2_INSTQUEUE_REG_7__7_ & ~n69184;
  assign n69186 = n68372 & n68388;
  assign n69187 = n68336 & n68391;
  assign n69188 = ~n69186 & ~n69187;
  assign n69189 = n68397 & n69180;
  assign n69190 = n69188 & ~n69189;
  assign n69191 = n68386 & n69181;
  assign n69192 = n68348 & ~n69191;
  assign n69193 = ~n69178 & ~n69192;
  assign n69194 = n68406 & n69193;
  assign n69195 = ~n69185 & n69190;
  assign n12916 = n69194 | ~n69195;
  assign n69197 = P2_P2_INSTQUEUE_REG_7__6_ & ~n69184;
  assign n69198 = n68372 & n68414;
  assign n69199 = n68336 & n68416;
  assign n69200 = ~n69198 & ~n69199;
  assign n69201 = n68422 & n69180;
  assign n69202 = n69200 & ~n69201;
  assign n69203 = n68428 & n69193;
  assign n69204 = ~n69197 & n69202;
  assign n12921 = n69203 | ~n69204;
  assign n69206 = P2_P2_INSTQUEUE_REG_7__5_ & ~n69184;
  assign n69207 = n68372 & n68436;
  assign n69208 = n68336 & n68438;
  assign n69209 = ~n69207 & ~n69208;
  assign n69210 = n68444 & n69180;
  assign n69211 = n69209 & ~n69210;
  assign n69212 = n68450 & n69193;
  assign n69213 = ~n69206 & n69211;
  assign n12926 = n69212 | ~n69213;
  assign n69215 = P2_P2_INSTQUEUE_REG_7__4_ & ~n69184;
  assign n69216 = n68372 & n68458;
  assign n69217 = n68336 & n68460;
  assign n69218 = ~n69216 & ~n69217;
  assign n69219 = n68466 & n69180;
  assign n69220 = n69218 & ~n69219;
  assign n69221 = n68472 & n69193;
  assign n69222 = ~n69215 & n69220;
  assign n12931 = n69221 | ~n69222;
  assign n69224 = P2_P2_INSTQUEUE_REG_7__3_ & ~n69184;
  assign n69225 = n68372 & n68480;
  assign n69226 = n68336 & n68482;
  assign n69227 = ~n69225 & ~n69226;
  assign n69228 = n68488 & n69180;
  assign n69229 = n69227 & ~n69228;
  assign n69230 = n68494 & n69193;
  assign n69231 = ~n69224 & n69229;
  assign n12936 = n69230 | ~n69231;
  assign n69233 = P2_P2_INSTQUEUE_REG_7__2_ & ~n69184;
  assign n69234 = n68372 & n68502;
  assign n69235 = n68336 & n68504;
  assign n69236 = ~n69234 & ~n69235;
  assign n69237 = n68510 & n69180;
  assign n69238 = n69236 & ~n69237;
  assign n69239 = n68516 & n69193;
  assign n69240 = ~n69233 & n69238;
  assign n12941 = n69239 | ~n69240;
  assign n69242 = P2_P2_INSTQUEUE_REG_7__1_ & ~n69184;
  assign n69243 = n68372 & n68524;
  assign n69244 = n68336 & n68526;
  assign n69245 = ~n69243 & ~n69244;
  assign n69246 = n68532 & n69180;
  assign n69247 = n69245 & ~n69246;
  assign n69248 = n68538 & n69193;
  assign n69249 = ~n69242 & n69247;
  assign n12946 = n69248 | ~n69249;
  assign n69251 = P2_P2_INSTQUEUE_REG_7__0_ & ~n69184;
  assign n69252 = n68372 & n68546;
  assign n69253 = n68336 & n68548;
  assign n69254 = ~n69252 & ~n69253;
  assign n69255 = n68554 & n69180;
  assign n69256 = n69254 & ~n69255;
  assign n69257 = n68560 & n69193;
  assign n69258 = ~n69251 & n69256;
  assign n12951 = n69257 | ~n69258;
  assign n69260 = ~P2_P2_INSTQUEUEWR_ADDR_REG_3_ & P2_P2_INSTQUEUEWR_ADDR_REG_1_;
  assign n69261 = n68565 & n69260;
  assign n69262 = P2_P2_STATE2_REG_3_ & ~n69261;
  assign n69263 = n68331 & ~n69262;
  assign n69264 = n68349 & n68363;
  assign n69265 = ~n69261 & ~n69264;
  assign n69266 = n68571 & n69179;
  assign n69267 = n68352 & n68371;
  assign n69268 = ~n69266 & ~n69267;
  assign n69269 = n68348 & ~n69268;
  assign n69270 = n69265 & ~n69269;
  assign n69271 = n69263 & ~n69270;
  assign n69272 = P2_P2_INSTQUEUE_REG_6__7_ & ~n69271;
  assign n69273 = n68388 & n69267;
  assign n69274 = n68391 & n69261;
  assign n69275 = ~n69273 & ~n69274;
  assign n69276 = n68397 & n69266;
  assign n69277 = n69275 & ~n69276;
  assign n69278 = n68386 & n69268;
  assign n69279 = n68348 & ~n69278;
  assign n69280 = ~n69265 & ~n69279;
  assign n69281 = n68406 & n69280;
  assign n69282 = ~n69272 & n69277;
  assign n12956 = n69281 | ~n69282;
  assign n69284 = P2_P2_INSTQUEUE_REG_6__6_ & ~n69271;
  assign n69285 = n68414 & n69267;
  assign n69286 = n68416 & n69261;
  assign n69287 = ~n69285 & ~n69286;
  assign n69288 = n68422 & n69266;
  assign n69289 = n69287 & ~n69288;
  assign n69290 = n68428 & n69280;
  assign n69291 = ~n69284 & n69289;
  assign n12961 = n69290 | ~n69291;
  assign n69293 = P2_P2_INSTQUEUE_REG_6__5_ & ~n69271;
  assign n69294 = n68436 & n69267;
  assign n69295 = n68438 & n69261;
  assign n69296 = ~n69294 & ~n69295;
  assign n69297 = n68444 & n69266;
  assign n69298 = n69296 & ~n69297;
  assign n69299 = n68450 & n69280;
  assign n69300 = ~n69293 & n69298;
  assign n12966 = n69299 | ~n69300;
  assign n69302 = P2_P2_INSTQUEUE_REG_6__4_ & ~n69271;
  assign n69303 = n68458 & n69267;
  assign n69304 = n68460 & n69261;
  assign n69305 = ~n69303 & ~n69304;
  assign n69306 = n68466 & n69266;
  assign n69307 = n69305 & ~n69306;
  assign n69308 = n68472 & n69280;
  assign n69309 = ~n69302 & n69307;
  assign n12971 = n69308 | ~n69309;
  assign n69311 = P2_P2_INSTQUEUE_REG_6__3_ & ~n69271;
  assign n69312 = n68480 & n69267;
  assign n69313 = n68482 & n69261;
  assign n69314 = ~n69312 & ~n69313;
  assign n69315 = n68488 & n69266;
  assign n69316 = n69314 & ~n69315;
  assign n69317 = n68494 & n69280;
  assign n69318 = ~n69311 & n69316;
  assign n12976 = n69317 | ~n69318;
  assign n69320 = P2_P2_INSTQUEUE_REG_6__2_ & ~n69271;
  assign n69321 = n68502 & n69267;
  assign n69322 = n68504 & n69261;
  assign n69323 = ~n69321 & ~n69322;
  assign n69324 = n68510 & n69266;
  assign n69325 = n69323 & ~n69324;
  assign n69326 = n68516 & n69280;
  assign n69327 = ~n69320 & n69325;
  assign n12981 = n69326 | ~n69327;
  assign n69329 = P2_P2_INSTQUEUE_REG_6__1_ & ~n69271;
  assign n69330 = n68524 & n69267;
  assign n69331 = n68526 & n69261;
  assign n69332 = ~n69330 & ~n69331;
  assign n69333 = n68532 & n69266;
  assign n69334 = n69332 & ~n69333;
  assign n69335 = n68538 & n69280;
  assign n69336 = ~n69329 & n69334;
  assign n12986 = n69335 | ~n69336;
  assign n69338 = P2_P2_INSTQUEUE_REG_6__0_ & ~n69271;
  assign n69339 = n68546 & n69267;
  assign n69340 = n68548 & n69261;
  assign n69341 = ~n69339 & ~n69340;
  assign n69342 = n68554 & n69266;
  assign n69343 = n69341 & ~n69342;
  assign n69344 = n68560 & n69280;
  assign n69345 = ~n69338 & n69343;
  assign n12991 = n69344 | ~n69345;
  assign n69347 = ~P2_P2_INSTQUEUEWR_ADDR_REG_3_ & P2_P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n69348 = n68340 & n69347;
  assign n69349 = P2_P2_STATE2_REG_3_ & ~n69348;
  assign n69350 = n68331 & ~n69349;
  assign n69351 = n68350 & n68363;
  assign n69352 = ~n69348 & ~n69351;
  assign n69353 = n68659 & n69179;
  assign n69354 = n68353 & n68371;
  assign n69355 = ~n69353 & ~n69354;
  assign n69356 = n68348 & ~n69355;
  assign n69357 = n69352 & ~n69356;
  assign n69358 = n69350 & ~n69357;
  assign n69359 = P2_P2_INSTQUEUE_REG_5__7_ & ~n69358;
  assign n69360 = n68388 & n69354;
  assign n69361 = n68391 & n69348;
  assign n69362 = ~n69360 & ~n69361;
  assign n69363 = n68397 & n69353;
  assign n69364 = n69362 & ~n69363;
  assign n69365 = n68386 & n69355;
  assign n69366 = n68348 & ~n69365;
  assign n69367 = ~n69352 & ~n69366;
  assign n69368 = n68406 & n69367;
  assign n69369 = ~n69359 & n69364;
  assign n12996 = n69368 | ~n69369;
  assign n69371 = P2_P2_INSTQUEUE_REG_5__6_ & ~n69358;
  assign n69372 = n68414 & n69354;
  assign n69373 = n68416 & n69348;
  assign n69374 = ~n69372 & ~n69373;
  assign n69375 = n68422 & n69353;
  assign n69376 = n69374 & ~n69375;
  assign n69377 = n68428 & n69367;
  assign n69378 = ~n69371 & n69376;
  assign n13001 = n69377 | ~n69378;
  assign n69380 = P2_P2_INSTQUEUE_REG_5__5_ & ~n69358;
  assign n69381 = n68436 & n69354;
  assign n69382 = n68438 & n69348;
  assign n69383 = ~n69381 & ~n69382;
  assign n69384 = n68444 & n69353;
  assign n69385 = n69383 & ~n69384;
  assign n69386 = n68450 & n69367;
  assign n69387 = ~n69380 & n69385;
  assign n13006 = n69386 | ~n69387;
  assign n69389 = P2_P2_INSTQUEUE_REG_5__4_ & ~n69358;
  assign n69390 = n68458 & n69354;
  assign n69391 = n68460 & n69348;
  assign n69392 = ~n69390 & ~n69391;
  assign n69393 = n68466 & n69353;
  assign n69394 = n69392 & ~n69393;
  assign n69395 = n68472 & n69367;
  assign n69396 = ~n69389 & n69394;
  assign n13011 = n69395 | ~n69396;
  assign n69398 = P2_P2_INSTQUEUE_REG_5__3_ & ~n69358;
  assign n69399 = n68480 & n69354;
  assign n69400 = n68482 & n69348;
  assign n69401 = ~n69399 & ~n69400;
  assign n69402 = n68488 & n69353;
  assign n69403 = n69401 & ~n69402;
  assign n69404 = n68494 & n69367;
  assign n69405 = ~n69398 & n69403;
  assign n13016 = n69404 | ~n69405;
  assign n69407 = P2_P2_INSTQUEUE_REG_5__2_ & ~n69358;
  assign n69408 = n68502 & n69354;
  assign n69409 = n68504 & n69348;
  assign n69410 = ~n69408 & ~n69409;
  assign n69411 = n68510 & n69353;
  assign n69412 = n69410 & ~n69411;
  assign n69413 = n68516 & n69367;
  assign n69414 = ~n69407 & n69412;
  assign n13021 = n69413 | ~n69414;
  assign n69416 = P2_P2_INSTQUEUE_REG_5__1_ & ~n69358;
  assign n69417 = n68524 & n69354;
  assign n69418 = n68526 & n69348;
  assign n69419 = ~n69417 & ~n69418;
  assign n69420 = n68532 & n69353;
  assign n69421 = n69419 & ~n69420;
  assign n69422 = n68538 & n69367;
  assign n69423 = ~n69416 & n69421;
  assign n13026 = n69422 | ~n69423;
  assign n69425 = P2_P2_INSTQUEUE_REG_5__0_ & ~n69358;
  assign n69426 = n68546 & n69354;
  assign n69427 = n68548 & n69348;
  assign n69428 = ~n69426 & ~n69427;
  assign n69429 = n68554 & n69353;
  assign n69430 = n69428 & ~n69429;
  assign n69431 = n68560 & n69367;
  assign n69432 = ~n69425 & n69430;
  assign n13031 = n69431 | ~n69432;
  assign n69434 = n68371 & n68747;
  assign n69435 = n68388 & n69434;
  assign n69436 = ~P2_P2_INSTQUEUEWR_ADDR_REG_3_ & ~P2_P2_INSTQUEUEWR_ADDR_REG_1_;
  assign n69437 = n68565 & n69436;
  assign n69438 = n68391 & n69437;
  assign n69439 = n68348 & ~n68386;
  assign n69440 = n68342 & n68363;
  assign n69441 = ~n69439 & n69440;
  assign n69442 = n68406 & n69441;
  assign n69443 = ~n69435 & ~n69438;
  assign n69444 = ~n69442 & n69443;
  assign n69445 = n68745 & n69179;
  assign n69446 = n68397 & n69445;
  assign n69447 = n69444 & ~n69446;
  assign n69448 = P2_P2_STATE2_REG_3_ & ~n69437;
  assign n69449 = n68331 & ~n69448;
  assign n69450 = ~n69434 & ~n69445;
  assign n69451 = n68348 & ~n69450;
  assign n69452 = ~n69440 & ~n69451;
  assign n69453 = n69449 & ~n69452;
  assign n69454 = P2_P2_INSTQUEUE_REG_4__7_ & ~n69453;
  assign n13036 = ~n69447 | n69454;
  assign n69456 = n68414 & n69434;
  assign n69457 = n68416 & n69437;
  assign n69458 = n68428 & n69441;
  assign n69459 = ~n69456 & ~n69457;
  assign n69460 = ~n69458 & n69459;
  assign n69461 = n68422 & n69445;
  assign n69462 = n69460 & ~n69461;
  assign n69463 = P2_P2_INSTQUEUE_REG_4__6_ & ~n69453;
  assign n13041 = ~n69462 | n69463;
  assign n69465 = n68436 & n69434;
  assign n69466 = n68438 & n69437;
  assign n69467 = n68450 & n69441;
  assign n69468 = ~n69465 & ~n69466;
  assign n69469 = ~n69467 & n69468;
  assign n69470 = n68444 & n69445;
  assign n69471 = n69469 & ~n69470;
  assign n69472 = P2_P2_INSTQUEUE_REG_4__5_ & ~n69453;
  assign n13046 = ~n69471 | n69472;
  assign n69474 = n68458 & n69434;
  assign n69475 = n68460 & n69437;
  assign n69476 = n68472 & n69441;
  assign n69477 = ~n69474 & ~n69475;
  assign n69478 = ~n69476 & n69477;
  assign n69479 = n68466 & n69445;
  assign n69480 = n69478 & ~n69479;
  assign n69481 = P2_P2_INSTQUEUE_REG_4__4_ & ~n69453;
  assign n13051 = ~n69480 | n69481;
  assign n69483 = n68480 & n69434;
  assign n69484 = n68482 & n69437;
  assign n69485 = n68494 & n69441;
  assign n69486 = ~n69483 & ~n69484;
  assign n69487 = ~n69485 & n69486;
  assign n69488 = n68488 & n69445;
  assign n69489 = n69487 & ~n69488;
  assign n69490 = P2_P2_INSTQUEUE_REG_4__3_ & ~n69453;
  assign n13056 = ~n69489 | n69490;
  assign n69492 = n68502 & n69434;
  assign n69493 = n68504 & n69437;
  assign n69494 = n68516 & n69441;
  assign n69495 = ~n69492 & ~n69493;
  assign n69496 = ~n69494 & n69495;
  assign n69497 = n68510 & n69445;
  assign n69498 = n69496 & ~n69497;
  assign n69499 = P2_P2_INSTQUEUE_REG_4__2_ & ~n69453;
  assign n13061 = ~n69498 | n69499;
  assign n69501 = n68524 & n69434;
  assign n69502 = n68526 & n69437;
  assign n69503 = n68538 & n69441;
  assign n69504 = ~n69501 & ~n69502;
  assign n69505 = ~n69503 & n69504;
  assign n69506 = n68532 & n69445;
  assign n69507 = n69505 & ~n69506;
  assign n69508 = P2_P2_INSTQUEUE_REG_4__1_ & ~n69453;
  assign n13066 = ~n69507 | n69508;
  assign n69510 = n68546 & n69434;
  assign n69511 = n68548 & n69437;
  assign n69512 = n68560 & n69441;
  assign n69513 = ~n69510 & ~n69511;
  assign n69514 = ~n69512 & n69513;
  assign n69515 = n68554 & n69445;
  assign n69516 = n69514 & ~n69515;
  assign n69517 = P2_P2_INSTQUEUE_REG_4__0_ & ~n69453;
  assign n13071 = ~n69516 | n69517;
  assign n69519 = n68358 & n68367;
  assign n69520 = n68359 & n69519;
  assign n69521 = n68388 & n69520;
  assign n69522 = ~P2_P2_INSTQUEUEWR_ADDR_REG_3_ & ~P2_P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n69523 = n68324 & n69522;
  assign n69524 = n68391 & n69523;
  assign n69525 = n68335 & n68338;
  assign n69526 = n68343 & n69525;
  assign n69527 = ~n69523 & ~n69526;
  assign n69528 = ~n69439 & ~n69527;
  assign n69529 = n68406 & n69528;
  assign n69530 = ~n69521 & ~n69524;
  assign n69531 = ~n69529 & n69530;
  assign n69532 = n68362 & n68373;
  assign n69533 = n68355 & n69532;
  assign n69534 = n68397 & n69533;
  assign n69535 = n69531 & ~n69534;
  assign n69536 = P2_P2_STATE2_REG_3_ & ~n69523;
  assign n69537 = n68331 & ~n69536;
  assign n69538 = ~n69520 & ~n69533;
  assign n69539 = n68348 & ~n69538;
  assign n69540 = n69527 & ~n69539;
  assign n69541 = n69537 & ~n69540;
  assign n69542 = P2_P2_INSTQUEUE_REG_3__7_ & ~n69541;
  assign n13076 = ~n69535 | n69542;
  assign n69544 = n68414 & n69520;
  assign n69545 = n68416 & n69523;
  assign n69546 = n68428 & n69528;
  assign n69547 = ~n69544 & ~n69545;
  assign n69548 = ~n69546 & n69547;
  assign n69549 = n68422 & n69533;
  assign n69550 = n69548 & ~n69549;
  assign n69551 = P2_P2_INSTQUEUE_REG_3__6_ & ~n69541;
  assign n13081 = ~n69550 | n69551;
  assign n69553 = n68436 & n69520;
  assign n69554 = n68438 & n69523;
  assign n69555 = n68450 & n69528;
  assign n69556 = ~n69553 & ~n69554;
  assign n69557 = ~n69555 & n69556;
  assign n69558 = n68444 & n69533;
  assign n69559 = n69557 & ~n69558;
  assign n69560 = P2_P2_INSTQUEUE_REG_3__5_ & ~n69541;
  assign n13086 = ~n69559 | n69560;
  assign n69562 = n68458 & n69520;
  assign n69563 = n68460 & n69523;
  assign n69564 = n68472 & n69528;
  assign n69565 = ~n69562 & ~n69563;
  assign n69566 = ~n69564 & n69565;
  assign n69567 = n68466 & n69533;
  assign n69568 = n69566 & ~n69567;
  assign n69569 = P2_P2_INSTQUEUE_REG_3__4_ & ~n69541;
  assign n13091 = ~n69568 | n69569;
  assign n69571 = n68480 & n69520;
  assign n69572 = n68482 & n69523;
  assign n69573 = n68494 & n69528;
  assign n69574 = ~n69571 & ~n69572;
  assign n69575 = ~n69573 & n69574;
  assign n69576 = n68488 & n69533;
  assign n69577 = n69575 & ~n69576;
  assign n69578 = P2_P2_INSTQUEUE_REG_3__3_ & ~n69541;
  assign n13096 = ~n69577 | n69578;
  assign n69580 = n68502 & n69520;
  assign n69581 = n68504 & n69523;
  assign n69582 = n68516 & n69528;
  assign n69583 = ~n69580 & ~n69581;
  assign n69584 = ~n69582 & n69583;
  assign n69585 = n68510 & n69533;
  assign n69586 = n69584 & ~n69585;
  assign n69587 = P2_P2_INSTQUEUE_REG_3__2_ & ~n69541;
  assign n13101 = ~n69586 | n69587;
  assign n69589 = n68524 & n69520;
  assign n69590 = n68526 & n69523;
  assign n69591 = n68538 & n69528;
  assign n69592 = ~n69589 & ~n69590;
  assign n69593 = ~n69591 & n69592;
  assign n69594 = n68532 & n69533;
  assign n69595 = n69593 & ~n69594;
  assign n69596 = P2_P2_INSTQUEUE_REG_3__1_ & ~n69541;
  assign n13106 = ~n69595 | n69596;
  assign n69598 = n68546 & n69520;
  assign n69599 = n68548 & n69523;
  assign n69600 = n68560 & n69528;
  assign n69601 = ~n69598 & ~n69599;
  assign n69602 = ~n69600 & n69601;
  assign n69603 = n68554 & n69533;
  assign n69604 = n69602 & ~n69603;
  assign n69605 = P2_P2_INSTQUEUE_REG_3__0_ & ~n69541;
  assign n13111 = ~n69604 | n69605;
  assign n69607 = n68352 & n69519;
  assign n69608 = n68388 & n69607;
  assign n69609 = n68918 & n69260;
  assign n69610 = n68391 & n69609;
  assign n69611 = n68349 & n69525;
  assign n69612 = ~n69609 & ~n69611;
  assign n69613 = ~n69439 & ~n69612;
  assign n69614 = n68406 & n69613;
  assign n69615 = ~n69608 & ~n69610;
  assign n69616 = ~n69614 & n69615;
  assign n69617 = n68571 & n69532;
  assign n69618 = n68397 & n69617;
  assign n69619 = n69616 & ~n69618;
  assign n69620 = P2_P2_STATE2_REG_3_ & ~n69609;
  assign n69621 = n68331 & ~n69620;
  assign n69622 = ~n69607 & ~n69617;
  assign n69623 = n68348 & ~n69622;
  assign n69624 = n69612 & ~n69623;
  assign n69625 = n69621 & ~n69624;
  assign n69626 = P2_P2_INSTQUEUE_REG_2__7_ & ~n69625;
  assign n13116 = ~n69619 | n69626;
  assign n69628 = n68414 & n69607;
  assign n69629 = n68416 & n69609;
  assign n69630 = n68428 & n69613;
  assign n69631 = ~n69628 & ~n69629;
  assign n69632 = ~n69630 & n69631;
  assign n69633 = n68422 & n69617;
  assign n69634 = n69632 & ~n69633;
  assign n69635 = P2_P2_INSTQUEUE_REG_2__6_ & ~n69625;
  assign n13121 = ~n69634 | n69635;
  assign n69637 = n68436 & n69607;
  assign n69638 = n68438 & n69609;
  assign n69639 = n68450 & n69613;
  assign n69640 = ~n69637 & ~n69638;
  assign n69641 = ~n69639 & n69640;
  assign n69642 = n68444 & n69617;
  assign n69643 = n69641 & ~n69642;
  assign n69644 = P2_P2_INSTQUEUE_REG_2__5_ & ~n69625;
  assign n13126 = ~n69643 | n69644;
  assign n69646 = n68458 & n69607;
  assign n69647 = n68460 & n69609;
  assign n69648 = n68472 & n69613;
  assign n69649 = ~n69646 & ~n69647;
  assign n69650 = ~n69648 & n69649;
  assign n69651 = n68466 & n69617;
  assign n69652 = n69650 & ~n69651;
  assign n69653 = P2_P2_INSTQUEUE_REG_2__4_ & ~n69625;
  assign n13131 = ~n69652 | n69653;
  assign n69655 = n68480 & n69607;
  assign n69656 = n68482 & n69609;
  assign n69657 = n68494 & n69613;
  assign n69658 = ~n69655 & ~n69656;
  assign n69659 = ~n69657 & n69658;
  assign n69660 = n68488 & n69617;
  assign n69661 = n69659 & ~n69660;
  assign n69662 = P2_P2_INSTQUEUE_REG_2__3_ & ~n69625;
  assign n13136 = ~n69661 | n69662;
  assign n69664 = n68502 & n69607;
  assign n69665 = n68504 & n69609;
  assign n69666 = n68516 & n69613;
  assign n69667 = ~n69664 & ~n69665;
  assign n69668 = ~n69666 & n69667;
  assign n69669 = n68510 & n69617;
  assign n69670 = n69668 & ~n69669;
  assign n69671 = P2_P2_INSTQUEUE_REG_2__2_ & ~n69625;
  assign n13141 = ~n69670 | n69671;
  assign n69673 = n68524 & n69607;
  assign n69674 = n68526 & n69609;
  assign n69675 = n68538 & n69613;
  assign n69676 = ~n69673 & ~n69674;
  assign n69677 = ~n69675 & n69676;
  assign n69678 = n68532 & n69617;
  assign n69679 = n69677 & ~n69678;
  assign n69680 = P2_P2_INSTQUEUE_REG_2__1_ & ~n69625;
  assign n13146 = ~n69679 | n69680;
  assign n69682 = n68546 & n69607;
  assign n69683 = n68548 & n69609;
  assign n69684 = n68560 & n69613;
  assign n69685 = ~n69682 & ~n69683;
  assign n69686 = ~n69684 & n69685;
  assign n69687 = n68554 & n69617;
  assign n69688 = n69686 & ~n69687;
  assign n69689 = P2_P2_INSTQUEUE_REG_2__0_ & ~n69625;
  assign n13151 = ~n69688 | n69689;
  assign n69691 = n68353 & n69519;
  assign n69692 = n68388 & n69691;
  assign n69693 = n68340 & n69522;
  assign n69694 = n68391 & n69693;
  assign n69695 = n68350 & n69525;
  assign n69696 = ~n69693 & ~n69695;
  assign n69697 = ~n69439 & ~n69696;
  assign n69698 = n68406 & n69697;
  assign n69699 = ~n69692 & ~n69694;
  assign n69700 = ~n69698 & n69699;
  assign n69701 = n68659 & n69532;
  assign n69702 = n68397 & n69701;
  assign n69703 = n69700 & ~n69702;
  assign n69704 = P2_P2_STATE2_REG_3_ & ~n69693;
  assign n69705 = n68331 & ~n69704;
  assign n69706 = ~n69691 & ~n69701;
  assign n69707 = n68348 & ~n69706;
  assign n69708 = n69696 & ~n69707;
  assign n69709 = n69705 & ~n69708;
  assign n69710 = P2_P2_INSTQUEUE_REG_1__7_ & ~n69709;
  assign n13156 = ~n69703 | n69710;
  assign n69712 = n68414 & n69691;
  assign n69713 = n68416 & n69693;
  assign n69714 = n68428 & n69697;
  assign n69715 = ~n69712 & ~n69713;
  assign n69716 = ~n69714 & n69715;
  assign n69717 = n68422 & n69701;
  assign n69718 = n69716 & ~n69717;
  assign n69719 = P2_P2_INSTQUEUE_REG_1__6_ & ~n69709;
  assign n13161 = ~n69718 | n69719;
  assign n69721 = n68436 & n69691;
  assign n69722 = n68438 & n69693;
  assign n69723 = n68450 & n69697;
  assign n69724 = ~n69721 & ~n69722;
  assign n69725 = ~n69723 & n69724;
  assign n69726 = n68444 & n69701;
  assign n69727 = n69725 & ~n69726;
  assign n69728 = P2_P2_INSTQUEUE_REG_1__5_ & ~n69709;
  assign n13166 = ~n69727 | n69728;
  assign n69730 = n68458 & n69691;
  assign n69731 = n68460 & n69693;
  assign n69732 = n68472 & n69697;
  assign n69733 = ~n69730 & ~n69731;
  assign n69734 = ~n69732 & n69733;
  assign n69735 = n68466 & n69701;
  assign n69736 = n69734 & ~n69735;
  assign n69737 = P2_P2_INSTQUEUE_REG_1__4_ & ~n69709;
  assign n13171 = ~n69736 | n69737;
  assign n69739 = n68480 & n69691;
  assign n69740 = n68482 & n69693;
  assign n69741 = n68494 & n69697;
  assign n69742 = ~n69739 & ~n69740;
  assign n69743 = ~n69741 & n69742;
  assign n69744 = n68488 & n69701;
  assign n69745 = n69743 & ~n69744;
  assign n69746 = P2_P2_INSTQUEUE_REG_1__3_ & ~n69709;
  assign n13176 = ~n69745 | n69746;
  assign n69748 = n68502 & n69691;
  assign n69749 = n68504 & n69693;
  assign n69750 = n68516 & n69697;
  assign n69751 = ~n69748 & ~n69749;
  assign n69752 = ~n69750 & n69751;
  assign n69753 = n68510 & n69701;
  assign n69754 = n69752 & ~n69753;
  assign n69755 = P2_P2_INSTQUEUE_REG_1__2_ & ~n69709;
  assign n13181 = ~n69754 | n69755;
  assign n69757 = n68524 & n69691;
  assign n69758 = n68526 & n69693;
  assign n69759 = n68538 & n69697;
  assign n69760 = ~n69757 & ~n69758;
  assign n69761 = ~n69759 & n69760;
  assign n69762 = n68532 & n69701;
  assign n69763 = n69761 & ~n69762;
  assign n69764 = P2_P2_INSTQUEUE_REG_1__1_ & ~n69709;
  assign n13186 = ~n69763 | n69764;
  assign n69766 = n68546 & n69691;
  assign n69767 = n68548 & n69693;
  assign n69768 = n68560 & n69697;
  assign n69769 = ~n69766 & ~n69767;
  assign n69770 = ~n69768 & n69769;
  assign n69771 = n68554 & n69701;
  assign n69772 = n69770 & ~n69771;
  assign n69773 = P2_P2_INSTQUEUE_REG_1__0_ & ~n69709;
  assign n13191 = ~n69772 | n69773;
  assign n69775 = n68747 & n69519;
  assign n69776 = n68388 & n69775;
  assign n69777 = n68918 & n69436;
  assign n69778 = n68391 & n69777;
  assign n69779 = n68342 & n69525;
  assign n69780 = ~n69439 & n69779;
  assign n69781 = n68406 & n69780;
  assign n69782 = ~n69776 & ~n69778;
  assign n69783 = ~n69781 & n69782;
  assign n69784 = n68745 & n69532;
  assign n69785 = n68397 & n69784;
  assign n69786 = n69783 & ~n69785;
  assign n69787 = P2_P2_STATE2_REG_3_ & ~n69777;
  assign n69788 = n68331 & ~n69787;
  assign n69789 = ~n69775 & ~n69784;
  assign n69790 = n68348 & ~n69789;
  assign n69791 = ~n69779 & ~n69790;
  assign n69792 = n69788 & ~n69791;
  assign n69793 = P2_P2_INSTQUEUE_REG_0__7_ & ~n69792;
  assign n13196 = ~n69786 | n69793;
  assign n69795 = n68414 & n69775;
  assign n69796 = n68416 & n69777;
  assign n69797 = n68428 & n69780;
  assign n69798 = ~n69795 & ~n69796;
  assign n69799 = ~n69797 & n69798;
  assign n69800 = n68422 & n69784;
  assign n69801 = n69799 & ~n69800;
  assign n69802 = P2_P2_INSTQUEUE_REG_0__6_ & ~n69792;
  assign n13201 = ~n69801 | n69802;
  assign n69804 = n68436 & n69775;
  assign n69805 = n68438 & n69777;
  assign n69806 = n68450 & n69780;
  assign n69807 = ~n69804 & ~n69805;
  assign n69808 = ~n69806 & n69807;
  assign n69809 = n68444 & n69784;
  assign n69810 = n69808 & ~n69809;
  assign n69811 = P2_P2_INSTQUEUE_REG_0__5_ & ~n69792;
  assign n13206 = ~n69810 | n69811;
  assign n69813 = n68458 & n69775;
  assign n69814 = n68460 & n69777;
  assign n69815 = n68472 & n69780;
  assign n69816 = ~n69813 & ~n69814;
  assign n69817 = ~n69815 & n69816;
  assign n69818 = n68466 & n69784;
  assign n69819 = n69817 & ~n69818;
  assign n69820 = P2_P2_INSTQUEUE_REG_0__4_ & ~n69792;
  assign n13211 = ~n69819 | n69820;
  assign n69822 = n68480 & n69775;
  assign n69823 = n68482 & n69777;
  assign n69824 = n68494 & n69780;
  assign n69825 = ~n69822 & ~n69823;
  assign n69826 = ~n69824 & n69825;
  assign n69827 = n68488 & n69784;
  assign n69828 = n69826 & ~n69827;
  assign n69829 = P2_P2_INSTQUEUE_REG_0__3_ & ~n69792;
  assign n13216 = ~n69828 | n69829;
  assign n69831 = n68502 & n69775;
  assign n69832 = n68504 & n69777;
  assign n69833 = n68516 & n69780;
  assign n69834 = ~n69831 & ~n69832;
  assign n69835 = ~n69833 & n69834;
  assign n69836 = n68510 & n69784;
  assign n69837 = n69835 & ~n69836;
  assign n69838 = P2_P2_INSTQUEUE_REG_0__2_ & ~n69792;
  assign n13221 = ~n69837 | n69838;
  assign n69840 = n68524 & n69775;
  assign n69841 = n68526 & n69777;
  assign n69842 = n68538 & n69780;
  assign n69843 = ~n69840 & ~n69841;
  assign n69844 = ~n69842 & n69843;
  assign n69845 = n68532 & n69784;
  assign n69846 = n69844 & ~n69845;
  assign n69847 = P2_P2_INSTQUEUE_REG_0__1_ & ~n69792;
  assign n13226 = ~n69846 | n69847;
  assign n69849 = n68546 & n69775;
  assign n69850 = n68548 & n69777;
  assign n69851 = n68560 & n69780;
  assign n69852 = ~n69849 & ~n69850;
  assign n69853 = ~n69851 & n69852;
  assign n69854 = n68554 & n69784;
  assign n69855 = n69853 & ~n69854;
  assign n69856 = P2_P2_INSTQUEUE_REG_0__0_ & ~n69792;
  assign n13231 = ~n69855 | n69856;
  assign n69858 = P2_P2_STATE2_REG_3_ & ~P2_P2_STATE2_REG_0_;
  assign n69859 = P2_P2_STATE2_REG_0_ & P2_P2_FLUSH_REG;
  assign n69860 = n67626 & n69859;
  assign n69861 = ~n69858 & ~n69860;
  assign n69862 = ~n68158 & n68268;
  assign n69863 = n69861 & ~n69862;
  assign n69864 = P2_P2_INSTQUEUERD_ADDR_REG_4_ & n69863;
  assign n69865 = ~n68201 & n68274;
  assign n69866 = n67993 & n69865;
  assign n69867 = ~n69863 & n69866;
  assign n13236 = n69864 | n69867;
  assign n69869 = ~n68192 & n68274;
  assign n69870 = ~n67665 & ~n68165;
  assign n69871 = n68283 & ~n69870;
  assign n69872 = ~n69869 & ~n69871;
  assign n69873 = ~n69863 & ~n69872;
  assign n69874 = P2_P2_INSTQUEUERD_ADDR_REG_3_ & n69863;
  assign n13241 = n69873 | n69874;
  assign n69876 = ~n68116 & n68283;
  assign n69877 = P2_P2_STATE2_REG_1_ & ~n68290;
  assign n69878 = ~n68299 & n69877;
  assign n69879 = ~n69876 & ~n69878;
  assign n69880 = ~n68132 & n68274;
  assign n69881 = n69879 & ~n69880;
  assign n69882 = ~n69863 & ~n69881;
  assign n69883 = P2_P2_INSTQUEUERD_ADDR_REG_2_ & n69863;
  assign n13246 = n69882 | n69883;
  assign n69885 = n68228 & n68283;
  assign n69886 = n68299 & n69877;
  assign n69887 = ~n69885 & ~n69886;
  assign n69888 = ~n68233 & n68274;
  assign n69889 = n69887 & ~n69888;
  assign n69890 = ~n69863 & ~n69889;
  assign n69891 = P2_P2_INSTQUEUERD_ADDR_REG_1_ & n69863;
  assign n13251 = n69890 | n69891;
  assign n69893 = P2_P2_STATE2_REG_1_ & n68290;
  assign n69894 = ~P2_P2_INSTQUEUERD_ADDR_REG_0_ & n68283;
  assign n69895 = ~n69893 & ~n69894;
  assign n69896 = ~n68219 & n68274;
  assign n69897 = n69895 & ~n69896;
  assign n69898 = ~n69863 & ~n69897;
  assign n69899 = P2_P2_INSTQUEUERD_ADDR_REG_0_ & n69863;
  assign n13256 = n69898 | n69899;
  assign n69901 = P2_P2_STATE2_REG_0_ & n67626;
  assign n69902 = ~n68313 & n69901;
  assign n69903 = ~n68331 & ~n69860;
  assign n69904 = ~n69902 & n69903;
  assign n13261 = P2_P2_INSTQUEUEWR_ADDR_REG_4_ & n69904;
  assign n69906 = P2_P2_STATE2_REG_3_ & ~n68325;
  assign n69907 = ~n69904 & ~n69906;
  assign n69908 = P2_P2_INSTQUEUEWR_ADDR_REG_3_ & ~n69907;
  assign n69909 = ~n68274 & ~n68347;
  assign n69910 = ~n68367 & ~n69909;
  assign n69911 = P2_P2_STATE2_REG_3_ & n68336;
  assign n69912 = ~n69910 & ~n69911;
  assign n69913 = n68355 & ~n68362;
  assign n69914 = ~n68373 & ~n69913;
  assign n69915 = ~n69180 & ~n69914;
  assign n69916 = n68386 & ~n69915;
  assign n69917 = n69912 & ~n69916;
  assign n69918 = ~n69904 & ~n69917;
  assign n13266 = n69908 | n69918;
  assign n69920 = ~n68358 & ~n69909;
  assign n69921 = P2_P2_STATE2_REG_3_ & ~P2_P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n69922 = n68324 & n69921;
  assign n69923 = ~n69920 & ~n69922;
  assign n69924 = ~n68355 & ~n68362;
  assign n69925 = n68355 & n68362;
  assign n69926 = ~n69924 & ~n69925;
  assign n69927 = n68386 & ~n69926;
  assign n69928 = n69923 & ~n69927;
  assign n69929 = ~n69904 & ~n69928;
  assign n69930 = P2_P2_STATE2_REG_3_ & ~n68324;
  assign n69931 = ~n69904 & ~n69930;
  assign n69932 = P2_P2_INSTQUEUEWR_ADDR_REG_2_ & ~n69931;
  assign n13271 = n69929 | n69932;
  assign n69934 = ~n68351 & ~n69909;
  assign n69935 = P2_P2_STATE2_REG_3_ & ~P2_P2_INSTQUEUEWR_ADDR_REG_1_;
  assign n69936 = ~n68354 & n68386;
  assign n69937 = ~n69935 & ~n69936;
  assign n69938 = P2_P2_INSTQUEUEWR_ADDR_REG_0_ & ~n69937;
  assign n69939 = n68386 & n68659;
  assign n69940 = ~n69934 & ~n69938;
  assign n69941 = ~n69939 & n69940;
  assign n69942 = ~n69904 & ~n69941;
  assign n69943 = P2_P2_STATE2_REG_3_ & ~P2_P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n69944 = ~n69904 & ~n69943;
  assign n69945 = P2_P2_INSTQUEUEWR_ADDR_REG_1_ & ~n69944;
  assign n13276 = n69942 | n69945;
  assign n69947 = ~n68274 & ~n68346;
  assign n69948 = ~n69904 & n69947;
  assign n69949 = P2_P2_INSTQUEUEWR_ADDR_REG_0_ & ~n69948;
  assign n69950 = ~n68314 & ~n69943;
  assign n69951 = ~n69904 & ~n69950;
  assign n13281 = n69949 | n69951;
  assign n69953 = ~P2_P2_STATE2_REG_1_ & n68346;
  assign n69954 = ~P2_P2_STATE2_REG_0_ & n69953;
  assign n69955 = n67922 & n67966;
  assign n69956 = ~n67754 & ~n67913;
  assign n69957 = n68011 & n69956;
  assign n69958 = n67920 & n67966;
  assign n69959 = ~n68150 & ~n69957;
  assign n69960 = ~n69958 & n69959;
  assign n69961 = n67971 & n68019;
  assign n69962 = n67723 & n67918;
  assign n69963 = n67966 & n69962;
  assign n69964 = ~n69961 & ~n69963;
  assign n69965 = n67882 & ~n69964;
  assign n69966 = ~n67722 & n68025;
  assign n69967 = ~n67541 & n67691;
  assign n69968 = n67966 & n69967;
  assign n69969 = ~n69966 & ~n69968;
  assign n69970 = ~n67882 & ~n69969;
  assign n69971 = n67913 & n68011;
  assign n69972 = ~n69965 & ~n69970;
  assign n69973 = ~n69971 & n69972;
  assign n69974 = n67847 & ~n69973;
  assign n69975 = n68142 & ~n69955;
  assign n69976 = n69960 & n69975;
  assign n69977 = ~n69974 & n69976;
  assign n69978 = n68268 & ~n69977;
  assign n69979 = ~n69954 & ~n69978;
  assign n69980 = P2_P2_STATE2_REG_2_ & ~n69979;
  assign n69981 = ~P2_P2_INSTADDRPOINTER_REG_0_ & n68212;
  assign n69982 = ~P2_P2_INSTADDRPOINTER_REG_0_ & n68055;
  assign n69983 = ~n69981 & ~n69982;
  assign n69984 = ~P2_P2_INSTADDRPOINTER_REG_0_ & ~n68102;
  assign n69985 = P2_P2_INSTADDRPOINTER_REG_0_ & n68173;
  assign n69986 = P2_P2_INSTADDRPOINTER_REG_0_ & n68174;
  assign n69987 = n67914 & n68045;
  assign n69988 = n68051 & n69987;
  assign n69989 = ~P2_P2_INSTADDRPOINTER_REG_0_ & n69988;
  assign n69990 = n67991 & n68045;
  assign n69991 = n68051 & n69990;
  assign n69992 = ~P2_P2_INSTADDRPOINTER_REG_0_ & n69991;
  assign n69993 = ~n69989 & ~n69992;
  assign n69994 = P2_P2_INSTADDRPOINTER_REG_0_ & n67989;
  assign n69995 = n69993 & ~n69994;
  assign n69996 = n68116 & n69870;
  assign n69997 = P2_P2_INSTQUEUERD_ADDR_REG_0_ & ~n68228;
  assign n69998 = n69996 & n69997;
  assign n69999 = P2_P2_INSTQUEUE_REG_0__0_ & n69998;
  assign n70000 = ~P2_P2_INSTQUEUERD_ADDR_REG_0_ & ~n68228;
  assign n70001 = n69996 & n70000;
  assign n70002 = P2_P2_INSTQUEUE_REG_1__0_ & n70001;
  assign n70003 = P2_P2_INSTQUEUERD_ADDR_REG_0_ & n68228;
  assign n70004 = n69996 & n70003;
  assign n70005 = P2_P2_INSTQUEUE_REG_2__0_ & n70004;
  assign n70006 = ~P2_P2_INSTQUEUERD_ADDR_REG_0_ & n68228;
  assign n70007 = n69996 & n70006;
  assign n70008 = P2_P2_INSTQUEUE_REG_3__0_ & n70007;
  assign n70009 = ~n69999 & ~n70002;
  assign n70010 = ~n70005 & n70009;
  assign n70011 = ~n70008 & n70010;
  assign n70012 = ~n68116 & n69870;
  assign n70013 = n69997 & n70012;
  assign n70014 = P2_P2_INSTQUEUE_REG_4__0_ & n70013;
  assign n70015 = n70000 & n70012;
  assign n70016 = P2_P2_INSTQUEUE_REG_5__0_ & n70015;
  assign n70017 = n70003 & n70012;
  assign n70018 = P2_P2_INSTQUEUE_REG_6__0_ & n70017;
  assign n70019 = n70006 & n70012;
  assign n70020 = P2_P2_INSTQUEUE_REG_7__0_ & n70019;
  assign n70021 = ~n70014 & ~n70016;
  assign n70022 = ~n70018 & n70021;
  assign n70023 = ~n70020 & n70022;
  assign n70024 = n68116 & ~n69870;
  assign n70025 = n69997 & n70024;
  assign n70026 = P2_P2_INSTQUEUE_REG_8__0_ & n70025;
  assign n70027 = n70000 & n70024;
  assign n70028 = P2_P2_INSTQUEUE_REG_9__0_ & n70027;
  assign n70029 = n70003 & n70024;
  assign n70030 = P2_P2_INSTQUEUE_REG_10__0_ & n70029;
  assign n70031 = n70006 & n70024;
  assign n70032 = P2_P2_INSTQUEUE_REG_11__0_ & n70031;
  assign n70033 = ~n70026 & ~n70028;
  assign n70034 = ~n70030 & n70033;
  assign n70035 = ~n70032 & n70034;
  assign n70036 = ~n68116 & ~n69870;
  assign n70037 = n69997 & n70036;
  assign n70038 = P2_P2_INSTQUEUE_REG_12__0_ & n70037;
  assign n70039 = n70000 & n70036;
  assign n70040 = P2_P2_INSTQUEUE_REG_13__0_ & n70039;
  assign n70041 = n70003 & n70036;
  assign n70042 = P2_P2_INSTQUEUE_REG_14__0_ & n70041;
  assign n70043 = n70006 & n70036;
  assign n70044 = P2_P2_INSTQUEUE_REG_15__0_ & n70043;
  assign n70045 = ~n70038 & ~n70040;
  assign n70046 = ~n70042 & n70045;
  assign n70047 = ~n70044 & n70046;
  assign n70048 = n70011 & n70023;
  assign n70049 = n70035 & n70048;
  assign n70050 = n70047 & n70049;
  assign n70051 = P2_P2_INSTADDRPOINTER_REG_0_ & n70050;
  assign n70052 = ~P2_P2_INSTADDRPOINTER_REG_0_ & ~n70050;
  assign n70053 = ~n70051 & ~n70052;
  assign n70054 = P2_P2_INSTQUEUE_REG_0__7_ & n69998;
  assign n70055 = P2_P2_INSTQUEUE_REG_1__7_ & n70001;
  assign n70056 = P2_P2_INSTQUEUE_REG_2__7_ & n70004;
  assign n70057 = P2_P2_INSTQUEUE_REG_3__7_ & n70007;
  assign n70058 = ~n70054 & ~n70055;
  assign n70059 = ~n70056 & n70058;
  assign n70060 = ~n70057 & n70059;
  assign n70061 = P2_P2_INSTQUEUE_REG_4__7_ & n70013;
  assign n70062 = P2_P2_INSTQUEUE_REG_5__7_ & n70015;
  assign n70063 = P2_P2_INSTQUEUE_REG_6__7_ & n70017;
  assign n70064 = P2_P2_INSTQUEUE_REG_7__7_ & n70019;
  assign n70065 = ~n70061 & ~n70062;
  assign n70066 = ~n70063 & n70065;
  assign n70067 = ~n70064 & n70066;
  assign n70068 = P2_P2_INSTQUEUE_REG_8__7_ & n70025;
  assign n70069 = P2_P2_INSTQUEUE_REG_9__7_ & n70027;
  assign n70070 = P2_P2_INSTQUEUE_REG_10__7_ & n70029;
  assign n70071 = P2_P2_INSTQUEUE_REG_11__7_ & n70031;
  assign n70072 = ~n70068 & ~n70069;
  assign n70073 = ~n70070 & n70072;
  assign n70074 = ~n70071 & n70073;
  assign n70075 = P2_P2_INSTQUEUE_REG_12__7_ & n70037;
  assign n70076 = P2_P2_INSTQUEUE_REG_13__7_ & n70039;
  assign n70077 = P2_P2_INSTQUEUE_REG_14__7_ & n70041;
  assign n70078 = P2_P2_INSTQUEUE_REG_15__7_ & n70043;
  assign n70079 = ~n70075 & ~n70076;
  assign n70080 = ~n70077 & n70079;
  assign n70081 = ~n70078 & n70080;
  assign n70082 = n70060 & n70067;
  assign n70083 = n70074 & n70082;
  assign n70084 = n70081 & n70083;
  assign n70085 = n68021 & ~n70084;
  assign n70086 = ~n70053 & n70085;
  assign n70087 = n68021 & n70084;
  assign n70088 = ~n70053 & n70087;
  assign n70089 = ~n69985 & ~n69986;
  assign n70090 = n69995 & n70089;
  assign n70091 = ~n70086 & n70090;
  assign n70092 = ~n70088 & n70091;
  assign n70093 = n67987 & n68015;
  assign n70094 = ~P2_P2_INSTADDRPOINTER_REG_0_ & n70093;
  assign n70095 = ~P2_P2_INSTADDRPOINTER_REG_0_ & n68059;
  assign n70096 = n67816 & n68002;
  assign n70097 = n68048 & n70096;
  assign n70098 = ~P2_P2_INSTADDRPOINTER_REG_0_ & n70097;
  assign n70099 = ~P2_P2_INSTADDRPOINTER_REG_0_ & n70050;
  assign n70100 = P2_P2_INSTADDRPOINTER_REG_0_ & ~n70050;
  assign n70101 = ~n70099 & ~n70100;
  assign n70102 = n68016 & ~n70101;
  assign n70103 = n67691 & n68045;
  assign n70104 = n68048 & n70103;
  assign n70105 = ~P2_P2_INSTADDRPOINTER_REG_0_ & n70104;
  assign n70106 = ~n70094 & ~n70095;
  assign n70107 = ~n70098 & n70106;
  assign n70108 = ~n70102 & n70107;
  assign n70109 = ~n70105 & n70108;
  assign n70110 = P2_P2_INSTADDRPOINTER_REG_0_ & n67915;
  assign n70111 = P2_P2_INSTADDRPOINTER_REG_0_ & n67993;
  assign n70112 = P2_P2_INSTADDRPOINTER_REG_0_ & n67997;
  assign n70113 = ~P2_P2_INSTADDRPOINTER_REG_0_ & n68013;
  assign n70114 = ~P2_P2_INSTADDRPOINTER_REG_0_ & n68005;
  assign n70115 = ~n70110 & ~n70111;
  assign n70116 = ~n70112 & n70115;
  assign n70117 = ~n70113 & n70116;
  assign n70118 = ~n70114 & n70117;
  assign n70119 = n70109 & n70118;
  assign n70120 = n69983 & ~n69984;
  assign n70121 = n70092 & n70120;
  assign n70122 = n70119 & n70121;
  assign n70123 = n69980 & ~n70122;
  assign n70124 = ~P2_P2_STATE2_REG_2_ & ~n69979;
  assign n70125 = P2_P2_REIP_REG_0_ & n70124;
  assign n70126 = P2_P2_INSTADDRPOINTER_REG_0_ & n69979;
  assign n70127 = ~n70123 & ~n70125;
  assign n13286 = n70126 | ~n70127;
  assign n70129 = P2_P2_INSTADDRPOINTER_REG_1_ & n69979;
  assign n70130 = P2_P2_REIP_REG_1_ & n70124;
  assign n70131 = ~n68102 & ~n68296;
  assign n70132 = n68212 & ~n68296;
  assign n70133 = n68055 & ~n68296;
  assign n70134 = ~n70132 & ~n70133;
  assign n70135 = ~P2_P2_INSTADDRPOINTER_REG_1_ & n70100;
  assign n70136 = P2_P2_INSTADDRPOINTER_REG_1_ & ~n70100;
  assign n70137 = ~n70135 & ~n70136;
  assign n70138 = P2_P2_INSTQUEUE_REG_0__1_ & n69998;
  assign n70139 = P2_P2_INSTQUEUE_REG_1__1_ & n70001;
  assign n70140 = P2_P2_INSTQUEUE_REG_2__1_ & n70004;
  assign n70141 = P2_P2_INSTQUEUE_REG_3__1_ & n70007;
  assign n70142 = ~n70138 & ~n70139;
  assign n70143 = ~n70140 & n70142;
  assign n70144 = ~n70141 & n70143;
  assign n70145 = P2_P2_INSTQUEUE_REG_4__1_ & n70013;
  assign n70146 = P2_P2_INSTQUEUE_REG_5__1_ & n70015;
  assign n70147 = P2_P2_INSTQUEUE_REG_6__1_ & n70017;
  assign n70148 = P2_P2_INSTQUEUE_REG_7__1_ & n70019;
  assign n70149 = ~n70145 & ~n70146;
  assign n70150 = ~n70147 & n70149;
  assign n70151 = ~n70148 & n70150;
  assign n70152 = P2_P2_INSTQUEUE_REG_8__1_ & n70025;
  assign n70153 = P2_P2_INSTQUEUE_REG_9__1_ & n70027;
  assign n70154 = P2_P2_INSTQUEUE_REG_10__1_ & n70029;
  assign n70155 = P2_P2_INSTQUEUE_REG_11__1_ & n70031;
  assign n70156 = ~n70152 & ~n70153;
  assign n70157 = ~n70154 & n70156;
  assign n70158 = ~n70155 & n70157;
  assign n70159 = P2_P2_INSTQUEUE_REG_12__1_ & n70037;
  assign n70160 = P2_P2_INSTQUEUE_REG_13__1_ & n70039;
  assign n70161 = P2_P2_INSTQUEUE_REG_14__1_ & n70041;
  assign n70162 = P2_P2_INSTQUEUE_REG_15__1_ & n70043;
  assign n70163 = ~n70159 & ~n70160;
  assign n70164 = ~n70161 & n70163;
  assign n70165 = ~n70162 & n70164;
  assign n70166 = n70144 & n70151;
  assign n70167 = n70158 & n70166;
  assign n70168 = n70165 & n70167;
  assign n70169 = ~n70137 & ~n70168;
  assign n70170 = ~P2_P2_INSTADDRPOINTER_REG_1_ & ~n70100;
  assign n70171 = n70168 & n70170;
  assign n70172 = n70100 & n70168;
  assign n70173 = P2_P2_INSTADDRPOINTER_REG_1_ & n70172;
  assign n70174 = ~n70169 & ~n70171;
  assign n70175 = ~n70173 & n70174;
  assign n70176 = n70087 & ~n70175;
  assign n70177 = ~n68296 & n70104;
  assign n70178 = ~n68296 & n70097;
  assign n70179 = ~n68296 & n70093;
  assign n70180 = n68059 & ~n68296;
  assign n70181 = ~n70177 & ~n70178;
  assign n70182 = ~n70179 & n70181;
  assign n70183 = ~n70180 & n70182;
  assign n70184 = ~P2_P2_INSTADDRPOINTER_REG_1_ & n67915;
  assign n70185 = ~P2_P2_INSTADDRPOINTER_REG_1_ & n67993;
  assign n70186 = ~P2_P2_INSTADDRPOINTER_REG_1_ & n67997;
  assign n70187 = n68013 & ~n68296;
  assign n70188 = n68005 & ~n68296;
  assign n70189 = ~n70184 & ~n70185;
  assign n70190 = ~n70186 & n70189;
  assign n70191 = ~n70187 & n70190;
  assign n70192 = ~n70188 & n70191;
  assign n70193 = ~P2_P2_INSTADDRPOINTER_REG_1_ & n70051;
  assign n70194 = P2_P2_INSTADDRPOINTER_REG_1_ & ~n70051;
  assign n70195 = ~n70193 & ~n70194;
  assign n70196 = ~n70050 & n70168;
  assign n70197 = n70050 & ~n70168;
  assign n70198 = ~n70196 & ~n70197;
  assign n70199 = ~n70195 & n70198;
  assign n70200 = ~P2_P2_INSTADDRPOINTER_REG_1_ & ~n70051;
  assign n70201 = ~n70198 & n70200;
  assign n70202 = n70051 & ~n70198;
  assign n70203 = P2_P2_INSTADDRPOINTER_REG_1_ & n70202;
  assign n70204 = ~n70199 & ~n70201;
  assign n70205 = ~n70203 & n70204;
  assign n70206 = n68016 & ~n70205;
  assign n70207 = n70183 & n70192;
  assign n70208 = ~n70206 & n70207;
  assign n70209 = ~P2_P2_INSTADDRPOINTER_REG_1_ & n68173;
  assign n70210 = ~P2_P2_INSTADDRPOINTER_REG_1_ & n68174;
  assign n70211 = ~n68296 & n69988;
  assign n70212 = ~n68296 & n69991;
  assign n70213 = ~n70211 & ~n70212;
  assign n70214 = ~P2_P2_INSTADDRPOINTER_REG_1_ & n67989;
  assign n70215 = n70213 & ~n70214;
  assign n70216 = n70100 & ~n70168;
  assign n70217 = ~n70100 & n70168;
  assign n70218 = ~n70216 & ~n70217;
  assign n70219 = ~P2_P2_INSTADDRPOINTER_REG_1_ & ~n70218;
  assign n70220 = ~n70100 & ~n70168;
  assign n70221 = P2_P2_INSTADDRPOINTER_REG_1_ & n70220;
  assign n70222 = P2_P2_INSTADDRPOINTER_REG_1_ & n70100;
  assign n70223 = n70168 & n70222;
  assign n70224 = ~n70219 & ~n70221;
  assign n70225 = ~n70223 & n70224;
  assign n70226 = n70085 & ~n70225;
  assign n70227 = ~n70209 & ~n70210;
  assign n70228 = n70215 & n70227;
  assign n70229 = ~n70226 & n70228;
  assign n70230 = ~n70131 & n70134;
  assign n70231 = ~n70176 & n70230;
  assign n70232 = n70208 & n70231;
  assign n70233 = n70229 & n70232;
  assign n70234 = n69980 & ~n70233;
  assign n70235 = ~n70129 & ~n70130;
  assign n13291 = n70234 | ~n70235;
  assign n70237 = P2_P2_INSTADDRPOINTER_REG_2_ & n69979;
  assign n70238 = P2_P2_REIP_REG_2_ & n70124;
  assign n70239 = P2_P2_INSTADDRPOINTER_REG_0_ & P2_P2_INSTADDRPOINTER_REG_1_;
  assign n70240 = ~P2_P2_INSTADDRPOINTER_REG_2_ & n70239;
  assign n70241 = P2_P2_INSTADDRPOINTER_REG_2_ & ~n70239;
  assign n70242 = ~n70240 & ~n70241;
  assign n70243 = ~n68102 & ~n70242;
  assign n70244 = P2_P2_INSTADDRPOINTER_REG_1_ & ~P2_P2_INSTADDRPOINTER_REG_2_;
  assign n70245 = ~P2_P2_INSTADDRPOINTER_REG_1_ & P2_P2_INSTADDRPOINTER_REG_2_;
  assign n70246 = ~n70244 & ~n70245;
  assign n70247 = n68173 & ~n70246;
  assign n70248 = n68174 & ~n70246;
  assign n70249 = n69988 & ~n70242;
  assign n70250 = n69991 & ~n70242;
  assign n70251 = ~n70249 & ~n70250;
  assign n70252 = n67989 & ~n70246;
  assign n70253 = n70251 & ~n70252;
  assign n70254 = ~n70247 & ~n70248;
  assign n70255 = n70253 & n70254;
  assign n70256 = P2_P2_INSTADDRPOINTER_REG_1_ & ~n70220;
  assign n70257 = ~n70172 & ~n70256;
  assign n70258 = P2_P2_INSTQUEUE_REG_0__2_ & n69998;
  assign n70259 = P2_P2_INSTQUEUE_REG_1__2_ & n70001;
  assign n70260 = P2_P2_INSTQUEUE_REG_2__2_ & n70004;
  assign n70261 = P2_P2_INSTQUEUE_REG_3__2_ & n70007;
  assign n70262 = ~n70258 & ~n70259;
  assign n70263 = ~n70260 & n70262;
  assign n70264 = ~n70261 & n70263;
  assign n70265 = P2_P2_INSTQUEUE_REG_4__2_ & n70013;
  assign n70266 = P2_P2_INSTQUEUE_REG_5__2_ & n70015;
  assign n70267 = P2_P2_INSTQUEUE_REG_6__2_ & n70017;
  assign n70268 = P2_P2_INSTQUEUE_REG_7__2_ & n70019;
  assign n70269 = ~n70265 & ~n70266;
  assign n70270 = ~n70267 & n70269;
  assign n70271 = ~n70268 & n70270;
  assign n70272 = P2_P2_INSTQUEUE_REG_8__2_ & n70025;
  assign n70273 = P2_P2_INSTQUEUE_REG_9__2_ & n70027;
  assign n70274 = P2_P2_INSTQUEUE_REG_10__2_ & n70029;
  assign n70275 = P2_P2_INSTQUEUE_REG_11__2_ & n70031;
  assign n70276 = ~n70272 & ~n70273;
  assign n70277 = ~n70274 & n70276;
  assign n70278 = ~n70275 & n70277;
  assign n70279 = P2_P2_INSTQUEUE_REG_12__2_ & n70037;
  assign n70280 = P2_P2_INSTQUEUE_REG_13__2_ & n70039;
  assign n70281 = P2_P2_INSTQUEUE_REG_14__2_ & n70041;
  assign n70282 = P2_P2_INSTQUEUE_REG_15__2_ & n70043;
  assign n70283 = ~n70279 & ~n70280;
  assign n70284 = ~n70281 & n70283;
  assign n70285 = ~n70282 & n70284;
  assign n70286 = n70264 & n70271;
  assign n70287 = n70278 & n70286;
  assign n70288 = n70285 & n70287;
  assign n70289 = ~n70168 & n70288;
  assign n70290 = n70168 & ~n70288;
  assign n70291 = ~n70289 & ~n70290;
  assign n70292 = ~P2_P2_INSTADDRPOINTER_REG_2_ & ~n70291;
  assign n70293 = P2_P2_INSTADDRPOINTER_REG_2_ & n70291;
  assign n70294 = ~n70292 & ~n70293;
  assign n70295 = n70257 & ~n70294;
  assign n70296 = ~n70257 & n70294;
  assign n70297 = ~n70295 & ~n70296;
  assign n70298 = n70087 & ~n70297;
  assign n70299 = n68212 & ~n70242;
  assign n70300 = n68055 & ~n70242;
  assign n70301 = ~n70299 & ~n70300;
  assign n70302 = P2_P2_INSTADDRPOINTER_REG_1_ & n70168;
  assign n70303 = ~n70172 & ~n70222;
  assign n70304 = ~n70302 & n70303;
  assign n70305 = ~n70294 & n70304;
  assign n70306 = ~P2_P2_INSTADDRPOINTER_REG_2_ & n70291;
  assign n70307 = P2_P2_INSTADDRPOINTER_REG_2_ & ~n70291;
  assign n70308 = ~n70306 & ~n70307;
  assign n70309 = ~n70304 & ~n70308;
  assign n70310 = ~n70305 & ~n70309;
  assign n70311 = n70085 & ~n70310;
  assign n70312 = n70301 & ~n70311;
  assign n70313 = n70104 & ~n70242;
  assign n70314 = n70097 & ~n70242;
  assign n70315 = n70093 & ~n70242;
  assign n70316 = n68059 & ~n70242;
  assign n70317 = ~n70313 & ~n70314;
  assign n70318 = ~n70315 & n70317;
  assign n70319 = ~n70316 & n70318;
  assign n70320 = n67915 & ~n70246;
  assign n70321 = n67993 & ~n70246;
  assign n70322 = n67997 & ~n70246;
  assign n70323 = ~P2_P2_INSTADDRPOINTER_REG_2_ & ~n70239;
  assign n70324 = P2_P2_INSTADDRPOINTER_REG_2_ & n70239;
  assign n70325 = ~n70323 & ~n70324;
  assign n70326 = n68013 & ~n70325;
  assign n70327 = n68005 & ~n70325;
  assign n70328 = ~n70320 & ~n70321;
  assign n70329 = ~n70322 & n70328;
  assign n70330 = ~n70326 & n70329;
  assign n70331 = ~n70327 & n70330;
  assign n70332 = ~n70050 & ~n70168;
  assign n70333 = n70288 & ~n70332;
  assign n70334 = ~n70288 & n70332;
  assign n70335 = ~n70333 & ~n70334;
  assign n70336 = ~P2_P2_INSTADDRPOINTER_REG_2_ & ~n70335;
  assign n70337 = P2_P2_INSTADDRPOINTER_REG_2_ & n70335;
  assign n70338 = ~n70336 & ~n70337;
  assign n70339 = ~n70051 & n70198;
  assign n70340 = P2_P2_INSTADDRPOINTER_REG_1_ & ~n70339;
  assign n70341 = ~n70202 & ~n70340;
  assign n70342 = ~n70338 & n70341;
  assign n70343 = ~P2_P2_INSTADDRPOINTER_REG_2_ & n70335;
  assign n70344 = P2_P2_INSTADDRPOINTER_REG_2_ & ~n70335;
  assign n70345 = ~n70343 & ~n70344;
  assign n70346 = ~n70341 & ~n70345;
  assign n70347 = ~n70342 & ~n70346;
  assign n70348 = n68016 & ~n70347;
  assign n70349 = n70319 & n70331;
  assign n70350 = ~n70348 & n70349;
  assign n70351 = ~n70243 & n70255;
  assign n70352 = ~n70298 & n70351;
  assign n70353 = n70312 & n70352;
  assign n70354 = n70350 & n70353;
  assign n70355 = n69980 & ~n70354;
  assign n70356 = ~n70237 & ~n70238;
  assign n13296 = n70355 | ~n70356;
  assign n70358 = P2_P2_INSTADDRPOINTER_REG_3_ & n69979;
  assign n70359 = P2_P2_REIP_REG_3_ & n70124;
  assign n70360 = ~P2_P2_INSTADDRPOINTER_REG_3_ & n70324;
  assign n70361 = P2_P2_INSTADDRPOINTER_REG_3_ & ~n70324;
  assign n70362 = ~n70360 & ~n70361;
  assign n70363 = n68212 & ~n70362;
  assign n70364 = n68055 & ~n70362;
  assign n70365 = ~n70363 & ~n70364;
  assign n70366 = ~n68102 & ~n70362;
  assign n70367 = P2_P2_INSTADDRPOINTER_REG_1_ & P2_P2_INSTADDRPOINTER_REG_2_;
  assign n70368 = ~P2_P2_INSTADDRPOINTER_REG_3_ & n70367;
  assign n70369 = P2_P2_INSTADDRPOINTER_REG_3_ & ~n70367;
  assign n70370 = ~n70368 & ~n70369;
  assign n70371 = n68173 & ~n70370;
  assign n70372 = n68174 & ~n70370;
  assign n70373 = n69988 & ~n70362;
  assign n70374 = n69991 & ~n70362;
  assign n70375 = ~n70373 & ~n70374;
  assign n70376 = n67989 & ~n70370;
  assign n70377 = n70375 & ~n70376;
  assign n70378 = ~n70371 & ~n70372;
  assign n70379 = n70377 & n70378;
  assign n70380 = ~n70304 & ~n70306;
  assign n70381 = ~n70307 & ~n70380;
  assign n70382 = P2_P2_INSTQUEUE_REG_0__3_ & n69998;
  assign n70383 = P2_P2_INSTQUEUE_REG_1__3_ & n70001;
  assign n70384 = P2_P2_INSTQUEUE_REG_2__3_ & n70004;
  assign n70385 = P2_P2_INSTQUEUE_REG_3__3_ & n70007;
  assign n70386 = ~n70382 & ~n70383;
  assign n70387 = ~n70384 & n70386;
  assign n70388 = ~n70385 & n70387;
  assign n70389 = P2_P2_INSTQUEUE_REG_4__3_ & n70013;
  assign n70390 = P2_P2_INSTQUEUE_REG_5__3_ & n70015;
  assign n70391 = P2_P2_INSTQUEUE_REG_6__3_ & n70017;
  assign n70392 = P2_P2_INSTQUEUE_REG_7__3_ & n70019;
  assign n70393 = ~n70389 & ~n70390;
  assign n70394 = ~n70391 & n70393;
  assign n70395 = ~n70392 & n70394;
  assign n70396 = P2_P2_INSTQUEUE_REG_8__3_ & n70025;
  assign n70397 = P2_P2_INSTQUEUE_REG_9__3_ & n70027;
  assign n70398 = P2_P2_INSTQUEUE_REG_10__3_ & n70029;
  assign n70399 = P2_P2_INSTQUEUE_REG_11__3_ & n70031;
  assign n70400 = ~n70396 & ~n70397;
  assign n70401 = ~n70398 & n70400;
  assign n70402 = ~n70399 & n70401;
  assign n70403 = P2_P2_INSTQUEUE_REG_12__3_ & n70037;
  assign n70404 = P2_P2_INSTQUEUE_REG_13__3_ & n70039;
  assign n70405 = P2_P2_INSTQUEUE_REG_14__3_ & n70041;
  assign n70406 = P2_P2_INSTQUEUE_REG_15__3_ & n70043;
  assign n70407 = ~n70403 & ~n70404;
  assign n70408 = ~n70405 & n70407;
  assign n70409 = ~n70406 & n70408;
  assign n70410 = n70388 & n70395;
  assign n70411 = n70402 & n70410;
  assign n70412 = n70409 & n70411;
  assign n70413 = ~n70168 & ~n70288;
  assign n70414 = n70412 & ~n70413;
  assign n70415 = ~n70412 & n70413;
  assign n70416 = ~n70414 & ~n70415;
  assign n70417 = P2_P2_INSTADDRPOINTER_REG_3_ & ~n70416;
  assign n70418 = ~P2_P2_INSTADDRPOINTER_REG_3_ & n70416;
  assign n70419 = ~n70417 & ~n70418;
  assign n70420 = n70381 & ~n70419;
  assign n70421 = P2_P2_INSTADDRPOINTER_REG_3_ & n70416;
  assign n70422 = ~P2_P2_INSTADDRPOINTER_REG_3_ & ~n70416;
  assign n70423 = ~n70421 & ~n70422;
  assign n70424 = ~n70381 & ~n70423;
  assign n70425 = ~n70420 & ~n70424;
  assign n70426 = n70085 & ~n70425;
  assign n70427 = ~n70257 & ~n70306;
  assign n70428 = ~n70307 & ~n70427;
  assign n70429 = n70412 & n70413;
  assign n70430 = ~n70412 & ~n70413;
  assign n70431 = ~n70429 & ~n70430;
  assign n70432 = ~P2_P2_INSTADDRPOINTER_REG_3_ & n70431;
  assign n70433 = ~n70428 & ~n70432;
  assign n70434 = P2_P2_INSTADDRPOINTER_REG_3_ & ~n70431;
  assign n70435 = n70433 & ~n70434;
  assign n70436 = ~P2_P2_INSTADDRPOINTER_REG_3_ & ~n70431;
  assign n70437 = P2_P2_INSTADDRPOINTER_REG_3_ & n70431;
  assign n70438 = ~n70436 & ~n70437;
  assign n70439 = n70428 & n70438;
  assign n70440 = ~n70435 & ~n70439;
  assign n70441 = n70087 & n70440;
  assign n70442 = ~n70426 & ~n70441;
  assign n70443 = n70104 & ~n70362;
  assign n70444 = n70097 & ~n70362;
  assign n70445 = n70093 & ~n70362;
  assign n70446 = n68059 & ~n70362;
  assign n70447 = ~n70443 & ~n70444;
  assign n70448 = ~n70445 & n70447;
  assign n70449 = ~n70446 & n70448;
  assign n70450 = n67915 & ~n70370;
  assign n70451 = n67993 & ~n70370;
  assign n70452 = n67997 & ~n70370;
  assign n70453 = ~P2_P2_INSTADDRPOINTER_REG_3_ & n70323;
  assign n70454 = P2_P2_INSTADDRPOINTER_REG_3_ & ~n70323;
  assign n70455 = ~n70453 & ~n70454;
  assign n70456 = n68013 & n70455;
  assign n70457 = n68005 & n70455;
  assign n70458 = ~n70450 & ~n70451;
  assign n70459 = ~n70452 & n70458;
  assign n70460 = ~n70456 & n70459;
  assign n70461 = ~n70457 & n70460;
  assign n70462 = n70341 & ~n70344;
  assign n70463 = n70333 & n70412;
  assign n70464 = ~n70333 & ~n70412;
  assign n70465 = ~n70463 & ~n70464;
  assign n70466 = P2_P2_INSTADDRPOINTER_REG_3_ & n70465;
  assign n70467 = ~n70343 & n70465;
  assign n70468 = P2_P2_INSTADDRPOINTER_REG_3_ & ~n70343;
  assign n70469 = ~n70467 & ~n70468;
  assign n70470 = ~n70462 & ~n70466;
  assign n70471 = ~n70469 & n70470;
  assign n70472 = ~P2_P2_INSTADDRPOINTER_REG_3_ & n70465;
  assign n70473 = P2_P2_INSTADDRPOINTER_REG_3_ & ~n70465;
  assign n70474 = ~n70472 & ~n70473;
  assign n70475 = ~n70344 & n70474;
  assign n70476 = ~n70341 & ~n70343;
  assign n70477 = n70475 & ~n70476;
  assign n70478 = ~n70471 & ~n70477;
  assign n70479 = n68016 & n70478;
  assign n70480 = n70449 & n70461;
  assign n70481 = ~n70479 & n70480;
  assign n70482 = n70365 & ~n70366;
  assign n70483 = n70379 & n70482;
  assign n70484 = n70442 & n70483;
  assign n70485 = n70481 & n70484;
  assign n70486 = n69980 & ~n70485;
  assign n70487 = ~n70358 & ~n70359;
  assign n13301 = n70486 | ~n70487;
  assign n70489 = P2_P2_INSTADDRPOINTER_REG_4_ & n69979;
  assign n70490 = P2_P2_REIP_REG_4_ & n70124;
  assign n70491 = P2_P2_INSTADDRPOINTER_REG_3_ & n70324;
  assign n70492 = ~P2_P2_INSTADDRPOINTER_REG_4_ & n70491;
  assign n70493 = P2_P2_INSTADDRPOINTER_REG_4_ & ~n70491;
  assign n70494 = ~n70492 & ~n70493;
  assign n70495 = ~n68102 & ~n70494;
  assign n70496 = P2_P2_INSTADDRPOINTER_REG_3_ & n70367;
  assign n70497 = ~P2_P2_INSTADDRPOINTER_REG_4_ & n70496;
  assign n70498 = P2_P2_INSTADDRPOINTER_REG_4_ & ~n70496;
  assign n70499 = ~n70497 & ~n70498;
  assign n70500 = n68173 & ~n70499;
  assign n70501 = n68174 & ~n70499;
  assign n70502 = n69988 & ~n70494;
  assign n70503 = n69991 & ~n70494;
  assign n70504 = ~n70502 & ~n70503;
  assign n70505 = n67989 & ~n70499;
  assign n70506 = n70504 & ~n70505;
  assign n70507 = ~n70500 & ~n70501;
  assign n70508 = n70506 & n70507;
  assign n70509 = P2_P2_INSTQUEUE_REG_0__4_ & n69998;
  assign n70510 = P2_P2_INSTQUEUE_REG_1__4_ & n70001;
  assign n70511 = P2_P2_INSTQUEUE_REG_2__4_ & n70004;
  assign n70512 = P2_P2_INSTQUEUE_REG_3__4_ & n70007;
  assign n70513 = ~n70509 & ~n70510;
  assign n70514 = ~n70511 & n70513;
  assign n70515 = ~n70512 & n70514;
  assign n70516 = P2_P2_INSTQUEUE_REG_4__4_ & n70013;
  assign n70517 = P2_P2_INSTQUEUE_REG_5__4_ & n70015;
  assign n70518 = P2_P2_INSTQUEUE_REG_6__4_ & n70017;
  assign n70519 = P2_P2_INSTQUEUE_REG_7__4_ & n70019;
  assign n70520 = ~n70516 & ~n70517;
  assign n70521 = ~n70518 & n70520;
  assign n70522 = ~n70519 & n70521;
  assign n70523 = P2_P2_INSTQUEUE_REG_8__4_ & n70025;
  assign n70524 = P2_P2_INSTQUEUE_REG_9__4_ & n70027;
  assign n70525 = P2_P2_INSTQUEUE_REG_10__4_ & n70029;
  assign n70526 = P2_P2_INSTQUEUE_REG_11__4_ & n70031;
  assign n70527 = ~n70523 & ~n70524;
  assign n70528 = ~n70525 & n70527;
  assign n70529 = ~n70526 & n70528;
  assign n70530 = P2_P2_INSTQUEUE_REG_12__4_ & n70037;
  assign n70531 = P2_P2_INSTQUEUE_REG_13__4_ & n70039;
  assign n70532 = P2_P2_INSTQUEUE_REG_14__4_ & n70041;
  assign n70533 = P2_P2_INSTQUEUE_REG_15__4_ & n70043;
  assign n70534 = ~n70530 & ~n70531;
  assign n70535 = ~n70532 & n70534;
  assign n70536 = ~n70533 & n70535;
  assign n70537 = n70515 & n70522;
  assign n70538 = n70529 & n70537;
  assign n70539 = n70536 & n70538;
  assign n70540 = n70415 & n70539;
  assign n70541 = ~n70415 & ~n70539;
  assign n70542 = ~n70540 & ~n70541;
  assign n70543 = P2_P2_INSTADDRPOINTER_REG_4_ & ~n70542;
  assign n70544 = ~P2_P2_INSTADDRPOINTER_REG_4_ & n70542;
  assign n70545 = ~n70543 & ~n70544;
  assign n70546 = ~n70433 & ~n70434;
  assign n70547 = n70545 & ~n70546;
  assign n70548 = ~P2_P2_INSTADDRPOINTER_REG_4_ & ~n70542;
  assign n70549 = P2_P2_INSTADDRPOINTER_REG_4_ & n70542;
  assign n70550 = ~n70548 & ~n70549;
  assign n70551 = ~n70434 & n70550;
  assign n70552 = ~n70433 & n70551;
  assign n70553 = ~n70547 & ~n70552;
  assign n70554 = n70087 & n70553;
  assign n70555 = n68212 & ~n70494;
  assign n70556 = n68055 & ~n70494;
  assign n70557 = ~n70555 & ~n70556;
  assign n70558 = ~n70306 & ~n70422;
  assign n70559 = ~n70172 & ~n70302;
  assign n70560 = ~n70307 & n70559;
  assign n70561 = ~n70222 & n70560;
  assign n70562 = n70558 & ~n70561;
  assign n70563 = ~n70421 & ~n70562;
  assign n70564 = n70415 & ~n70539;
  assign n70565 = ~n70415 & n70539;
  assign n70566 = ~n70564 & ~n70565;
  assign n70567 = P2_P2_INSTADDRPOINTER_REG_4_ & ~n70566;
  assign n70568 = ~P2_P2_INSTADDRPOINTER_REG_4_ & n70566;
  assign n70569 = ~n70567 & ~n70568;
  assign n70570 = n70563 & ~n70569;
  assign n70571 = P2_P2_INSTADDRPOINTER_REG_4_ & n70566;
  assign n70572 = ~P2_P2_INSTADDRPOINTER_REG_4_ & ~n70566;
  assign n70573 = ~n70571 & ~n70572;
  assign n70574 = ~n70563 & ~n70573;
  assign n70575 = ~n70570 & ~n70574;
  assign n70576 = n70085 & ~n70575;
  assign n70577 = n70557 & ~n70576;
  assign n70578 = n70104 & ~n70494;
  assign n70579 = n70097 & ~n70494;
  assign n70580 = n70093 & ~n70494;
  assign n70581 = n68059 & ~n70494;
  assign n70582 = ~n70578 & ~n70579;
  assign n70583 = ~n70580 & n70582;
  assign n70584 = ~n70581 & n70583;
  assign n70585 = n67915 & ~n70499;
  assign n70586 = n67993 & ~n70499;
  assign n70587 = n67997 & ~n70499;
  assign n70588 = ~P2_P2_INSTADDRPOINTER_REG_4_ & n70454;
  assign n70589 = P2_P2_INSTADDRPOINTER_REG_4_ & ~n70454;
  assign n70590 = ~n70588 & ~n70589;
  assign n70591 = n68013 & ~n70590;
  assign n70592 = n68005 & ~n70590;
  assign n70593 = ~n70585 & ~n70586;
  assign n70594 = ~n70587 & n70593;
  assign n70595 = ~n70591 & n70594;
  assign n70596 = ~n70592 & n70595;
  assign n70597 = n70464 & n70539;
  assign n70598 = ~n70464 & ~n70539;
  assign n70599 = ~n70597 & ~n70598;
  assign n70600 = ~P2_P2_INSTADDRPOINTER_REG_4_ & ~n70599;
  assign n70601 = P2_P2_INSTADDRPOINTER_REG_4_ & n70599;
  assign n70602 = ~n70600 & ~n70601;
  assign n70603 = n70344 & n70465;
  assign n70604 = ~n70344 & ~n70465;
  assign n70605 = P2_P2_INSTADDRPOINTER_REG_3_ & ~n70604;
  assign n70606 = ~n70603 & ~n70605;
  assign n70607 = ~n70341 & ~n70469;
  assign n70608 = n70606 & ~n70607;
  assign n70609 = ~n70602 & n70608;
  assign n70610 = ~P2_P2_INSTADDRPOINTER_REG_4_ & n70599;
  assign n70611 = P2_P2_INSTADDRPOINTER_REG_4_ & ~n70599;
  assign n70612 = ~n70610 & ~n70611;
  assign n70613 = ~n70608 & ~n70612;
  assign n70614 = ~n70609 & ~n70613;
  assign n70615 = n68016 & ~n70614;
  assign n70616 = n70584 & n70596;
  assign n70617 = ~n70615 & n70616;
  assign n70618 = ~n70495 & n70508;
  assign n70619 = ~n70554 & n70618;
  assign n70620 = n70577 & n70619;
  assign n70621 = n70617 & n70620;
  assign n70622 = n69980 & ~n70621;
  assign n70623 = ~n70489 & ~n70490;
  assign n13306 = n70622 | ~n70623;
  assign n70625 = P2_P2_INSTADDRPOINTER_REG_5_ & n69979;
  assign n70626 = P2_P2_REIP_REG_5_ & n70124;
  assign n70627 = P2_P2_INSTADDRPOINTER_REG_4_ & n70496;
  assign n70628 = ~P2_P2_INSTADDRPOINTER_REG_5_ & n70627;
  assign n70629 = P2_P2_INSTADDRPOINTER_REG_5_ & ~n70627;
  assign n70630 = ~n70628 & ~n70629;
  assign n70631 = n68173 & ~n70630;
  assign n70632 = n68174 & ~n70630;
  assign n70633 = P2_P2_INSTADDRPOINTER_REG_4_ & n70491;
  assign n70634 = ~P2_P2_INSTADDRPOINTER_REG_5_ & n70633;
  assign n70635 = P2_P2_INSTADDRPOINTER_REG_5_ & ~n70633;
  assign n70636 = ~n70634 & ~n70635;
  assign n70637 = n69988 & ~n70636;
  assign n70638 = n69991 & ~n70636;
  assign n70639 = ~n70637 & ~n70638;
  assign n70640 = n67989 & ~n70630;
  assign n70641 = n70639 & ~n70640;
  assign n70642 = ~n70631 & ~n70632;
  assign n70643 = n70641 & n70642;
  assign n70644 = ~n68102 & ~n70636;
  assign n70645 = n70421 & ~n70572;
  assign n70646 = ~n70571 & ~n70645;
  assign n70647 = n70558 & ~n70572;
  assign n70648 = ~n70561 & n70647;
  assign n70649 = n70646 & ~n70648;
  assign n70650 = P2_P2_INSTQUEUE_REG_0__5_ & n69998;
  assign n70651 = P2_P2_INSTQUEUE_REG_1__5_ & n70001;
  assign n70652 = P2_P2_INSTQUEUE_REG_2__5_ & n70004;
  assign n70653 = P2_P2_INSTQUEUE_REG_3__5_ & n70007;
  assign n70654 = ~n70650 & ~n70651;
  assign n70655 = ~n70652 & n70654;
  assign n70656 = ~n70653 & n70655;
  assign n70657 = P2_P2_INSTQUEUE_REG_4__5_ & n70013;
  assign n70658 = P2_P2_INSTQUEUE_REG_5__5_ & n70015;
  assign n70659 = P2_P2_INSTQUEUE_REG_6__5_ & n70017;
  assign n70660 = P2_P2_INSTQUEUE_REG_7__5_ & n70019;
  assign n70661 = ~n70657 & ~n70658;
  assign n70662 = ~n70659 & n70661;
  assign n70663 = ~n70660 & n70662;
  assign n70664 = P2_P2_INSTQUEUE_REG_8__5_ & n70025;
  assign n70665 = P2_P2_INSTQUEUE_REG_9__5_ & n70027;
  assign n70666 = P2_P2_INSTQUEUE_REG_10__5_ & n70029;
  assign n70667 = P2_P2_INSTQUEUE_REG_11__5_ & n70031;
  assign n70668 = ~n70664 & ~n70665;
  assign n70669 = ~n70666 & n70668;
  assign n70670 = ~n70667 & n70669;
  assign n70671 = P2_P2_INSTQUEUE_REG_12__5_ & n70037;
  assign n70672 = P2_P2_INSTQUEUE_REG_13__5_ & n70039;
  assign n70673 = P2_P2_INSTQUEUE_REG_14__5_ & n70041;
  assign n70674 = P2_P2_INSTQUEUE_REG_15__5_ & n70043;
  assign n70675 = ~n70671 & ~n70672;
  assign n70676 = ~n70673 & n70675;
  assign n70677 = ~n70674 & n70676;
  assign n70678 = n70656 & n70663;
  assign n70679 = n70670 & n70678;
  assign n70680 = n70677 & n70679;
  assign n70681 = ~n70564 & n70680;
  assign n70682 = ~n70539 & ~n70680;
  assign n70683 = n70415 & n70682;
  assign n70684 = ~n70681 & ~n70683;
  assign n70685 = P2_P2_INSTADDRPOINTER_REG_5_ & ~n70684;
  assign n70686 = ~P2_P2_INSTADDRPOINTER_REG_5_ & n70684;
  assign n70687 = ~n70685 & ~n70686;
  assign n70688 = n70649 & ~n70687;
  assign n70689 = ~n70649 & n70687;
  assign n70690 = ~n70688 & ~n70689;
  assign n70691 = n70085 & ~n70690;
  assign n70692 = n68212 & ~n70636;
  assign n70693 = n68055 & ~n70636;
  assign n70694 = ~n70692 & ~n70693;
  assign n70695 = n70434 & ~n70544;
  assign n70696 = ~n70543 & ~n70695;
  assign n70697 = ~n70432 & ~n70544;
  assign n70698 = ~n70428 & n70697;
  assign n70699 = n70696 & ~n70698;
  assign n70700 = n70564 & n70680;
  assign n70701 = ~n70564 & ~n70680;
  assign n70702 = ~n70700 & ~n70701;
  assign n70703 = ~P2_P2_INSTADDRPOINTER_REG_5_ & ~n70702;
  assign n70704 = P2_P2_INSTADDRPOINTER_REG_5_ & n70702;
  assign n70705 = ~n70703 & ~n70704;
  assign n70706 = n70699 & ~n70705;
  assign n70707 = ~n70699 & n70705;
  assign n70708 = ~n70706 & ~n70707;
  assign n70709 = n70087 & ~n70708;
  assign n70710 = n70694 & ~n70709;
  assign n70711 = n70104 & ~n70636;
  assign n70712 = n70097 & ~n70636;
  assign n70713 = n70093 & ~n70636;
  assign n70714 = n68059 & ~n70636;
  assign n70715 = ~n70711 & ~n70712;
  assign n70716 = ~n70713 & n70715;
  assign n70717 = ~n70714 & n70716;
  assign n70718 = n67915 & ~n70630;
  assign n70719 = n67993 & ~n70630;
  assign n70720 = n67997 & ~n70630;
  assign n70721 = P2_P2_INSTADDRPOINTER_REG_4_ & n70454;
  assign n70722 = ~P2_P2_INSTADDRPOINTER_REG_5_ & n70721;
  assign n70723 = P2_P2_INSTADDRPOINTER_REG_5_ & ~n70721;
  assign n70724 = ~n70722 & ~n70723;
  assign n70725 = n68013 & ~n70724;
  assign n70726 = n68005 & ~n70724;
  assign n70727 = ~n70718 & ~n70719;
  assign n70728 = ~n70720 & n70727;
  assign n70729 = ~n70725 & n70728;
  assign n70730 = ~n70726 & n70729;
  assign n70731 = n70464 & ~n70539;
  assign n70732 = n70680 & n70731;
  assign n70733 = ~n70680 & ~n70731;
  assign n70734 = ~n70732 & ~n70733;
  assign n70735 = P2_P2_INSTADDRPOINTER_REG_5_ & ~n70734;
  assign n70736 = ~P2_P2_INSTADDRPOINTER_REG_5_ & n70734;
  assign n70737 = ~n70610 & ~n70736;
  assign n70738 = ~n70735 & n70737;
  assign n70739 = n70608 & ~n70611;
  assign n70740 = n70738 & ~n70739;
  assign n70741 = ~P2_P2_INSTADDRPOINTER_REG_5_ & ~n70734;
  assign n70742 = P2_P2_INSTADDRPOINTER_REG_5_ & n70734;
  assign n70743 = ~n70741 & ~n70742;
  assign n70744 = ~n70611 & n70743;
  assign n70745 = ~n70608 & ~n70610;
  assign n70746 = n70744 & ~n70745;
  assign n70747 = ~n70740 & ~n70746;
  assign n70748 = n68016 & n70747;
  assign n70749 = n70717 & n70730;
  assign n70750 = ~n70748 & n70749;
  assign n70751 = n70643 & ~n70644;
  assign n70752 = ~n70691 & n70751;
  assign n70753 = n70710 & n70752;
  assign n70754 = n70750 & n70753;
  assign n70755 = n69980 & ~n70754;
  assign n70756 = ~n70625 & ~n70626;
  assign n13311 = n70755 | ~n70756;
  assign n70758 = P2_P2_INSTADDRPOINTER_REG_6_ & n69979;
  assign n70759 = P2_P2_REIP_REG_6_ & n70124;
  assign n70760 = P2_P2_INSTADDRPOINTER_REG_5_ & n70627;
  assign n70761 = ~P2_P2_INSTADDRPOINTER_REG_6_ & n70760;
  assign n70762 = P2_P2_INSTADDRPOINTER_REG_6_ & ~n70760;
  assign n70763 = ~n70761 & ~n70762;
  assign n70764 = n68173 & ~n70763;
  assign n70765 = n68174 & ~n70763;
  assign n70766 = P2_P2_INSTADDRPOINTER_REG_5_ & n70633;
  assign n70767 = ~P2_P2_INSTADDRPOINTER_REG_6_ & n70766;
  assign n70768 = P2_P2_INSTADDRPOINTER_REG_6_ & ~n70766;
  assign n70769 = ~n70767 & ~n70768;
  assign n70770 = n69988 & ~n70769;
  assign n70771 = n69991 & ~n70769;
  assign n70772 = ~n70770 & ~n70771;
  assign n70773 = n67989 & ~n70763;
  assign n70774 = n70772 & ~n70773;
  assign n70775 = ~n70764 & ~n70765;
  assign n70776 = n70774 & n70775;
  assign n70777 = ~n68102 & ~n70769;
  assign n70778 = ~P2_P2_INSTADDRPOINTER_REG_5_ & ~n70684;
  assign n70779 = ~n70649 & ~n70778;
  assign n70780 = P2_P2_INSTADDRPOINTER_REG_5_ & n70684;
  assign n70781 = ~n70779 & ~n70780;
  assign n70782 = P2_P2_INSTQUEUE_REG_0__6_ & n69998;
  assign n70783 = P2_P2_INSTQUEUE_REG_1__6_ & n70001;
  assign n70784 = P2_P2_INSTQUEUE_REG_2__6_ & n70004;
  assign n70785 = P2_P2_INSTQUEUE_REG_3__6_ & n70007;
  assign n70786 = ~n70782 & ~n70783;
  assign n70787 = ~n70784 & n70786;
  assign n70788 = ~n70785 & n70787;
  assign n70789 = P2_P2_INSTQUEUE_REG_4__6_ & n70013;
  assign n70790 = P2_P2_INSTQUEUE_REG_5__6_ & n70015;
  assign n70791 = P2_P2_INSTQUEUE_REG_6__6_ & n70017;
  assign n70792 = P2_P2_INSTQUEUE_REG_7__6_ & n70019;
  assign n70793 = ~n70789 & ~n70790;
  assign n70794 = ~n70791 & n70793;
  assign n70795 = ~n70792 & n70794;
  assign n70796 = P2_P2_INSTQUEUE_REG_8__6_ & n70025;
  assign n70797 = P2_P2_INSTQUEUE_REG_9__6_ & n70027;
  assign n70798 = P2_P2_INSTQUEUE_REG_10__6_ & n70029;
  assign n70799 = P2_P2_INSTQUEUE_REG_11__6_ & n70031;
  assign n70800 = ~n70796 & ~n70797;
  assign n70801 = ~n70798 & n70800;
  assign n70802 = ~n70799 & n70801;
  assign n70803 = P2_P2_INSTQUEUE_REG_12__6_ & n70037;
  assign n70804 = P2_P2_INSTQUEUE_REG_13__6_ & n70039;
  assign n70805 = P2_P2_INSTQUEUE_REG_14__6_ & n70041;
  assign n70806 = P2_P2_INSTQUEUE_REG_15__6_ & n70043;
  assign n70807 = ~n70803 & ~n70804;
  assign n70808 = ~n70805 & n70807;
  assign n70809 = ~n70806 & n70808;
  assign n70810 = n70788 & n70795;
  assign n70811 = n70802 & n70810;
  assign n70812 = n70809 & n70811;
  assign n70813 = n70683 & ~n70812;
  assign n70814 = ~n70683 & n70812;
  assign n70815 = ~n70813 & ~n70814;
  assign n70816 = P2_P2_INSTADDRPOINTER_REG_6_ & ~n70815;
  assign n70817 = ~P2_P2_INSTADDRPOINTER_REG_6_ & n70815;
  assign n70818 = ~n70816 & ~n70817;
  assign n70819 = n70781 & ~n70818;
  assign n70820 = ~n70781 & n70818;
  assign n70821 = ~n70819 & ~n70820;
  assign n70822 = n70085 & ~n70821;
  assign n70823 = n68212 & ~n70769;
  assign n70824 = n68055 & ~n70769;
  assign n70825 = ~n70823 & ~n70824;
  assign n70826 = ~n70699 & ~n70702;
  assign n70827 = P2_P2_INSTADDRPOINTER_REG_5_ & ~n70699;
  assign n70828 = P2_P2_INSTADDRPOINTER_REG_5_ & ~n70702;
  assign n70829 = ~n70826 & ~n70827;
  assign n70830 = ~n70828 & n70829;
  assign n70831 = n70564 & ~n70680;
  assign n70832 = n70812 & n70831;
  assign n70833 = ~n70812 & ~n70831;
  assign n70834 = ~n70832 & ~n70833;
  assign n70835 = ~P2_P2_INSTADDRPOINTER_REG_6_ & ~n70834;
  assign n70836 = P2_P2_INSTADDRPOINTER_REG_6_ & n70834;
  assign n70837 = ~n70835 & ~n70836;
  assign n70838 = n70830 & ~n70837;
  assign n70839 = ~n70830 & n70837;
  assign n70840 = ~n70838 & ~n70839;
  assign n70841 = n70087 & ~n70840;
  assign n70842 = n70825 & ~n70841;
  assign n70843 = n70104 & ~n70769;
  assign n70844 = n70097 & ~n70769;
  assign n70845 = n70093 & ~n70769;
  assign n70846 = n68059 & ~n70769;
  assign n70847 = ~n70843 & ~n70844;
  assign n70848 = ~n70845 & n70847;
  assign n70849 = ~n70846 & n70848;
  assign n70850 = n67915 & ~n70763;
  assign n70851 = n67993 & ~n70763;
  assign n70852 = n67997 & ~n70763;
  assign n70853 = P2_P2_INSTADDRPOINTER_REG_5_ & n70721;
  assign n70854 = ~P2_P2_INSTADDRPOINTER_REG_6_ & n70853;
  assign n70855 = P2_P2_INSTADDRPOINTER_REG_6_ & ~n70853;
  assign n70856 = ~n70854 & ~n70855;
  assign n70857 = n68013 & ~n70856;
  assign n70858 = n68005 & ~n70856;
  assign n70859 = ~n70850 & ~n70851;
  assign n70860 = ~n70852 & n70859;
  assign n70861 = ~n70857 & n70860;
  assign n70862 = ~n70858 & n70861;
  assign n70863 = n70611 & ~n70734;
  assign n70864 = ~n70611 & n70734;
  assign n70865 = P2_P2_INSTADDRPOINTER_REG_5_ & ~n70864;
  assign n70866 = ~n70863 & ~n70865;
  assign n70867 = ~n70608 & n70737;
  assign n70868 = n70866 & ~n70867;
  assign n70869 = ~n70680 & n70731;
  assign n70870 = n70812 & n70869;
  assign n70871 = ~n70812 & ~n70869;
  assign n70872 = ~n70870 & ~n70871;
  assign n70873 = ~P2_P2_INSTADDRPOINTER_REG_6_ & ~n70872;
  assign n70874 = P2_P2_INSTADDRPOINTER_REG_6_ & n70872;
  assign n70875 = ~n70873 & ~n70874;
  assign n70876 = n70868 & ~n70875;
  assign n70877 = ~n70868 & n70875;
  assign n70878 = ~n70876 & ~n70877;
  assign n70879 = n68016 & ~n70878;
  assign n70880 = n70849 & n70862;
  assign n70881 = ~n70879 & n70880;
  assign n70882 = n70776 & ~n70777;
  assign n70883 = ~n70822 & n70882;
  assign n70884 = n70842 & n70883;
  assign n70885 = n70881 & n70884;
  assign n70886 = n69980 & ~n70885;
  assign n70887 = ~n70758 & ~n70759;
  assign n13316 = n70886 | ~n70887;
  assign n70889 = P2_P2_INSTADDRPOINTER_REG_7_ & n69979;
  assign n70890 = P2_P2_REIP_REG_7_ & n70124;
  assign n70891 = P2_P2_INSTADDRPOINTER_REG_6_ & n70760;
  assign n70892 = ~P2_P2_INSTADDRPOINTER_REG_7_ & n70891;
  assign n70893 = P2_P2_INSTADDRPOINTER_REG_7_ & ~n70891;
  assign n70894 = ~n70892 & ~n70893;
  assign n70895 = n68173 & ~n70894;
  assign n70896 = n68174 & ~n70894;
  assign n70897 = P2_P2_INSTADDRPOINTER_REG_6_ & n70766;
  assign n70898 = ~P2_P2_INSTADDRPOINTER_REG_7_ & n70897;
  assign n70899 = P2_P2_INSTADDRPOINTER_REG_7_ & ~n70897;
  assign n70900 = ~n70898 & ~n70899;
  assign n70901 = n69988 & ~n70900;
  assign n70902 = n69991 & ~n70900;
  assign n70903 = ~n70901 & ~n70902;
  assign n70904 = n67989 & ~n70894;
  assign n70905 = n70903 & ~n70904;
  assign n70906 = ~n70895 & ~n70896;
  assign n70907 = n70905 & n70906;
  assign n70908 = ~n68102 & ~n70900;
  assign n70909 = P2_P2_INSTADDRPOINTER_REG_6_ & n70815;
  assign n70910 = ~P2_P2_INSTADDRPOINTER_REG_6_ & ~n70815;
  assign n70911 = ~n70781 & ~n70910;
  assign n70912 = ~n70909 & ~n70911;
  assign n70913 = n70084 & ~n70813;
  assign n70914 = ~n70084 & ~n70812;
  assign n70915 = n70683 & n70914;
  assign n70916 = ~n70913 & ~n70915;
  assign n70917 = P2_P2_INSTADDRPOINTER_REG_7_ & ~n70916;
  assign n70918 = ~P2_P2_INSTADDRPOINTER_REG_7_ & n70916;
  assign n70919 = ~n70917 & ~n70918;
  assign n70920 = n70912 & ~n70919;
  assign n70921 = ~n70912 & n70919;
  assign n70922 = ~n70920 & ~n70921;
  assign n70923 = n70085 & ~n70922;
  assign n70924 = n68212 & ~n70900;
  assign n70925 = n68055 & ~n70900;
  assign n70926 = ~n70924 & ~n70925;
  assign n70927 = P2_P2_INSTADDRPOINTER_REG_6_ & ~n70834;
  assign n70928 = ~P2_P2_INSTADDRPOINTER_REG_6_ & n70834;
  assign n70929 = ~n70830 & ~n70928;
  assign n70930 = ~n70927 & ~n70929;
  assign n70931 = ~n70812 & n70831;
  assign n70932 = n70084 & n70931;
  assign n70933 = ~n70084 & ~n70931;
  assign n70934 = ~n70932 & ~n70933;
  assign n70935 = ~P2_P2_INSTADDRPOINTER_REG_7_ & ~n70934;
  assign n70936 = P2_P2_INSTADDRPOINTER_REG_7_ & n70934;
  assign n70937 = ~n70935 & ~n70936;
  assign n70938 = n70930 & ~n70937;
  assign n70939 = ~n70930 & n70937;
  assign n70940 = ~n70938 & ~n70939;
  assign n70941 = n70087 & ~n70940;
  assign n70942 = n70926 & ~n70941;
  assign n70943 = n70104 & ~n70900;
  assign n70944 = n70097 & ~n70900;
  assign n70945 = n70093 & ~n70900;
  assign n70946 = n68059 & ~n70900;
  assign n70947 = ~n70943 & ~n70944;
  assign n70948 = ~n70945 & n70947;
  assign n70949 = ~n70946 & n70948;
  assign n70950 = n67915 & ~n70894;
  assign n70951 = n67993 & ~n70894;
  assign n70952 = n67997 & ~n70894;
  assign n70953 = P2_P2_INSTADDRPOINTER_REG_6_ & n70853;
  assign n70954 = ~P2_P2_INSTADDRPOINTER_REG_7_ & n70953;
  assign n70955 = P2_P2_INSTADDRPOINTER_REG_7_ & ~n70953;
  assign n70956 = ~n70954 & ~n70955;
  assign n70957 = n68013 & ~n70956;
  assign n70958 = n68005 & ~n70956;
  assign n70959 = ~n70950 & ~n70951;
  assign n70960 = ~n70952 & n70959;
  assign n70961 = ~n70957 & n70960;
  assign n70962 = ~n70958 & n70961;
  assign n70963 = P2_P2_INSTADDRPOINTER_REG_6_ & ~n70872;
  assign n70964 = ~P2_P2_INSTADDRPOINTER_REG_6_ & n70872;
  assign n70965 = ~n70868 & ~n70964;
  assign n70966 = ~n70963 & ~n70965;
  assign n70967 = ~n70812 & n70869;
  assign n70968 = n70084 & n70967;
  assign n70969 = ~n70084 & ~n70967;
  assign n70970 = ~n70968 & ~n70969;
  assign n70971 = ~P2_P2_INSTADDRPOINTER_REG_7_ & ~n70970;
  assign n70972 = P2_P2_INSTADDRPOINTER_REG_7_ & n70970;
  assign n70973 = ~n70971 & ~n70972;
  assign n70974 = n70966 & ~n70973;
  assign n70975 = ~n70966 & n70973;
  assign n70976 = ~n70974 & ~n70975;
  assign n70977 = n68016 & ~n70976;
  assign n70978 = n70949 & n70962;
  assign n70979 = ~n70977 & n70978;
  assign n70980 = n70907 & ~n70908;
  assign n70981 = ~n70923 & n70980;
  assign n70982 = n70942 & n70981;
  assign n70983 = n70979 & n70982;
  assign n70984 = n69980 & ~n70983;
  assign n70985 = ~n70889 & ~n70890;
  assign n13321 = n70984 | ~n70985;
  assign n70987 = P2_P2_INSTADDRPOINTER_REG_8_ & n69979;
  assign n70988 = P2_P2_REIP_REG_8_ & n70124;
  assign n70989 = P2_P2_INSTADDRPOINTER_REG_7_ & n70891;
  assign n70990 = ~P2_P2_INSTADDRPOINTER_REG_8_ & n70989;
  assign n70991 = P2_P2_INSTADDRPOINTER_REG_8_ & ~n70989;
  assign n70992 = ~n70990 & ~n70991;
  assign n70993 = n68173 & ~n70992;
  assign n70994 = n68174 & ~n70992;
  assign n70995 = n67989 & ~n70992;
  assign n70996 = P2_P2_INSTADDRPOINTER_REG_7_ & n70897;
  assign n70997 = ~P2_P2_INSTADDRPOINTER_REG_8_ & n70996;
  assign n70998 = P2_P2_INSTADDRPOINTER_REG_8_ & ~n70996;
  assign n70999 = ~n70997 & ~n70998;
  assign n71000 = n69991 & ~n70999;
  assign n71001 = n69988 & ~n70999;
  assign n71002 = ~n70995 & ~n71000;
  assign n71003 = ~n71001 & n71002;
  assign n71004 = ~n70993 & ~n70994;
  assign n71005 = n71003 & n71004;
  assign n71006 = ~n68102 & ~n70999;
  assign n71007 = ~P2_P2_INSTADDRPOINTER_REG_7_ & ~n70916;
  assign n71008 = ~n70912 & ~n71007;
  assign n71009 = P2_P2_INSTADDRPOINTER_REG_7_ & n70916;
  assign n71010 = ~n71008 & ~n71009;
  assign n71011 = ~P2_P2_INSTADDRPOINTER_REG_8_ & ~n70915;
  assign n71012 = P2_P2_INSTADDRPOINTER_REG_8_ & n70915;
  assign n71013 = ~n71011 & ~n71012;
  assign n71014 = n71010 & ~n71013;
  assign n71015 = ~n71010 & n71013;
  assign n71016 = ~n71014 & ~n71015;
  assign n71017 = n70085 & ~n71016;
  assign n71018 = n68212 & ~n70999;
  assign n71019 = n68055 & ~n70999;
  assign n71020 = ~n71018 & ~n71019;
  assign n71021 = ~n70930 & ~n70934;
  assign n71022 = P2_P2_INSTADDRPOINTER_REG_7_ & ~n70930;
  assign n71023 = P2_P2_INSTADDRPOINTER_REG_7_ & ~n70934;
  assign n71024 = ~n71021 & ~n71022;
  assign n71025 = ~n71023 & n71024;
  assign n71026 = n70831 & n70914;
  assign n71027 = ~P2_P2_INSTADDRPOINTER_REG_8_ & n71026;
  assign n71028 = P2_P2_INSTADDRPOINTER_REG_8_ & ~n71026;
  assign n71029 = ~n71027 & ~n71028;
  assign n71030 = n71025 & ~n71029;
  assign n71031 = ~n71025 & n71029;
  assign n71032 = ~n71030 & ~n71031;
  assign n71033 = n70087 & ~n71032;
  assign n71034 = n71020 & ~n71033;
  assign n71035 = n70104 & ~n70999;
  assign n71036 = n68059 & ~n70999;
  assign n71037 = n70093 & ~n70999;
  assign n71038 = n70097 & ~n70999;
  assign n71039 = ~n71035 & ~n71036;
  assign n71040 = ~n71037 & n71039;
  assign n71041 = ~n71038 & n71040;
  assign n71042 = n67915 & ~n70992;
  assign n71043 = n67993 & ~n70992;
  assign n71044 = n67997 & ~n70992;
  assign n71045 = P2_P2_INSTADDRPOINTER_REG_7_ & n70953;
  assign n71046 = ~P2_P2_INSTADDRPOINTER_REG_8_ & n71045;
  assign n71047 = P2_P2_INSTADDRPOINTER_REG_8_ & ~n71045;
  assign n71048 = ~n71046 & ~n71047;
  assign n71049 = n68013 & ~n71048;
  assign n71050 = n68005 & ~n71048;
  assign n71051 = ~n71042 & ~n71043;
  assign n71052 = ~n71044 & n71051;
  assign n71053 = ~n71049 & n71052;
  assign n71054 = ~n71050 & n71053;
  assign n71055 = ~n70966 & ~n70970;
  assign n71056 = P2_P2_INSTADDRPOINTER_REG_7_ & ~n70966;
  assign n71057 = P2_P2_INSTADDRPOINTER_REG_7_ & ~n70970;
  assign n71058 = ~n71055 & ~n71056;
  assign n71059 = ~n71057 & n71058;
  assign n71060 = n70869 & n70914;
  assign n71061 = ~P2_P2_INSTADDRPOINTER_REG_8_ & n71060;
  assign n71062 = P2_P2_INSTADDRPOINTER_REG_8_ & ~n71060;
  assign n71063 = ~n71061 & ~n71062;
  assign n71064 = n71059 & ~n71063;
  assign n71065 = ~n71059 & n71063;
  assign n71066 = ~n71064 & ~n71065;
  assign n71067 = n68016 & ~n71066;
  assign n71068 = n71041 & n71054;
  assign n71069 = ~n71067 & n71068;
  assign n71070 = n71005 & ~n71006;
  assign n71071 = ~n71017 & n71070;
  assign n71072 = n71034 & n71071;
  assign n71073 = n71069 & n71072;
  assign n71074 = n69980 & ~n71073;
  assign n71075 = ~n70987 & ~n70988;
  assign n13326 = n71074 | ~n71075;
  assign n71077 = P2_P2_INSTADDRPOINTER_REG_9_ & n69979;
  assign n71078 = P2_P2_REIP_REG_9_ & n70124;
  assign n71079 = P2_P2_INSTADDRPOINTER_REG_8_ & n70989;
  assign n71080 = ~P2_P2_INSTADDRPOINTER_REG_9_ & n71079;
  assign n71081 = P2_P2_INSTADDRPOINTER_REG_9_ & ~n71079;
  assign n71082 = ~n71080 & ~n71081;
  assign n71083 = n68173 & ~n71082;
  assign n71084 = n68174 & ~n71082;
  assign n71085 = P2_P2_INSTADDRPOINTER_REG_8_ & n70996;
  assign n71086 = ~P2_P2_INSTADDRPOINTER_REG_9_ & n71085;
  assign n71087 = P2_P2_INSTADDRPOINTER_REG_9_ & ~n71085;
  assign n71088 = ~n71086 & ~n71087;
  assign n71089 = n69988 & ~n71088;
  assign n71090 = n67989 & ~n71082;
  assign n71091 = n69991 & ~n71088;
  assign n71092 = ~n71090 & ~n71091;
  assign n71093 = ~n71083 & ~n71084;
  assign n71094 = ~n71089 & n71093;
  assign n71095 = n71092 & n71094;
  assign n71096 = ~n68102 & ~n71088;
  assign n71097 = ~P2_P2_INSTADDRPOINTER_REG_8_ & n70915;
  assign n71098 = ~n71010 & ~n71097;
  assign n71099 = P2_P2_INSTADDRPOINTER_REG_8_ & ~n70915;
  assign n71100 = ~n71098 & ~n71099;
  assign n71101 = P2_P2_INSTADDRPOINTER_REG_9_ & n70915;
  assign n71102 = ~P2_P2_INSTADDRPOINTER_REG_9_ & ~n70915;
  assign n71103 = ~n71101 & ~n71102;
  assign n71104 = n71100 & ~n71103;
  assign n71105 = P2_P2_INSTADDRPOINTER_REG_9_ & ~n70915;
  assign n71106 = ~P2_P2_INSTADDRPOINTER_REG_9_ & n70915;
  assign n71107 = ~n71105 & ~n71106;
  assign n71108 = ~n71100 & ~n71107;
  assign n71109 = ~n71104 & ~n71108;
  assign n71110 = n70085 & ~n71109;
  assign n71111 = n68212 & ~n71088;
  assign n71112 = n68055 & ~n71088;
  assign n71113 = ~n71111 & ~n71112;
  assign n71114 = P2_P2_INSTADDRPOINTER_REG_8_ & n71026;
  assign n71115 = ~P2_P2_INSTADDRPOINTER_REG_8_ & ~n71026;
  assign n71116 = ~n71025 & ~n71115;
  assign n71117 = ~n71114 & ~n71116;
  assign n71118 = ~P2_P2_INSTADDRPOINTER_REG_9_ & n71117;
  assign n71119 = P2_P2_INSTADDRPOINTER_REG_9_ & ~n71117;
  assign n71120 = ~n71118 & ~n71119;
  assign n71121 = n70087 & n71120;
  assign n71122 = n71113 & ~n71121;
  assign n71123 = n70104 & ~n71088;
  assign n71124 = n68059 & ~n71088;
  assign n71125 = n70093 & ~n71088;
  assign n71126 = n70097 & ~n71088;
  assign n71127 = ~n71123 & ~n71124;
  assign n71128 = ~n71125 & n71127;
  assign n71129 = ~n71126 & n71128;
  assign n71130 = n67915 & ~n71082;
  assign n71131 = n67993 & ~n71082;
  assign n71132 = n67997 & ~n71082;
  assign n71133 = P2_P2_INSTADDRPOINTER_REG_8_ & n71045;
  assign n71134 = ~P2_P2_INSTADDRPOINTER_REG_9_ & n71133;
  assign n71135 = P2_P2_INSTADDRPOINTER_REG_9_ & ~n71133;
  assign n71136 = ~n71134 & ~n71135;
  assign n71137 = n68013 & ~n71136;
  assign n71138 = n68005 & ~n71136;
  assign n71139 = ~n71130 & ~n71131;
  assign n71140 = ~n71132 & n71139;
  assign n71141 = ~n71137 & n71140;
  assign n71142 = ~n71138 & n71141;
  assign n71143 = P2_P2_INSTADDRPOINTER_REG_8_ & n71060;
  assign n71144 = ~P2_P2_INSTADDRPOINTER_REG_8_ & ~n71060;
  assign n71145 = ~n71059 & ~n71144;
  assign n71146 = ~n71143 & ~n71145;
  assign n71147 = ~P2_P2_INSTADDRPOINTER_REG_9_ & n71146;
  assign n71148 = P2_P2_INSTADDRPOINTER_REG_9_ & ~n71146;
  assign n71149 = ~n71147 & ~n71148;
  assign n71150 = n68016 & n71149;
  assign n71151 = n71129 & n71142;
  assign n71152 = ~n71150 & n71151;
  assign n71153 = n71095 & ~n71096;
  assign n71154 = ~n71110 & n71153;
  assign n71155 = n71122 & n71154;
  assign n71156 = n71152 & n71155;
  assign n71157 = n69980 & ~n71156;
  assign n71158 = ~n71077 & ~n71078;
  assign n13331 = n71157 | ~n71158;
  assign n71160 = P2_P2_INSTADDRPOINTER_REG_10_ & n69979;
  assign n71161 = P2_P2_REIP_REG_10_ & n70124;
  assign n71162 = P2_P2_INSTADDRPOINTER_REG_9_ & n71079;
  assign n71163 = ~P2_P2_INSTADDRPOINTER_REG_10_ & n71162;
  assign n71164 = P2_P2_INSTADDRPOINTER_REG_10_ & ~n71162;
  assign n71165 = ~n71163 & ~n71164;
  assign n71166 = n68173 & ~n71165;
  assign n71167 = n68174 & ~n71165;
  assign n71168 = P2_P2_INSTADDRPOINTER_REG_9_ & n71085;
  assign n71169 = ~P2_P2_INSTADDRPOINTER_REG_10_ & n71168;
  assign n71170 = P2_P2_INSTADDRPOINTER_REG_10_ & ~n71168;
  assign n71171 = ~n71169 & ~n71170;
  assign n71172 = n69988 & ~n71171;
  assign n71173 = n67989 & ~n71165;
  assign n71174 = n69991 & ~n71171;
  assign n71175 = ~n71173 & ~n71174;
  assign n71176 = ~n71166 & ~n71167;
  assign n71177 = ~n71172 & n71176;
  assign n71178 = n71175 & n71177;
  assign n71179 = ~n68102 & ~n71171;
  assign n71180 = ~n71097 & ~n71106;
  assign n71181 = ~n71010 & n71180;
  assign n71182 = ~n71099 & ~n71105;
  assign n71183 = ~n71181 & n71182;
  assign n71184 = ~P2_P2_INSTADDRPOINTER_REG_10_ & ~n70915;
  assign n71185 = P2_P2_INSTADDRPOINTER_REG_10_ & n70915;
  assign n71186 = ~n71184 & ~n71185;
  assign n71187 = n71183 & ~n71186;
  assign n71188 = P2_P2_INSTADDRPOINTER_REG_10_ & ~n70915;
  assign n71189 = ~P2_P2_INSTADDRPOINTER_REG_10_ & n70915;
  assign n71190 = ~n71188 & ~n71189;
  assign n71191 = ~n71183 & ~n71190;
  assign n71192 = ~n71187 & ~n71191;
  assign n71193 = n70085 & ~n71192;
  assign n71194 = n68212 & ~n71171;
  assign n71195 = n68055 & ~n71171;
  assign n71196 = ~n71194 & ~n71195;
  assign n71197 = ~P2_P2_INSTADDRPOINTER_REG_10_ & ~n71119;
  assign n71198 = P2_P2_INSTADDRPOINTER_REG_9_ & P2_P2_INSTADDRPOINTER_REG_10_;
  assign n71199 = ~n71117 & n71198;
  assign n71200 = ~n71197 & ~n71199;
  assign n71201 = n70087 & n71200;
  assign n71202 = n71196 & ~n71201;
  assign n71203 = n70104 & ~n71171;
  assign n71204 = n68059 & ~n71171;
  assign n71205 = n70093 & ~n71171;
  assign n71206 = n70097 & ~n71171;
  assign n71207 = ~n71203 & ~n71204;
  assign n71208 = ~n71205 & n71207;
  assign n71209 = ~n71206 & n71208;
  assign n71210 = n67915 & ~n71165;
  assign n71211 = n67993 & ~n71165;
  assign n71212 = n67997 & ~n71165;
  assign n71213 = P2_P2_INSTADDRPOINTER_REG_9_ & n71133;
  assign n71214 = ~P2_P2_INSTADDRPOINTER_REG_10_ & n71213;
  assign n71215 = P2_P2_INSTADDRPOINTER_REG_10_ & ~n71213;
  assign n71216 = ~n71214 & ~n71215;
  assign n71217 = n68013 & ~n71216;
  assign n71218 = n68005 & ~n71216;
  assign n71219 = ~n71210 & ~n71211;
  assign n71220 = ~n71212 & n71219;
  assign n71221 = ~n71217 & n71220;
  assign n71222 = ~n71218 & n71221;
  assign n71223 = ~P2_P2_INSTADDRPOINTER_REG_10_ & ~n71148;
  assign n71224 = ~n71146 & n71198;
  assign n71225 = ~n71223 & ~n71224;
  assign n71226 = n68016 & n71225;
  assign n71227 = n71209 & n71222;
  assign n71228 = ~n71226 & n71227;
  assign n71229 = n71178 & ~n71179;
  assign n71230 = ~n71193 & n71229;
  assign n71231 = n71202 & n71230;
  assign n71232 = n71228 & n71231;
  assign n71233 = n69980 & ~n71232;
  assign n71234 = ~n71160 & ~n71161;
  assign n13336 = n71233 | ~n71234;
  assign n71236 = P2_P2_INSTADDRPOINTER_REG_11_ & n69979;
  assign n71237 = P2_P2_REIP_REG_11_ & n70124;
  assign n71238 = ~n71236 & ~n71237;
  assign n71239 = P2_P2_INSTADDRPOINTER_REG_10_ & n71168;
  assign n71240 = ~P2_P2_INSTADDRPOINTER_REG_11_ & n71239;
  assign n71241 = P2_P2_INSTADDRPOINTER_REG_11_ & ~n71239;
  assign n71242 = ~n71240 & ~n71241;
  assign n71243 = n70104 & ~n71242;
  assign n71244 = n68059 & ~n71242;
  assign n71245 = n70093 & ~n71242;
  assign n71246 = n70097 & ~n71242;
  assign n71247 = ~n71243 & ~n71244;
  assign n71248 = ~n71245 & n71247;
  assign n71249 = ~n71246 & n71248;
  assign n71250 = P2_P2_INSTADDRPOINTER_REG_10_ & n71162;
  assign n71251 = ~P2_P2_INSTADDRPOINTER_REG_11_ & n71250;
  assign n71252 = P2_P2_INSTADDRPOINTER_REG_11_ & ~n71250;
  assign n71253 = ~n71251 & ~n71252;
  assign n71254 = n67915 & ~n71253;
  assign n71255 = n67993 & ~n71253;
  assign n71256 = n67997 & ~n71253;
  assign n71257 = P2_P2_INSTADDRPOINTER_REG_10_ & n71213;
  assign n71258 = ~P2_P2_INSTADDRPOINTER_REG_11_ & n71257;
  assign n71259 = P2_P2_INSTADDRPOINTER_REG_11_ & ~n71257;
  assign n71260 = ~n71258 & ~n71259;
  assign n71261 = n68013 & ~n71260;
  assign n71262 = n68005 & ~n71260;
  assign n71263 = ~n71254 & ~n71255;
  assign n71264 = ~n71256 & n71263;
  assign n71265 = ~n71261 & n71264;
  assign n71266 = ~n71262 & n71265;
  assign n71267 = P2_P2_INSTADDRPOINTER_REG_11_ & ~n71224;
  assign n71268 = ~P2_P2_INSTADDRPOINTER_REG_11_ & n71224;
  assign n71269 = ~n71267 & ~n71268;
  assign n71270 = n68016 & ~n71269;
  assign n71271 = n71249 & n71266;
  assign n71272 = ~n71270 & n71271;
  assign n71273 = n68212 & ~n71242;
  assign n71274 = n68055 & ~n71242;
  assign n71275 = ~n71273 & ~n71274;
  assign n71276 = ~n68102 & ~n71242;
  assign n71277 = n71182 & ~n71188;
  assign n71278 = n71180 & ~n71189;
  assign n71279 = ~n71010 & n71278;
  assign n71280 = n71277 & ~n71279;
  assign n71281 = ~P2_P2_INSTADDRPOINTER_REG_11_ & ~n70915;
  assign n71282 = P2_P2_INSTADDRPOINTER_REG_11_ & n70915;
  assign n71283 = ~n71281 & ~n71282;
  assign n71284 = n71280 & ~n71283;
  assign n71285 = ~n71280 & n71283;
  assign n71286 = ~n71284 & ~n71285;
  assign n71287 = n70085 & ~n71286;
  assign n71288 = n68173 & ~n71253;
  assign n71289 = n68174 & ~n71253;
  assign n71290 = n69988 & ~n71242;
  assign n71291 = n67989 & ~n71253;
  assign n71292 = n69991 & ~n71242;
  assign n71293 = ~n71291 & ~n71292;
  assign n71294 = ~n71288 & ~n71289;
  assign n71295 = ~n71290 & n71294;
  assign n71296 = n71293 & n71295;
  assign n71297 = P2_P2_INSTADDRPOINTER_REG_11_ & ~n71199;
  assign n71298 = ~P2_P2_INSTADDRPOINTER_REG_11_ & n71199;
  assign n71299 = ~n71297 & ~n71298;
  assign n71300 = n70087 & ~n71299;
  assign n71301 = n71275 & ~n71276;
  assign n71302 = ~n71287 & n71301;
  assign n71303 = n71296 & n71302;
  assign n71304 = ~n71300 & n71303;
  assign n71305 = n71272 & n71304;
  assign n71306 = n69980 & ~n71305;
  assign n13341 = ~n71238 | n71306;
  assign n71308 = P2_P2_INSTADDRPOINTER_REG_12_ & n69979;
  assign n71309 = P2_P2_REIP_REG_12_ & n70124;
  assign n71310 = P2_P2_INSTADDRPOINTER_REG_11_ & n71250;
  assign n71311 = ~P2_P2_INSTADDRPOINTER_REG_12_ & n71310;
  assign n71312 = P2_P2_INSTADDRPOINTER_REG_12_ & ~n71310;
  assign n71313 = ~n71311 & ~n71312;
  assign n71314 = n68173 & ~n71313;
  assign n71315 = n68174 & ~n71313;
  assign n71316 = P2_P2_INSTADDRPOINTER_REG_11_ & n71239;
  assign n71317 = ~P2_P2_INSTADDRPOINTER_REG_12_ & n71316;
  assign n71318 = P2_P2_INSTADDRPOINTER_REG_12_ & ~n71316;
  assign n71319 = ~n71317 & ~n71318;
  assign n71320 = n69988 & ~n71319;
  assign n71321 = n67989 & ~n71313;
  assign n71322 = n69991 & ~n71319;
  assign n71323 = ~n71321 & ~n71322;
  assign n71324 = ~n71314 & ~n71315;
  assign n71325 = ~n71320 & n71324;
  assign n71326 = n71323 & n71325;
  assign n71327 = ~n68102 & ~n71319;
  assign n71328 = ~P2_P2_INSTADDRPOINTER_REG_12_ & ~n70915;
  assign n71329 = P2_P2_INSTADDRPOINTER_REG_12_ & n70915;
  assign n71330 = ~n71328 & ~n71329;
  assign n71331 = P2_P2_INSTADDRPOINTER_REG_11_ & ~n70915;
  assign n71332 = ~P2_P2_INSTADDRPOINTER_REG_11_ & n70915;
  assign n71333 = ~n71280 & ~n71332;
  assign n71334 = ~n71331 & ~n71333;
  assign n71335 = ~n71330 & n71334;
  assign n71336 = ~P2_P2_INSTADDRPOINTER_REG_12_ & n70915;
  assign n71337 = P2_P2_INSTADDRPOINTER_REG_12_ & ~n70915;
  assign n71338 = ~n71336 & ~n71337;
  assign n71339 = ~n71334 & ~n71338;
  assign n71340 = ~n71335 & ~n71339;
  assign n71341 = n70085 & ~n71340;
  assign n71342 = n68212 & ~n71319;
  assign n71343 = n68055 & ~n71319;
  assign n71344 = ~n71342 & ~n71343;
  assign n71345 = P2_P2_INSTADDRPOINTER_REG_11_ & n71199;
  assign n71346 = ~P2_P2_INSTADDRPOINTER_REG_12_ & ~n71345;
  assign n71347 = P2_P2_INSTADDRPOINTER_REG_11_ & P2_P2_INSTADDRPOINTER_REG_12_;
  assign n71348 = n71199 & n71347;
  assign n71349 = ~n71346 & ~n71348;
  assign n71350 = n70087 & n71349;
  assign n71351 = n71344 & ~n71350;
  assign n71352 = n70104 & ~n71319;
  assign n71353 = n68059 & ~n71319;
  assign n71354 = n70093 & ~n71319;
  assign n71355 = n70097 & ~n71319;
  assign n71356 = ~n71352 & ~n71353;
  assign n71357 = ~n71354 & n71356;
  assign n71358 = ~n71355 & n71357;
  assign n71359 = n67915 & ~n71313;
  assign n71360 = n67993 & ~n71313;
  assign n71361 = n67997 & ~n71313;
  assign n71362 = P2_P2_INSTADDRPOINTER_REG_11_ & n71257;
  assign n71363 = ~P2_P2_INSTADDRPOINTER_REG_12_ & n71362;
  assign n71364 = P2_P2_INSTADDRPOINTER_REG_12_ & ~n71362;
  assign n71365 = ~n71363 & ~n71364;
  assign n71366 = n68013 & ~n71365;
  assign n71367 = n68005 & ~n71365;
  assign n71368 = ~n71359 & ~n71360;
  assign n71369 = ~n71361 & n71368;
  assign n71370 = ~n71366 & n71369;
  assign n71371 = ~n71367 & n71370;
  assign n71372 = P2_P2_INSTADDRPOINTER_REG_11_ & n71224;
  assign n71373 = ~P2_P2_INSTADDRPOINTER_REG_12_ & ~n71372;
  assign n71374 = n71224 & n71347;
  assign n71375 = ~n71373 & ~n71374;
  assign n71376 = n68016 & n71375;
  assign n71377 = n71358 & n71371;
  assign n71378 = ~n71376 & n71377;
  assign n71379 = n71326 & ~n71327;
  assign n71380 = ~n71341 & n71379;
  assign n71381 = n71351 & n71380;
  assign n71382 = n71378 & n71381;
  assign n71383 = n69980 & ~n71382;
  assign n71384 = ~n71308 & ~n71309;
  assign n13346 = n71383 | ~n71384;
  assign n71386 = P2_P2_INSTADDRPOINTER_REG_13_ & n69979;
  assign n71387 = P2_P2_REIP_REG_13_ & n70124;
  assign n71388 = P2_P2_INSTADDRPOINTER_REG_12_ & n71310;
  assign n71389 = ~P2_P2_INSTADDRPOINTER_REG_13_ & n71388;
  assign n71390 = P2_P2_INSTADDRPOINTER_REG_13_ & ~n71388;
  assign n71391 = ~n71389 & ~n71390;
  assign n71392 = n68173 & ~n71391;
  assign n71393 = n68174 & ~n71391;
  assign n71394 = P2_P2_INSTADDRPOINTER_REG_12_ & n71316;
  assign n71395 = ~P2_P2_INSTADDRPOINTER_REG_13_ & n71394;
  assign n71396 = P2_P2_INSTADDRPOINTER_REG_13_ & ~n71394;
  assign n71397 = ~n71395 & ~n71396;
  assign n71398 = n69988 & ~n71397;
  assign n71399 = n67989 & ~n71391;
  assign n71400 = n69991 & ~n71397;
  assign n71401 = ~n71399 & ~n71400;
  assign n71402 = ~n71392 & ~n71393;
  assign n71403 = ~n71398 & n71402;
  assign n71404 = n71401 & n71403;
  assign n71405 = ~n68102 & ~n71397;
  assign n71406 = P2_P2_INSTADDRPOINTER_REG_13_ & ~n70915;
  assign n71407 = P2_P2_INSTADDRPOINTER_REG_12_ & P2_P2_INSTADDRPOINTER_REG_13_;
  assign n71408 = n70915 & ~n71407;
  assign n71409 = ~n71406 & ~n71408;
  assign n71410 = n71334 & ~n71337;
  assign n71411 = n71409 & ~n71410;
  assign n71412 = ~P2_P2_INSTADDRPOINTER_REG_13_ & ~n70915;
  assign n71413 = P2_P2_INSTADDRPOINTER_REG_13_ & n70915;
  assign n71414 = ~n71412 & ~n71413;
  assign n71415 = ~n71337 & n71414;
  assign n71416 = ~n71334 & ~n71336;
  assign n71417 = n71415 & ~n71416;
  assign n71418 = ~n71411 & ~n71417;
  assign n71419 = n70085 & n71418;
  assign n71420 = n68212 & ~n71397;
  assign n71421 = n68055 & ~n71397;
  assign n71422 = ~n71420 & ~n71421;
  assign n71423 = ~P2_P2_INSTADDRPOINTER_REG_13_ & ~n71348;
  assign n71424 = P2_P2_INSTADDRPOINTER_REG_13_ & n71348;
  assign n71425 = ~n71423 & ~n71424;
  assign n71426 = n70087 & n71425;
  assign n71427 = n71422 & ~n71426;
  assign n71428 = n70104 & ~n71397;
  assign n71429 = n68059 & ~n71397;
  assign n71430 = n70093 & ~n71397;
  assign n71431 = n70097 & ~n71397;
  assign n71432 = ~n71428 & ~n71429;
  assign n71433 = ~n71430 & n71432;
  assign n71434 = ~n71431 & n71433;
  assign n71435 = n67915 & ~n71391;
  assign n71436 = n67993 & ~n71391;
  assign n71437 = n67997 & ~n71391;
  assign n71438 = P2_P2_INSTADDRPOINTER_REG_12_ & n71362;
  assign n71439 = ~P2_P2_INSTADDRPOINTER_REG_13_ & n71438;
  assign n71440 = P2_P2_INSTADDRPOINTER_REG_13_ & ~n71438;
  assign n71441 = ~n71439 & ~n71440;
  assign n71442 = n68013 & ~n71441;
  assign n71443 = n68005 & ~n71441;
  assign n71444 = ~n71435 & ~n71436;
  assign n71445 = ~n71437 & n71444;
  assign n71446 = ~n71442 & n71445;
  assign n71447 = ~n71443 & n71446;
  assign n71448 = ~P2_P2_INSTADDRPOINTER_REG_13_ & ~n71374;
  assign n71449 = P2_P2_INSTADDRPOINTER_REG_13_ & n71374;
  assign n71450 = ~n71448 & ~n71449;
  assign n71451 = n68016 & n71450;
  assign n71452 = n71434 & n71447;
  assign n71453 = ~n71451 & n71452;
  assign n71454 = n71404 & ~n71405;
  assign n71455 = ~n71419 & n71454;
  assign n71456 = n71427 & n71455;
  assign n71457 = n71453 & n71456;
  assign n71458 = n69980 & ~n71457;
  assign n71459 = ~n71386 & ~n71387;
  assign n13351 = n71458 | ~n71459;
  assign n71461 = P2_P2_INSTADDRPOINTER_REG_14_ & n69979;
  assign n71462 = P2_P2_REIP_REG_14_ & n70124;
  assign n71463 = ~n71461 & ~n71462;
  assign n71464 = P2_P2_INSTADDRPOINTER_REG_13_ & n71394;
  assign n71465 = ~P2_P2_INSTADDRPOINTER_REG_14_ & n71464;
  assign n71466 = P2_P2_INSTADDRPOINTER_REG_14_ & ~n71464;
  assign n71467 = ~n71465 & ~n71466;
  assign n71468 = n70104 & ~n71467;
  assign n71469 = n68059 & ~n71467;
  assign n71470 = n70093 & ~n71467;
  assign n71471 = n70097 & ~n71467;
  assign n71472 = ~n71468 & ~n71469;
  assign n71473 = ~n71470 & n71472;
  assign n71474 = ~n71471 & n71473;
  assign n71475 = P2_P2_INSTADDRPOINTER_REG_13_ & n71388;
  assign n71476 = ~P2_P2_INSTADDRPOINTER_REG_14_ & n71475;
  assign n71477 = P2_P2_INSTADDRPOINTER_REG_14_ & ~n71475;
  assign n71478 = ~n71476 & ~n71477;
  assign n71479 = n67915 & ~n71478;
  assign n71480 = n67993 & ~n71478;
  assign n71481 = n67997 & ~n71478;
  assign n71482 = P2_P2_INSTADDRPOINTER_REG_13_ & n71438;
  assign n71483 = ~P2_P2_INSTADDRPOINTER_REG_14_ & n71482;
  assign n71484 = P2_P2_INSTADDRPOINTER_REG_14_ & ~n71482;
  assign n71485 = ~n71483 & ~n71484;
  assign n71486 = n68013 & ~n71485;
  assign n71487 = n68005 & ~n71485;
  assign n71488 = ~n71479 & ~n71480;
  assign n71489 = ~n71481 & n71488;
  assign n71490 = ~n71486 & n71489;
  assign n71491 = ~n71487 & n71490;
  assign n71492 = ~P2_P2_INSTADDRPOINTER_REG_14_ & n71449;
  assign n71493 = P2_P2_INSTADDRPOINTER_REG_14_ & ~n71449;
  assign n71494 = ~n71492 & ~n71493;
  assign n71495 = n68016 & ~n71494;
  assign n71496 = n71474 & n71491;
  assign n71497 = ~n71495 & n71496;
  assign n71498 = n68212 & ~n71467;
  assign n71499 = n68055 & ~n71467;
  assign n71500 = ~n71498 & ~n71499;
  assign n71501 = ~n68102 & ~n71467;
  assign n71502 = n68173 & ~n71478;
  assign n71503 = n68174 & ~n71478;
  assign n71504 = n69988 & ~n71467;
  assign n71505 = n67989 & ~n71478;
  assign n71506 = n69991 & ~n71467;
  assign n71507 = ~n71505 & ~n71506;
  assign n71508 = ~n71502 & ~n71503;
  assign n71509 = ~n71504 & n71508;
  assign n71510 = n71507 & n71509;
  assign n71511 = ~n71337 & ~n71406;
  assign n71512 = ~n71331 & n71511;
  assign n71513 = ~n71332 & ~n71408;
  assign n71514 = ~n71280 & n71513;
  assign n71515 = n71512 & ~n71514;
  assign n71516 = ~P2_P2_INSTADDRPOINTER_REG_14_ & ~n70915;
  assign n71517 = P2_P2_INSTADDRPOINTER_REG_14_ & n70915;
  assign n71518 = ~n71516 & ~n71517;
  assign n71519 = n71515 & ~n71518;
  assign n71520 = ~n71515 & n71518;
  assign n71521 = ~n71519 & ~n71520;
  assign n71522 = n70085 & ~n71521;
  assign n71523 = ~P2_P2_INSTADDRPOINTER_REG_14_ & n71424;
  assign n71524 = P2_P2_INSTADDRPOINTER_REG_14_ & ~n71424;
  assign n71525 = ~n71523 & ~n71524;
  assign n71526 = n70087 & ~n71525;
  assign n71527 = n71500 & ~n71501;
  assign n71528 = n71510 & n71527;
  assign n71529 = ~n71522 & n71528;
  assign n71530 = ~n71526 & n71529;
  assign n71531 = n71497 & n71530;
  assign n71532 = n69980 & ~n71531;
  assign n13356 = ~n71463 | n71532;
  assign n71534 = P2_P2_INSTADDRPOINTER_REG_15_ & n69979;
  assign n71535 = P2_P2_REIP_REG_15_ & n70124;
  assign n71536 = ~n71534 & ~n71535;
  assign n71537 = P2_P2_INSTADDRPOINTER_REG_14_ & n71464;
  assign n71538 = ~P2_P2_INSTADDRPOINTER_REG_15_ & n71537;
  assign n71539 = P2_P2_INSTADDRPOINTER_REG_15_ & ~n71537;
  assign n71540 = ~n71538 & ~n71539;
  assign n71541 = n70104 & ~n71540;
  assign n71542 = n68059 & ~n71540;
  assign n71543 = n70093 & ~n71540;
  assign n71544 = n70097 & ~n71540;
  assign n71545 = ~n71541 & ~n71542;
  assign n71546 = ~n71543 & n71545;
  assign n71547 = ~n71544 & n71546;
  assign n71548 = P2_P2_INSTADDRPOINTER_REG_14_ & n71475;
  assign n71549 = ~P2_P2_INSTADDRPOINTER_REG_15_ & n71548;
  assign n71550 = P2_P2_INSTADDRPOINTER_REG_15_ & ~n71548;
  assign n71551 = ~n71549 & ~n71550;
  assign n71552 = n67915 & ~n71551;
  assign n71553 = n67993 & ~n71551;
  assign n71554 = n67997 & ~n71551;
  assign n71555 = P2_P2_INSTADDRPOINTER_REG_14_ & n71482;
  assign n71556 = ~P2_P2_INSTADDRPOINTER_REG_15_ & n71555;
  assign n71557 = P2_P2_INSTADDRPOINTER_REG_15_ & ~n71555;
  assign n71558 = ~n71556 & ~n71557;
  assign n71559 = n68013 & ~n71558;
  assign n71560 = n68005 & ~n71558;
  assign n71561 = ~n71552 & ~n71553;
  assign n71562 = ~n71554 & n71561;
  assign n71563 = ~n71559 & n71562;
  assign n71564 = ~n71560 & n71563;
  assign n71565 = P2_P2_INSTADDRPOINTER_REG_14_ & n71449;
  assign n71566 = ~P2_P2_INSTADDRPOINTER_REG_15_ & ~n71565;
  assign n71567 = P2_P2_INSTADDRPOINTER_REG_14_ & P2_P2_INSTADDRPOINTER_REG_15_;
  assign n71568 = P2_P2_INSTADDRPOINTER_REG_13_ & n71567;
  assign n71569 = n71374 & n71568;
  assign n71570 = ~n71566 & ~n71569;
  assign n71571 = n68016 & n71570;
  assign n71572 = n71547 & n71564;
  assign n71573 = ~n71571 & n71572;
  assign n71574 = n68212 & ~n71540;
  assign n71575 = n68055 & ~n71540;
  assign n71576 = ~n71574 & ~n71575;
  assign n71577 = ~n68102 & ~n71540;
  assign n71578 = n68173 & ~n71551;
  assign n71579 = n68174 & ~n71551;
  assign n71580 = n69988 & ~n71540;
  assign n71581 = n67989 & ~n71551;
  assign n71582 = n69991 & ~n71540;
  assign n71583 = ~n71581 & ~n71582;
  assign n71584 = ~n71578 & ~n71579;
  assign n71585 = ~n71580 & n71584;
  assign n71586 = n71583 & n71585;
  assign n71587 = P2_P2_INSTADDRPOINTER_REG_14_ & ~n70915;
  assign n71588 = n71512 & ~n71587;
  assign n71589 = ~P2_P2_INSTADDRPOINTER_REG_14_ & n70915;
  assign n71590 = n71513 & ~n71589;
  assign n71591 = ~n71280 & n71590;
  assign n71592 = n71588 & ~n71591;
  assign n71593 = ~P2_P2_INSTADDRPOINTER_REG_15_ & ~n70915;
  assign n71594 = P2_P2_INSTADDRPOINTER_REG_15_ & n70915;
  assign n71595 = ~n71593 & ~n71594;
  assign n71596 = n71592 & ~n71595;
  assign n71597 = ~n71592 & n71595;
  assign n71598 = ~n71596 & ~n71597;
  assign n71599 = n70085 & ~n71598;
  assign n71600 = P2_P2_INSTADDRPOINTER_REG_14_ & n71424;
  assign n71601 = ~P2_P2_INSTADDRPOINTER_REG_15_ & ~n71600;
  assign n71602 = n71348 & n71568;
  assign n71603 = ~n71601 & ~n71602;
  assign n71604 = n70087 & n71603;
  assign n71605 = n71576 & ~n71577;
  assign n71606 = n71586 & n71605;
  assign n71607 = ~n71599 & n71606;
  assign n71608 = ~n71604 & n71607;
  assign n71609 = n71573 & n71608;
  assign n71610 = n69980 & ~n71609;
  assign n13361 = ~n71536 | n71610;
  assign n71612 = P2_P2_INSTADDRPOINTER_REG_16_ & n69979;
  assign n71613 = P2_P2_REIP_REG_16_ & n70124;
  assign n71614 = ~n71612 & ~n71613;
  assign n71615 = P2_P2_INSTADDRPOINTER_REG_15_ & n71537;
  assign n71616 = ~P2_P2_INSTADDRPOINTER_REG_16_ & n71615;
  assign n71617 = P2_P2_INSTADDRPOINTER_REG_16_ & ~n71615;
  assign n71618 = ~n71616 & ~n71617;
  assign n71619 = n70104 & ~n71618;
  assign n71620 = n68059 & ~n71618;
  assign n71621 = n70093 & ~n71618;
  assign n71622 = n70097 & ~n71618;
  assign n71623 = ~n71619 & ~n71620;
  assign n71624 = ~n71621 & n71623;
  assign n71625 = ~n71622 & n71624;
  assign n71626 = P2_P2_INSTADDRPOINTER_REG_15_ & n71548;
  assign n71627 = ~P2_P2_INSTADDRPOINTER_REG_16_ & n71626;
  assign n71628 = P2_P2_INSTADDRPOINTER_REG_16_ & ~n71626;
  assign n71629 = ~n71627 & ~n71628;
  assign n71630 = n67915 & ~n71629;
  assign n71631 = n67993 & ~n71629;
  assign n71632 = n67997 & ~n71629;
  assign n71633 = P2_P2_INSTADDRPOINTER_REG_15_ & n71555;
  assign n71634 = ~P2_P2_INSTADDRPOINTER_REG_16_ & n71633;
  assign n71635 = P2_P2_INSTADDRPOINTER_REG_16_ & ~n71633;
  assign n71636 = ~n71634 & ~n71635;
  assign n71637 = n68013 & ~n71636;
  assign n71638 = n68005 & ~n71636;
  assign n71639 = ~n71630 & ~n71631;
  assign n71640 = ~n71632 & n71639;
  assign n71641 = ~n71637 & n71640;
  assign n71642 = ~n71638 & n71641;
  assign n71643 = ~P2_P2_INSTADDRPOINTER_REG_16_ & n71569;
  assign n71644 = P2_P2_INSTADDRPOINTER_REG_16_ & ~n71569;
  assign n71645 = ~n71643 & ~n71644;
  assign n71646 = n68016 & ~n71645;
  assign n71647 = n71625 & n71642;
  assign n71648 = ~n71646 & n71647;
  assign n71649 = n68212 & ~n71618;
  assign n71650 = n68055 & ~n71618;
  assign n71651 = ~n71649 & ~n71650;
  assign n71652 = ~n68102 & ~n71618;
  assign n71653 = P2_P2_INSTADDRPOINTER_REG_15_ & ~n70915;
  assign n71654 = ~P2_P2_INSTADDRPOINTER_REG_15_ & n70915;
  assign n71655 = ~n71592 & ~n71654;
  assign n71656 = ~n71653 & ~n71655;
  assign n71657 = ~P2_P2_INSTADDRPOINTER_REG_16_ & ~n70915;
  assign n71658 = P2_P2_INSTADDRPOINTER_REG_16_ & n70915;
  assign n71659 = ~n71657 & ~n71658;
  assign n71660 = n71656 & ~n71659;
  assign n71661 = ~n71656 & n71659;
  assign n71662 = ~n71660 & ~n71661;
  assign n71663 = n70085 & ~n71662;
  assign n71664 = n68173 & ~n71629;
  assign n71665 = n68174 & ~n71629;
  assign n71666 = n69988 & ~n71618;
  assign n71667 = n67989 & ~n71629;
  assign n71668 = n69991 & ~n71618;
  assign n71669 = ~n71667 & ~n71668;
  assign n71670 = ~n71664 & ~n71665;
  assign n71671 = ~n71666 & n71670;
  assign n71672 = n71669 & n71671;
  assign n71673 = ~P2_P2_INSTADDRPOINTER_REG_16_ & n71602;
  assign n71674 = P2_P2_INSTADDRPOINTER_REG_16_ & ~n71602;
  assign n71675 = ~n71673 & ~n71674;
  assign n71676 = n70087 & ~n71675;
  assign n71677 = n71651 & ~n71652;
  assign n71678 = ~n71663 & n71677;
  assign n71679 = n71672 & n71678;
  assign n71680 = ~n71676 & n71679;
  assign n71681 = n71648 & n71680;
  assign n71682 = n69980 & ~n71681;
  assign n13366 = ~n71614 | n71682;
  assign n71684 = P2_P2_INSTADDRPOINTER_REG_17_ & n69979;
  assign n71685 = P2_P2_REIP_REG_17_ & n70124;
  assign n71686 = P2_P2_INSTADDRPOINTER_REG_16_ & n71626;
  assign n71687 = ~P2_P2_INSTADDRPOINTER_REG_17_ & n71686;
  assign n71688 = P2_P2_INSTADDRPOINTER_REG_17_ & ~n71686;
  assign n71689 = ~n71687 & ~n71688;
  assign n71690 = n68173 & ~n71689;
  assign n71691 = n68174 & ~n71689;
  assign n71692 = P2_P2_INSTADDRPOINTER_REG_16_ & n71615;
  assign n71693 = ~P2_P2_INSTADDRPOINTER_REG_17_ & n71692;
  assign n71694 = P2_P2_INSTADDRPOINTER_REG_17_ & ~n71692;
  assign n71695 = ~n71693 & ~n71694;
  assign n71696 = n69988 & ~n71695;
  assign n71697 = n67989 & ~n71689;
  assign n71698 = n69991 & ~n71695;
  assign n71699 = ~n71697 & ~n71698;
  assign n71700 = ~n71690 & ~n71691;
  assign n71701 = ~n71696 & n71700;
  assign n71702 = n71699 & n71701;
  assign n71703 = ~n68102 & ~n71695;
  assign n71704 = P2_P2_INSTADDRPOINTER_REG_16_ & P2_P2_INSTADDRPOINTER_REG_17_;
  assign n71705 = ~n71656 & n71704;
  assign n71706 = n70915 & ~n71705;
  assign n71707 = P2_P2_INSTADDRPOINTER_REG_17_ & ~n70915;
  assign n71708 = ~P2_P2_INSTADDRPOINTER_REG_16_ & ~n71653;
  assign n71709 = ~n71655 & n71708;
  assign n71710 = ~n71706 & ~n71707;
  assign n71711 = ~n71709 & n71710;
  assign n71712 = P2_P2_INSTADDRPOINTER_REG_17_ & n71709;
  assign n71713 = ~n70915 & ~n71712;
  assign n71714 = P2_P2_INSTADDRPOINTER_REG_17_ & n70915;
  assign n71715 = P2_P2_INSTADDRPOINTER_REG_16_ & ~n71656;
  assign n71716 = ~n71713 & ~n71714;
  assign n71717 = ~n71715 & n71716;
  assign n71718 = ~n71711 & ~n71717;
  assign n71719 = n70085 & n71718;
  assign n71720 = n68212 & ~n71695;
  assign n71721 = n68055 & ~n71695;
  assign n71722 = ~n71720 & ~n71721;
  assign n71723 = P2_P2_INSTADDRPOINTER_REG_16_ & n71602;
  assign n71724 = ~P2_P2_INSTADDRPOINTER_REG_17_ & ~n71723;
  assign n71725 = n71602 & n71704;
  assign n71726 = ~n71724 & ~n71725;
  assign n71727 = n70087 & n71726;
  assign n71728 = n71722 & ~n71727;
  assign n71729 = n70104 & ~n71695;
  assign n71730 = n68059 & ~n71695;
  assign n71731 = n70093 & ~n71695;
  assign n71732 = n70097 & ~n71695;
  assign n71733 = ~n71729 & ~n71730;
  assign n71734 = ~n71731 & n71733;
  assign n71735 = ~n71732 & n71734;
  assign n71736 = n67915 & ~n71689;
  assign n71737 = n67993 & ~n71689;
  assign n71738 = n67997 & ~n71689;
  assign n71739 = P2_P2_INSTADDRPOINTER_REG_16_ & n71633;
  assign n71740 = ~P2_P2_INSTADDRPOINTER_REG_17_ & n71739;
  assign n71741 = P2_P2_INSTADDRPOINTER_REG_17_ & ~n71739;
  assign n71742 = ~n71740 & ~n71741;
  assign n71743 = n68013 & ~n71742;
  assign n71744 = n68005 & ~n71742;
  assign n71745 = ~n71736 & ~n71737;
  assign n71746 = ~n71738 & n71745;
  assign n71747 = ~n71743 & n71746;
  assign n71748 = ~n71744 & n71747;
  assign n71749 = P2_P2_INSTADDRPOINTER_REG_16_ & n71569;
  assign n71750 = ~P2_P2_INSTADDRPOINTER_REG_17_ & ~n71749;
  assign n71751 = n71569 & n71704;
  assign n71752 = ~n71750 & ~n71751;
  assign n71753 = n68016 & n71752;
  assign n71754 = n71735 & n71748;
  assign n71755 = ~n71753 & n71754;
  assign n71756 = n71702 & ~n71703;
  assign n71757 = ~n71719 & n71756;
  assign n71758 = n71728 & n71757;
  assign n71759 = n71755 & n71758;
  assign n71760 = n69980 & ~n71759;
  assign n71761 = ~n71684 & ~n71685;
  assign n13371 = n71760 | ~n71761;
  assign n71763 = P2_P2_INSTADDRPOINTER_REG_18_ & n69979;
  assign n71764 = P2_P2_REIP_REG_18_ & n70124;
  assign n71765 = ~n71763 & ~n71764;
  assign n71766 = P2_P2_INSTADDRPOINTER_REG_17_ & n71692;
  assign n71767 = ~P2_P2_INSTADDRPOINTER_REG_18_ & n71766;
  assign n71768 = P2_P2_INSTADDRPOINTER_REG_18_ & ~n71766;
  assign n71769 = ~n71767 & ~n71768;
  assign n71770 = n70104 & ~n71769;
  assign n71771 = n68059 & ~n71769;
  assign n71772 = n70093 & ~n71769;
  assign n71773 = n70097 & ~n71769;
  assign n71774 = ~n71770 & ~n71771;
  assign n71775 = ~n71772 & n71774;
  assign n71776 = ~n71773 & n71775;
  assign n71777 = P2_P2_INSTADDRPOINTER_REG_17_ & n71686;
  assign n71778 = ~P2_P2_INSTADDRPOINTER_REG_18_ & n71777;
  assign n71779 = P2_P2_INSTADDRPOINTER_REG_18_ & ~n71777;
  assign n71780 = ~n71778 & ~n71779;
  assign n71781 = n67915 & ~n71780;
  assign n71782 = n67993 & ~n71780;
  assign n71783 = n67997 & ~n71780;
  assign n71784 = P2_P2_INSTADDRPOINTER_REG_17_ & n71739;
  assign n71785 = ~P2_P2_INSTADDRPOINTER_REG_18_ & n71784;
  assign n71786 = P2_P2_INSTADDRPOINTER_REG_18_ & ~n71784;
  assign n71787 = ~n71785 & ~n71786;
  assign n71788 = n68013 & ~n71787;
  assign n71789 = n68005 & ~n71787;
  assign n71790 = ~n71781 & ~n71782;
  assign n71791 = ~n71783 & n71790;
  assign n71792 = ~n71788 & n71791;
  assign n71793 = ~n71789 & n71792;
  assign n71794 = ~P2_P2_INSTADDRPOINTER_REG_18_ & n71751;
  assign n71795 = P2_P2_INSTADDRPOINTER_REG_18_ & ~n71751;
  assign n71796 = ~n71794 & ~n71795;
  assign n71797 = n68016 & ~n71796;
  assign n71798 = n71776 & n71793;
  assign n71799 = ~n71797 & n71798;
  assign n71800 = n68212 & ~n71769;
  assign n71801 = n68055 & ~n71769;
  assign n71802 = ~n71800 & ~n71801;
  assign n71803 = ~n68102 & ~n71769;
  assign n71804 = ~n70915 & ~n71709;
  assign n71805 = ~n71705 & ~n71804;
  assign n71806 = ~n71707 & n71805;
  assign n71807 = ~P2_P2_INSTADDRPOINTER_REG_18_ & ~n70915;
  assign n71808 = P2_P2_INSTADDRPOINTER_REG_18_ & n70915;
  assign n71809 = ~n71807 & ~n71808;
  assign n71810 = n71806 & ~n71809;
  assign n71811 = ~n71806 & n71809;
  assign n71812 = ~n71810 & ~n71811;
  assign n71813 = n70085 & ~n71812;
  assign n71814 = n68173 & ~n71780;
  assign n71815 = n68174 & ~n71780;
  assign n71816 = n69988 & ~n71769;
  assign n71817 = n67989 & ~n71780;
  assign n71818 = n69991 & ~n71769;
  assign n71819 = ~n71817 & ~n71818;
  assign n71820 = ~n71814 & ~n71815;
  assign n71821 = ~n71816 & n71820;
  assign n71822 = n71819 & n71821;
  assign n71823 = ~P2_P2_INSTADDRPOINTER_REG_18_ & n71725;
  assign n71824 = P2_P2_INSTADDRPOINTER_REG_18_ & ~n71725;
  assign n71825 = ~n71823 & ~n71824;
  assign n71826 = n70087 & ~n71825;
  assign n71827 = n71802 & ~n71803;
  assign n71828 = ~n71813 & n71827;
  assign n71829 = n71822 & n71828;
  assign n71830 = ~n71826 & n71829;
  assign n71831 = n71799 & n71830;
  assign n71832 = n69980 & ~n71831;
  assign n13376 = ~n71765 | n71832;
  assign n71834 = P2_P2_INSTADDRPOINTER_REG_19_ & n69979;
  assign n71835 = P2_P2_REIP_REG_19_ & n70124;
  assign n71836 = P2_P2_INSTADDRPOINTER_REG_18_ & n71777;
  assign n71837 = ~P2_P2_INSTADDRPOINTER_REG_19_ & n71836;
  assign n71838 = P2_P2_INSTADDRPOINTER_REG_19_ & ~n71836;
  assign n71839 = ~n71837 & ~n71838;
  assign n71840 = n68173 & ~n71839;
  assign n71841 = n68174 & ~n71839;
  assign n71842 = P2_P2_INSTADDRPOINTER_REG_18_ & n71766;
  assign n71843 = ~P2_P2_INSTADDRPOINTER_REG_19_ & n71842;
  assign n71844 = P2_P2_INSTADDRPOINTER_REG_19_ & ~n71842;
  assign n71845 = ~n71843 & ~n71844;
  assign n71846 = n69988 & ~n71845;
  assign n71847 = n67989 & ~n71839;
  assign n71848 = n69991 & ~n71845;
  assign n71849 = ~n71847 & ~n71848;
  assign n71850 = ~n71840 & ~n71841;
  assign n71851 = ~n71846 & n71850;
  assign n71852 = n71849 & n71851;
  assign n71853 = ~n68102 & ~n71845;
  assign n71854 = ~P2_P2_INSTADDRPOINTER_REG_19_ & ~n70915;
  assign n71855 = P2_P2_INSTADDRPOINTER_REG_19_ & n70915;
  assign n71856 = ~n71854 & ~n71855;
  assign n71857 = ~P2_P2_INSTADDRPOINTER_REG_18_ & n70915;
  assign n71858 = ~n71806 & ~n71857;
  assign n71859 = P2_P2_INSTADDRPOINTER_REG_18_ & ~n70915;
  assign n71860 = ~n71858 & ~n71859;
  assign n71861 = ~n71856 & n71860;
  assign n71862 = ~P2_P2_INSTADDRPOINTER_REG_19_ & n70915;
  assign n71863 = P2_P2_INSTADDRPOINTER_REG_19_ & ~n70915;
  assign n71864 = ~n71862 & ~n71863;
  assign n71865 = ~n71860 & ~n71864;
  assign n71866 = ~n71861 & ~n71865;
  assign n71867 = n70085 & ~n71866;
  assign n71868 = n68212 & ~n71845;
  assign n71869 = n68055 & ~n71845;
  assign n71870 = ~n71868 & ~n71869;
  assign n71871 = P2_P2_INSTADDRPOINTER_REG_18_ & n71725;
  assign n71872 = ~P2_P2_INSTADDRPOINTER_REG_19_ & ~n71871;
  assign n71873 = P2_P2_INSTADDRPOINTER_REG_18_ & P2_P2_INSTADDRPOINTER_REG_19_;
  assign n71874 = n71725 & n71873;
  assign n71875 = ~n71872 & ~n71874;
  assign n71876 = n70087 & n71875;
  assign n71877 = n71870 & ~n71876;
  assign n71878 = n70104 & ~n71845;
  assign n71879 = n68059 & ~n71845;
  assign n71880 = n70093 & ~n71845;
  assign n71881 = n70097 & ~n71845;
  assign n71882 = ~n71878 & ~n71879;
  assign n71883 = ~n71880 & n71882;
  assign n71884 = ~n71881 & n71883;
  assign n71885 = n67915 & ~n71839;
  assign n71886 = n67993 & ~n71839;
  assign n71887 = n67997 & ~n71839;
  assign n71888 = P2_P2_INSTADDRPOINTER_REG_18_ & n71784;
  assign n71889 = ~P2_P2_INSTADDRPOINTER_REG_19_ & n71888;
  assign n71890 = P2_P2_INSTADDRPOINTER_REG_19_ & ~n71888;
  assign n71891 = ~n71889 & ~n71890;
  assign n71892 = n68013 & ~n71891;
  assign n71893 = n68005 & ~n71891;
  assign n71894 = ~n71885 & ~n71886;
  assign n71895 = ~n71887 & n71894;
  assign n71896 = ~n71892 & n71895;
  assign n71897 = ~n71893 & n71896;
  assign n71898 = P2_P2_INSTADDRPOINTER_REG_18_ & n71751;
  assign n71899 = ~P2_P2_INSTADDRPOINTER_REG_19_ & ~n71898;
  assign n71900 = n71751 & n71873;
  assign n71901 = ~n71899 & ~n71900;
  assign n71902 = n68016 & n71901;
  assign n71903 = n71884 & n71897;
  assign n71904 = ~n71902 & n71903;
  assign n71905 = n71852 & ~n71853;
  assign n71906 = ~n71867 & n71905;
  assign n71907 = n71877 & n71906;
  assign n71908 = n71904 & n71907;
  assign n71909 = n69980 & ~n71908;
  assign n71910 = ~n71834 & ~n71835;
  assign n13381 = n71909 | ~n71910;
  assign n71912 = P2_P2_INSTADDRPOINTER_REG_20_ & n69979;
  assign n71913 = P2_P2_REIP_REG_20_ & n70124;
  assign n71914 = ~n71912 & ~n71913;
  assign n71915 = P2_P2_INSTADDRPOINTER_REG_19_ & P2_P2_INSTADDRPOINTER_REG_20_;
  assign n71916 = n70915 & ~n71915;
  assign n71917 = P2_P2_INSTADDRPOINTER_REG_20_ & ~n70915;
  assign n71918 = ~n71916 & ~n71917;
  assign n71919 = n71860 & ~n71863;
  assign n71920 = n71918 & ~n71919;
  assign n71921 = ~P2_P2_INSTADDRPOINTER_REG_19_ & n71860;
  assign n71922 = P2_P2_INSTADDRPOINTER_REG_20_ & n71921;
  assign n71923 = ~n70915 & ~n71922;
  assign n71924 = P2_P2_INSTADDRPOINTER_REG_20_ & n70915;
  assign n71925 = P2_P2_INSTADDRPOINTER_REG_19_ & ~n71860;
  assign n71926 = ~n71923 & ~n71924;
  assign n71927 = ~n71925 & n71926;
  assign n71928 = ~n71920 & ~n71927;
  assign n71929 = n70085 & n71928;
  assign n71930 = P2_P2_INSTADDRPOINTER_REG_19_ & n71842;
  assign n71931 = ~P2_P2_INSTADDRPOINTER_REG_20_ & n71930;
  assign n71932 = P2_P2_INSTADDRPOINTER_REG_20_ & ~n71930;
  assign n71933 = ~n71931 & ~n71932;
  assign n71934 = ~n68102 & ~n71933;
  assign n71935 = n68212 & ~n71933;
  assign n71936 = n68055 & ~n71933;
  assign n71937 = ~n71935 & ~n71936;
  assign n71938 = P2_P2_INSTADDRPOINTER_REG_19_ & n71836;
  assign n71939 = ~P2_P2_INSTADDRPOINTER_REG_20_ & n71938;
  assign n71940 = P2_P2_INSTADDRPOINTER_REG_20_ & ~n71938;
  assign n71941 = ~n71939 & ~n71940;
  assign n71942 = n68173 & ~n71941;
  assign n71943 = n68174 & ~n71941;
  assign n71944 = n69988 & ~n71933;
  assign n71945 = n67989 & ~n71941;
  assign n71946 = n69991 & ~n71933;
  assign n71947 = ~n71945 & ~n71946;
  assign n71948 = ~n71942 & ~n71943;
  assign n71949 = ~n71944 & n71948;
  assign n71950 = n71947 & n71949;
  assign n71951 = ~P2_P2_INSTADDRPOINTER_REG_20_ & ~n71874;
  assign n71952 = P2_P2_INSTADDRPOINTER_REG_20_ & n71874;
  assign n71953 = ~n71951 & ~n71952;
  assign n71954 = n70087 & n71953;
  assign n71955 = n70104 & ~n71933;
  assign n71956 = n68059 & ~n71933;
  assign n71957 = n70093 & ~n71933;
  assign n71958 = n70097 & ~n71933;
  assign n71959 = ~n71955 & ~n71956;
  assign n71960 = ~n71957 & n71959;
  assign n71961 = ~n71958 & n71960;
  assign n71962 = n67915 & ~n71941;
  assign n71963 = n67993 & ~n71941;
  assign n71964 = n67997 & ~n71941;
  assign n71965 = P2_P2_INSTADDRPOINTER_REG_19_ & n71888;
  assign n71966 = ~P2_P2_INSTADDRPOINTER_REG_20_ & n71965;
  assign n71967 = P2_P2_INSTADDRPOINTER_REG_20_ & ~n71965;
  assign n71968 = ~n71966 & ~n71967;
  assign n71969 = n68013 & ~n71968;
  assign n71970 = n68005 & ~n71968;
  assign n71971 = ~n71962 & ~n71963;
  assign n71972 = ~n71964 & n71971;
  assign n71973 = ~n71969 & n71972;
  assign n71974 = ~n71970 & n71973;
  assign n71975 = ~P2_P2_INSTADDRPOINTER_REG_20_ & ~n71900;
  assign n71976 = P2_P2_INSTADDRPOINTER_REG_20_ & n71900;
  assign n71977 = ~n71975 & ~n71976;
  assign n71978 = n68016 & n71977;
  assign n71979 = n71961 & n71974;
  assign n71980 = ~n71978 & n71979;
  assign n71981 = ~n71934 & n71937;
  assign n71982 = n71950 & n71981;
  assign n71983 = ~n71954 & n71982;
  assign n71984 = n71980 & n71983;
  assign n71985 = ~n71929 & n71984;
  assign n71986 = n69980 & ~n71985;
  assign n13386 = ~n71914 | n71986;
  assign n71988 = P2_P2_INSTADDRPOINTER_REG_21_ & n69979;
  assign n71989 = P2_P2_REIP_REG_21_ & n70124;
  assign n71990 = P2_P2_INSTADDRPOINTER_REG_20_ & n71930;
  assign n71991 = ~P2_P2_INSTADDRPOINTER_REG_21_ & n71990;
  assign n71992 = P2_P2_INSTADDRPOINTER_REG_21_ & ~n71990;
  assign n71993 = ~n71991 & ~n71992;
  assign n71994 = ~n68102 & ~n71993;
  assign n71995 = P2_P2_INSTADDRPOINTER_REG_20_ & n71938;
  assign n71996 = ~P2_P2_INSTADDRPOINTER_REG_21_ & n71995;
  assign n71997 = P2_P2_INSTADDRPOINTER_REG_21_ & ~n71995;
  assign n71998 = ~n71996 & ~n71997;
  assign n71999 = n68173 & ~n71998;
  assign n72000 = n68174 & ~n71998;
  assign n72001 = n69988 & ~n71993;
  assign n72002 = n67989 & ~n71998;
  assign n72003 = n69991 & ~n71993;
  assign n72004 = ~n72002 & ~n72003;
  assign n72005 = ~n71999 & ~n72000;
  assign n72006 = ~n72001 & n72005;
  assign n72007 = n72004 & n72006;
  assign n72008 = ~P2_P2_INSTADDRPOINTER_REG_21_ & ~n71952;
  assign n72009 = P2_P2_INSTADDRPOINTER_REG_21_ & n71952;
  assign n72010 = ~n72008 & ~n72009;
  assign n72011 = n70087 & n72010;
  assign n72012 = n67915 & ~n71998;
  assign n72013 = n67993 & ~n71998;
  assign n72014 = n67997 & ~n71998;
  assign n72015 = P2_P2_INSTADDRPOINTER_REG_20_ & n71965;
  assign n72016 = ~P2_P2_INSTADDRPOINTER_REG_21_ & n72015;
  assign n72017 = P2_P2_INSTADDRPOINTER_REG_21_ & ~n72015;
  assign n72018 = ~n72016 & ~n72017;
  assign n72019 = n68013 & ~n72018;
  assign n72020 = n68005 & ~n72018;
  assign n72021 = ~n72012 & ~n72013;
  assign n72022 = ~n72014 & n72021;
  assign n72023 = ~n72019 & n72022;
  assign n72024 = ~n72020 & n72023;
  assign n72025 = n70104 & ~n71993;
  assign n72026 = n68059 & ~n71993;
  assign n72027 = n70093 & ~n71993;
  assign n72028 = n70097 & ~n71993;
  assign n72029 = ~n72025 & ~n72026;
  assign n72030 = ~n72027 & n72029;
  assign n72031 = ~n72028 & n72030;
  assign n72032 = ~P2_P2_INSTADDRPOINTER_REG_21_ & ~n71976;
  assign n72033 = P2_P2_INSTADDRPOINTER_REG_20_ & P2_P2_INSTADDRPOINTER_REG_21_;
  assign n72034 = n71900 & n72033;
  assign n72035 = ~n72032 & ~n72034;
  assign n72036 = n68016 & n72035;
  assign n72037 = n72024 & n72031;
  assign n72038 = ~n72036 & n72037;
  assign n72039 = n68212 & ~n71993;
  assign n72040 = n68055 & ~n71993;
  assign n72041 = ~n72039 & ~n72040;
  assign n72042 = ~n71860 & n71915;
  assign n72043 = ~n71917 & ~n72042;
  assign n72044 = ~n70915 & ~n71921;
  assign n72045 = n72043 & ~n72044;
  assign n72046 = ~P2_P2_INSTADDRPOINTER_REG_21_ & ~n70915;
  assign n72047 = P2_P2_INSTADDRPOINTER_REG_21_ & n70915;
  assign n72048 = ~n72046 & ~n72047;
  assign n72049 = n72045 & ~n72048;
  assign n72050 = ~n72045 & n72048;
  assign n72051 = ~n72049 & ~n72050;
  assign n72052 = n70085 & ~n72051;
  assign n72053 = n72041 & ~n72052;
  assign n72054 = ~n71994 & n72007;
  assign n72055 = ~n72011 & n72054;
  assign n72056 = n72038 & n72055;
  assign n72057 = n72053 & n72056;
  assign n72058 = n69980 & ~n72057;
  assign n72059 = ~n71988 & ~n71989;
  assign n13391 = n72058 | ~n72059;
  assign n72061 = P2_P2_INSTADDRPOINTER_REG_22_ & n69979;
  assign n72062 = P2_P2_REIP_REG_22_ & n70124;
  assign n72063 = ~n72061 & ~n72062;
  assign n72064 = P2_P2_INSTADDRPOINTER_REG_21_ & n72015;
  assign n72065 = ~P2_P2_INSTADDRPOINTER_REG_22_ & n72064;
  assign n72066 = P2_P2_INSTADDRPOINTER_REG_22_ & ~n72064;
  assign n72067 = ~n72065 & ~n72066;
  assign n72068 = n68013 & ~n72067;
  assign n72069 = n68005 & ~n72067;
  assign n72070 = ~n72068 & ~n72069;
  assign n72071 = P2_P2_INSTADDRPOINTER_REG_21_ & n71995;
  assign n72072 = ~P2_P2_INSTADDRPOINTER_REG_22_ & n72071;
  assign n72073 = P2_P2_INSTADDRPOINTER_REG_22_ & ~n72071;
  assign n72074 = ~n72072 & ~n72073;
  assign n72075 = n67915 & ~n72074;
  assign n72076 = n67993 & ~n72074;
  assign n72077 = n67997 & ~n72074;
  assign n72078 = ~n72075 & ~n72076;
  assign n72079 = ~n72077 & n72078;
  assign n72080 = P2_P2_INSTADDRPOINTER_REG_21_ & n71990;
  assign n72081 = ~P2_P2_INSTADDRPOINTER_REG_22_ & n72080;
  assign n72082 = P2_P2_INSTADDRPOINTER_REG_22_ & ~n72080;
  assign n72083 = ~n72081 & ~n72082;
  assign n72084 = n70093 & ~n72083;
  assign n72085 = n70097 & ~n72083;
  assign n72086 = n68059 & ~n72083;
  assign n72087 = ~n72084 & ~n72085;
  assign n72088 = ~n72086 & n72087;
  assign n72089 = ~P2_P2_INSTADDRPOINTER_REG_22_ & n72034;
  assign n72090 = P2_P2_INSTADDRPOINTER_REG_22_ & ~n72034;
  assign n72091 = ~n72089 & ~n72090;
  assign n72092 = n68016 & ~n72091;
  assign n72093 = n70104 & ~n72083;
  assign n72094 = ~n72092 & ~n72093;
  assign n72095 = n72070 & n72079;
  assign n72096 = n72088 & n72095;
  assign n72097 = n72094 & n72096;
  assign n72098 = P2_P2_INSTADDRPOINTER_REG_21_ & n71915;
  assign n72099 = n70915 & ~n72098;
  assign n72100 = ~n71857 & ~n72099;
  assign n72101 = ~n71806 & n72100;
  assign n72102 = P2_P2_INSTADDRPOINTER_REG_21_ & ~n70915;
  assign n72103 = ~n71859 & ~n72102;
  assign n72104 = ~n71863 & n72103;
  assign n72105 = ~n71917 & n72104;
  assign n72106 = ~n72101 & n72105;
  assign n72107 = ~P2_P2_INSTADDRPOINTER_REG_22_ & ~n70915;
  assign n72108 = P2_P2_INSTADDRPOINTER_REG_22_ & n70915;
  assign n72109 = ~n72107 & ~n72108;
  assign n72110 = n72106 & ~n72109;
  assign n72111 = ~n72106 & n72109;
  assign n72112 = ~n72110 & ~n72111;
  assign n72113 = n70085 & ~n72112;
  assign n72114 = ~n68102 & ~n72083;
  assign n72115 = n68212 & ~n72083;
  assign n72116 = n68055 & ~n72083;
  assign n72117 = ~n72115 & ~n72116;
  assign n72118 = n68173 & ~n72074;
  assign n72119 = n68174 & ~n72074;
  assign n72120 = n69988 & ~n72083;
  assign n72121 = n67989 & ~n72074;
  assign n72122 = n69991 & ~n72083;
  assign n72123 = ~n72121 & ~n72122;
  assign n72124 = ~n72118 & ~n72119;
  assign n72125 = ~n72120 & n72124;
  assign n72126 = n72123 & n72125;
  assign n72127 = ~P2_P2_INSTADDRPOINTER_REG_22_ & n72009;
  assign n72128 = P2_P2_INSTADDRPOINTER_REG_22_ & ~n72009;
  assign n72129 = ~n72127 & ~n72128;
  assign n72130 = n70087 & ~n72129;
  assign n72131 = ~n72113 & ~n72114;
  assign n72132 = n72117 & n72131;
  assign n72133 = n72126 & n72132;
  assign n72134 = ~n72130 & n72133;
  assign n72135 = n72097 & n72134;
  assign n72136 = n69980 & ~n72135;
  assign n13396 = ~n72063 | n72136;
  assign n72138 = P2_P2_INSTADDRPOINTER_REG_23_ & n69979;
  assign n72139 = P2_P2_REIP_REG_23_ & n70124;
  assign n72140 = ~n72138 & ~n72139;
  assign n72141 = P2_P2_INSTADDRPOINTER_REG_22_ & n72064;
  assign n72142 = ~P2_P2_INSTADDRPOINTER_REG_23_ & n72141;
  assign n72143 = P2_P2_INSTADDRPOINTER_REG_23_ & ~n72141;
  assign n72144 = ~n72142 & ~n72143;
  assign n72145 = n68013 & ~n72144;
  assign n72146 = n68005 & ~n72144;
  assign n72147 = ~n72145 & ~n72146;
  assign n72148 = P2_P2_INSTADDRPOINTER_REG_22_ & n72071;
  assign n72149 = ~P2_P2_INSTADDRPOINTER_REG_23_ & n72148;
  assign n72150 = P2_P2_INSTADDRPOINTER_REG_23_ & ~n72148;
  assign n72151 = ~n72149 & ~n72150;
  assign n72152 = n67915 & ~n72151;
  assign n72153 = n67993 & ~n72151;
  assign n72154 = n67997 & ~n72151;
  assign n72155 = ~n72152 & ~n72153;
  assign n72156 = ~n72154 & n72155;
  assign n72157 = P2_P2_INSTADDRPOINTER_REG_22_ & n72080;
  assign n72158 = ~P2_P2_INSTADDRPOINTER_REG_23_ & n72157;
  assign n72159 = P2_P2_INSTADDRPOINTER_REG_23_ & ~n72157;
  assign n72160 = ~n72158 & ~n72159;
  assign n72161 = n70093 & ~n72160;
  assign n72162 = n70097 & ~n72160;
  assign n72163 = n68059 & ~n72160;
  assign n72164 = ~n72161 & ~n72162;
  assign n72165 = ~n72163 & n72164;
  assign n72166 = P2_P2_INSTADDRPOINTER_REG_22_ & n72034;
  assign n72167 = ~P2_P2_INSTADDRPOINTER_REG_23_ & ~n72166;
  assign n72168 = P2_P2_INSTADDRPOINTER_REG_22_ & P2_P2_INSTADDRPOINTER_REG_23_;
  assign n72169 = n72034 & n72168;
  assign n72170 = ~n72167 & ~n72169;
  assign n72171 = n68016 & n72170;
  assign n72172 = n70104 & ~n72160;
  assign n72173 = ~n72171 & ~n72172;
  assign n72174 = n72147 & n72156;
  assign n72175 = n72165 & n72174;
  assign n72176 = n72173 & n72175;
  assign n72177 = ~P2_P2_INSTADDRPOINTER_REG_22_ & n70915;
  assign n72178 = n72100 & ~n72177;
  assign n72179 = ~n71806 & n72178;
  assign n72180 = P2_P2_INSTADDRPOINTER_REG_22_ & ~n70915;
  assign n72181 = n72105 & ~n72180;
  assign n72182 = ~n72179 & n72181;
  assign n72183 = ~P2_P2_INSTADDRPOINTER_REG_23_ & ~n70915;
  assign n72184 = P2_P2_INSTADDRPOINTER_REG_23_ & n70915;
  assign n72185 = ~n72183 & ~n72184;
  assign n72186 = n72182 & ~n72185;
  assign n72187 = ~n72182 & n72185;
  assign n72188 = ~n72186 & ~n72187;
  assign n72189 = n70085 & ~n72188;
  assign n72190 = ~n68102 & ~n72160;
  assign n72191 = n68212 & ~n72160;
  assign n72192 = n68055 & ~n72160;
  assign n72193 = ~n72191 & ~n72192;
  assign n72194 = n68173 & ~n72151;
  assign n72195 = n68174 & ~n72151;
  assign n72196 = n69988 & ~n72160;
  assign n72197 = n67989 & ~n72151;
  assign n72198 = n69991 & ~n72160;
  assign n72199 = ~n72197 & ~n72198;
  assign n72200 = ~n72194 & ~n72195;
  assign n72201 = ~n72196 & n72200;
  assign n72202 = n72199 & n72201;
  assign n72203 = P2_P2_INSTADDRPOINTER_REG_22_ & n72009;
  assign n72204 = ~P2_P2_INSTADDRPOINTER_REG_23_ & ~n72203;
  assign n72205 = n72009 & n72168;
  assign n72206 = ~n72204 & ~n72205;
  assign n72207 = n70087 & n72206;
  assign n72208 = ~n72189 & ~n72190;
  assign n72209 = n72193 & n72208;
  assign n72210 = n72202 & n72209;
  assign n72211 = ~n72207 & n72210;
  assign n72212 = n72176 & n72211;
  assign n72213 = n69980 & ~n72212;
  assign n13401 = ~n72140 | n72213;
  assign n72215 = P2_P2_INSTADDRPOINTER_REG_24_ & n69979;
  assign n72216 = P2_P2_REIP_REG_24_ & n70124;
  assign n72217 = ~n72215 & ~n72216;
  assign n72218 = P2_P2_INSTADDRPOINTER_REG_23_ & n72141;
  assign n72219 = ~P2_P2_INSTADDRPOINTER_REG_24_ & n72218;
  assign n72220 = P2_P2_INSTADDRPOINTER_REG_24_ & ~n72218;
  assign n72221 = ~n72219 & ~n72220;
  assign n72222 = n68013 & ~n72221;
  assign n72223 = n68005 & ~n72221;
  assign n72224 = ~n72222 & ~n72223;
  assign n72225 = P2_P2_INSTADDRPOINTER_REG_23_ & n72148;
  assign n72226 = ~P2_P2_INSTADDRPOINTER_REG_24_ & n72225;
  assign n72227 = P2_P2_INSTADDRPOINTER_REG_24_ & ~n72225;
  assign n72228 = ~n72226 & ~n72227;
  assign n72229 = n67915 & ~n72228;
  assign n72230 = n67993 & ~n72228;
  assign n72231 = n67997 & ~n72228;
  assign n72232 = ~n72229 & ~n72230;
  assign n72233 = ~n72231 & n72232;
  assign n72234 = ~P2_P2_INSTADDRPOINTER_REG_24_ & n72169;
  assign n72235 = P2_P2_INSTADDRPOINTER_REG_24_ & ~n72169;
  assign n72236 = ~n72234 & ~n72235;
  assign n72237 = n68016 & ~n72236;
  assign n72238 = P2_P2_INSTADDRPOINTER_REG_23_ & n72157;
  assign n72239 = ~P2_P2_INSTADDRPOINTER_REG_24_ & n72238;
  assign n72240 = P2_P2_INSTADDRPOINTER_REG_24_ & ~n72238;
  assign n72241 = ~n72239 & ~n72240;
  assign n72242 = n70104 & ~n72241;
  assign n72243 = ~n72237 & ~n72242;
  assign n72244 = n70093 & ~n72241;
  assign n72245 = n70097 & ~n72241;
  assign n72246 = n68059 & ~n72241;
  assign n72247 = ~n72244 & ~n72245;
  assign n72248 = ~n72246 & n72247;
  assign n72249 = n72224 & n72233;
  assign n72250 = n72243 & n72249;
  assign n72251 = n72248 & n72250;
  assign n72252 = P2_P2_INSTADDRPOINTER_REG_23_ & ~n70915;
  assign n72253 = n72181 & ~n72252;
  assign n72254 = ~P2_P2_INSTADDRPOINTER_REG_23_ & n70915;
  assign n72255 = n72178 & ~n72254;
  assign n72256 = ~n71806 & n72255;
  assign n72257 = n72253 & ~n72256;
  assign n72258 = ~P2_P2_INSTADDRPOINTER_REG_24_ & ~n70915;
  assign n72259 = P2_P2_INSTADDRPOINTER_REG_24_ & n70915;
  assign n72260 = ~n72258 & ~n72259;
  assign n72261 = n72257 & ~n72260;
  assign n72262 = ~n72257 & n72260;
  assign n72263 = ~n72261 & ~n72262;
  assign n72264 = n70085 & ~n72263;
  assign n72265 = ~n68102 & ~n72241;
  assign n72266 = n68212 & ~n72241;
  assign n72267 = n68055 & ~n72241;
  assign n72268 = ~n72266 & ~n72267;
  assign n72269 = ~P2_P2_INSTADDRPOINTER_REG_24_ & n72205;
  assign n72270 = P2_P2_INSTADDRPOINTER_REG_24_ & ~n72205;
  assign n72271 = ~n72269 & ~n72270;
  assign n72272 = n70087 & ~n72271;
  assign n72273 = n68173 & ~n72228;
  assign n72274 = n68174 & ~n72228;
  assign n72275 = n69988 & ~n72241;
  assign n72276 = n67989 & ~n72228;
  assign n72277 = n69991 & ~n72241;
  assign n72278 = ~n72276 & ~n72277;
  assign n72279 = ~n72273 & ~n72274;
  assign n72280 = ~n72275 & n72279;
  assign n72281 = n72278 & n72280;
  assign n72282 = ~n72264 & ~n72265;
  assign n72283 = n72268 & n72282;
  assign n72284 = ~n72272 & n72283;
  assign n72285 = n72281 & n72284;
  assign n72286 = n72251 & n72285;
  assign n72287 = n69980 & ~n72286;
  assign n13406 = ~n72217 | n72287;
  assign n72289 = P2_P2_INSTADDRPOINTER_REG_25_ & n69979;
  assign n72290 = P2_P2_REIP_REG_25_ & n70124;
  assign n72291 = ~n72289 & ~n72290;
  assign n72292 = P2_P2_INSTADDRPOINTER_REG_24_ & n72218;
  assign n72293 = ~P2_P2_INSTADDRPOINTER_REG_25_ & n72292;
  assign n72294 = P2_P2_INSTADDRPOINTER_REG_25_ & ~n72292;
  assign n72295 = ~n72293 & ~n72294;
  assign n72296 = n68013 & ~n72295;
  assign n72297 = n68005 & ~n72295;
  assign n72298 = ~n72296 & ~n72297;
  assign n72299 = P2_P2_INSTADDRPOINTER_REG_24_ & n72225;
  assign n72300 = ~P2_P2_INSTADDRPOINTER_REG_25_ & n72299;
  assign n72301 = P2_P2_INSTADDRPOINTER_REG_25_ & ~n72299;
  assign n72302 = ~n72300 & ~n72301;
  assign n72303 = n67915 & ~n72302;
  assign n72304 = n67993 & ~n72302;
  assign n72305 = n67997 & ~n72302;
  assign n72306 = ~n72303 & ~n72304;
  assign n72307 = ~n72305 & n72306;
  assign n72308 = P2_P2_INSTADDRPOINTER_REG_24_ & n72169;
  assign n72309 = ~P2_P2_INSTADDRPOINTER_REG_25_ & ~n72308;
  assign n72310 = P2_P2_INSTADDRPOINTER_REG_24_ & P2_P2_INSTADDRPOINTER_REG_25_;
  assign n72311 = n72169 & n72310;
  assign n72312 = ~n72309 & ~n72311;
  assign n72313 = n68016 & n72312;
  assign n72314 = P2_P2_INSTADDRPOINTER_REG_24_ & n72238;
  assign n72315 = ~P2_P2_INSTADDRPOINTER_REG_25_ & n72314;
  assign n72316 = P2_P2_INSTADDRPOINTER_REG_25_ & ~n72314;
  assign n72317 = ~n72315 & ~n72316;
  assign n72318 = n70104 & ~n72317;
  assign n72319 = ~n72313 & ~n72318;
  assign n72320 = n70093 & ~n72317;
  assign n72321 = n70097 & ~n72317;
  assign n72322 = n68059 & ~n72317;
  assign n72323 = ~n72320 & ~n72321;
  assign n72324 = ~n72322 & n72323;
  assign n72325 = n72298 & n72307;
  assign n72326 = n72319 & n72325;
  assign n72327 = n72324 & n72326;
  assign n72328 = ~P2_P2_INSTADDRPOINTER_REG_25_ & ~n70915;
  assign n72329 = P2_P2_INSTADDRPOINTER_REG_25_ & n70915;
  assign n72330 = ~n72328 & ~n72329;
  assign n72331 = P2_P2_INSTADDRPOINTER_REG_24_ & ~n70915;
  assign n72332 = ~P2_P2_INSTADDRPOINTER_REG_24_ & n70915;
  assign n72333 = ~n72257 & ~n72332;
  assign n72334 = ~n72331 & ~n72333;
  assign n72335 = ~n72330 & n72334;
  assign n72336 = ~P2_P2_INSTADDRPOINTER_REG_25_ & n70915;
  assign n72337 = P2_P2_INSTADDRPOINTER_REG_25_ & ~n70915;
  assign n72338 = ~n72336 & ~n72337;
  assign n72339 = ~n72334 & ~n72338;
  assign n72340 = ~n72335 & ~n72339;
  assign n72341 = n70085 & ~n72340;
  assign n72342 = ~n68102 & ~n72317;
  assign n72343 = P2_P2_INSTADDRPOINTER_REG_24_ & n72205;
  assign n72344 = ~P2_P2_INSTADDRPOINTER_REG_25_ & ~n72343;
  assign n72345 = n72205 & n72310;
  assign n72346 = ~n72344 & ~n72345;
  assign n72347 = n70087 & n72346;
  assign n72348 = n68212 & ~n72317;
  assign n72349 = n68055 & ~n72317;
  assign n72350 = ~n72348 & ~n72349;
  assign n72351 = n68173 & ~n72302;
  assign n72352 = n68174 & ~n72302;
  assign n72353 = n69988 & ~n72317;
  assign n72354 = n67989 & ~n72302;
  assign n72355 = n69991 & ~n72317;
  assign n72356 = ~n72354 & ~n72355;
  assign n72357 = ~n72351 & ~n72352;
  assign n72358 = ~n72353 & n72357;
  assign n72359 = n72356 & n72358;
  assign n72360 = ~n72341 & ~n72342;
  assign n72361 = ~n72347 & n72360;
  assign n72362 = n72350 & n72361;
  assign n72363 = n72359 & n72362;
  assign n72364 = n72327 & n72363;
  assign n72365 = n69980 & ~n72364;
  assign n13411 = ~n72291 | n72365;
  assign n72367 = P2_P2_INSTADDRPOINTER_REG_26_ & n69979;
  assign n72368 = P2_P2_REIP_REG_26_ & n70124;
  assign n72369 = P2_P2_INSTADDRPOINTER_REG_26_ & ~n70915;
  assign n72370 = P2_P2_INSTADDRPOINTER_REG_25_ & P2_P2_INSTADDRPOINTER_REG_26_;
  assign n72371 = n70915 & ~n72370;
  assign n72372 = ~n72369 & ~n72371;
  assign n72373 = n72334 & ~n72337;
  assign n72374 = n72372 & ~n72373;
  assign n72375 = ~P2_P2_INSTADDRPOINTER_REG_26_ & ~n70915;
  assign n72376 = P2_P2_INSTADDRPOINTER_REG_26_ & n70915;
  assign n72377 = ~n72375 & ~n72376;
  assign n72378 = ~n72337 & n72377;
  assign n72379 = ~n72334 & ~n72336;
  assign n72380 = n72378 & ~n72379;
  assign n72381 = ~n72374 & ~n72380;
  assign n72382 = n70085 & n72381;
  assign n72383 = ~P2_P2_INSTADDRPOINTER_REG_26_ & ~n72345;
  assign n72384 = P2_P2_INSTADDRPOINTER_REG_26_ & n72345;
  assign n72385 = ~n72383 & ~n72384;
  assign n72386 = n70087 & n72385;
  assign n72387 = ~n72382 & ~n72386;
  assign n72388 = P2_P2_INSTADDRPOINTER_REG_25_ & n72314;
  assign n72389 = ~P2_P2_INSTADDRPOINTER_REG_26_ & n72388;
  assign n72390 = P2_P2_INSTADDRPOINTER_REG_26_ & ~n72388;
  assign n72391 = ~n72389 & ~n72390;
  assign n72392 = ~n68102 & ~n72391;
  assign n72393 = n68212 & ~n72391;
  assign n72394 = n68055 & ~n72391;
  assign n72395 = ~n72393 & ~n72394;
  assign n72396 = P2_P2_INSTADDRPOINTER_REG_25_ & n72299;
  assign n72397 = ~P2_P2_INSTADDRPOINTER_REG_26_ & n72396;
  assign n72398 = P2_P2_INSTADDRPOINTER_REG_26_ & ~n72396;
  assign n72399 = ~n72397 & ~n72398;
  assign n72400 = n68173 & ~n72399;
  assign n72401 = n68174 & ~n72399;
  assign n72402 = n69988 & ~n72391;
  assign n72403 = n67989 & ~n72399;
  assign n72404 = n69991 & ~n72391;
  assign n72405 = ~n72403 & ~n72404;
  assign n72406 = ~n72400 & ~n72401;
  assign n72407 = ~n72402 & n72406;
  assign n72408 = n72405 & n72407;
  assign n72409 = P2_P2_INSTADDRPOINTER_REG_25_ & n72292;
  assign n72410 = ~P2_P2_INSTADDRPOINTER_REG_26_ & n72409;
  assign n72411 = P2_P2_INSTADDRPOINTER_REG_26_ & ~n72409;
  assign n72412 = ~n72410 & ~n72411;
  assign n72413 = n68013 & ~n72412;
  assign n72414 = n68005 & ~n72412;
  assign n72415 = ~n72413 & ~n72414;
  assign n72416 = n67915 & ~n72399;
  assign n72417 = n67993 & ~n72399;
  assign n72418 = n67997 & ~n72399;
  assign n72419 = ~n72416 & ~n72417;
  assign n72420 = ~n72418 & n72419;
  assign n72421 = ~P2_P2_INSTADDRPOINTER_REG_26_ & ~n72311;
  assign n72422 = P2_P2_INSTADDRPOINTER_REG_26_ & n72311;
  assign n72423 = ~n72421 & ~n72422;
  assign n72424 = n68016 & n72423;
  assign n72425 = n70104 & ~n72391;
  assign n72426 = ~n72424 & ~n72425;
  assign n72427 = n70093 & ~n72391;
  assign n72428 = n70097 & ~n72391;
  assign n72429 = n68059 & ~n72391;
  assign n72430 = ~n72427 & ~n72428;
  assign n72431 = ~n72429 & n72430;
  assign n72432 = n72415 & n72420;
  assign n72433 = n72426 & n72432;
  assign n72434 = n72431 & n72433;
  assign n72435 = n72387 & ~n72392;
  assign n72436 = n72395 & n72435;
  assign n72437 = n72408 & n72436;
  assign n72438 = n72434 & n72437;
  assign n72439 = n69980 & ~n72438;
  assign n72440 = ~n72367 & ~n72368;
  assign n13416 = n72439 | ~n72440;
  assign n72442 = P2_P2_INSTADDRPOINTER_REG_27_ & n69979;
  assign n72443 = P2_P2_REIP_REG_27_ & n70124;
  assign n72444 = ~n72337 & ~n72369;
  assign n72445 = ~n72334 & ~n72371;
  assign n72446 = n72444 & ~n72445;
  assign n72447 = ~P2_P2_INSTADDRPOINTER_REG_27_ & ~n70915;
  assign n72448 = P2_P2_INSTADDRPOINTER_REG_27_ & n70915;
  assign n72449 = ~n72447 & ~n72448;
  assign n72450 = n72446 & ~n72449;
  assign n72451 = ~n72446 & n72449;
  assign n72452 = ~n72450 & ~n72451;
  assign n72453 = n70085 & ~n72452;
  assign n72454 = ~P2_P2_INSTADDRPOINTER_REG_27_ & n72384;
  assign n72455 = P2_P2_INSTADDRPOINTER_REG_27_ & ~n72384;
  assign n72456 = ~n72454 & ~n72455;
  assign n72457 = n70087 & ~n72456;
  assign n72458 = ~n72453 & ~n72457;
  assign n72459 = P2_P2_INSTADDRPOINTER_REG_26_ & n72388;
  assign n72460 = ~P2_P2_INSTADDRPOINTER_REG_27_ & n72459;
  assign n72461 = P2_P2_INSTADDRPOINTER_REG_27_ & ~n72459;
  assign n72462 = ~n72460 & ~n72461;
  assign n72463 = ~n68102 & ~n72462;
  assign n72464 = n68212 & ~n72462;
  assign n72465 = n68055 & ~n72462;
  assign n72466 = ~n72464 & ~n72465;
  assign n72467 = P2_P2_INSTADDRPOINTER_REG_26_ & n72396;
  assign n72468 = ~P2_P2_INSTADDRPOINTER_REG_27_ & n72467;
  assign n72469 = P2_P2_INSTADDRPOINTER_REG_27_ & ~n72467;
  assign n72470 = ~n72468 & ~n72469;
  assign n72471 = n68173 & ~n72470;
  assign n72472 = n68174 & ~n72470;
  assign n72473 = n69988 & ~n72462;
  assign n72474 = n67989 & ~n72470;
  assign n72475 = n69991 & ~n72462;
  assign n72476 = ~n72474 & ~n72475;
  assign n72477 = ~n72471 & ~n72472;
  assign n72478 = ~n72473 & n72477;
  assign n72479 = n72476 & n72478;
  assign n72480 = P2_P2_INSTADDRPOINTER_REG_26_ & n72409;
  assign n72481 = ~P2_P2_INSTADDRPOINTER_REG_27_ & n72480;
  assign n72482 = P2_P2_INSTADDRPOINTER_REG_27_ & ~n72480;
  assign n72483 = ~n72481 & ~n72482;
  assign n72484 = n68013 & ~n72483;
  assign n72485 = n68005 & ~n72483;
  assign n72486 = ~n72484 & ~n72485;
  assign n72487 = n67915 & ~n72470;
  assign n72488 = n67993 & ~n72470;
  assign n72489 = n67997 & ~n72470;
  assign n72490 = ~n72487 & ~n72488;
  assign n72491 = ~n72489 & n72490;
  assign n72492 = ~P2_P2_INSTADDRPOINTER_REG_27_ & n72422;
  assign n72493 = P2_P2_INSTADDRPOINTER_REG_27_ & ~n72422;
  assign n72494 = ~n72492 & ~n72493;
  assign n72495 = n68016 & ~n72494;
  assign n72496 = n70104 & ~n72462;
  assign n72497 = ~n72495 & ~n72496;
  assign n72498 = n70093 & ~n72462;
  assign n72499 = n70097 & ~n72462;
  assign n72500 = n68059 & ~n72462;
  assign n72501 = ~n72498 & ~n72499;
  assign n72502 = ~n72500 & n72501;
  assign n72503 = n72486 & n72491;
  assign n72504 = n72497 & n72503;
  assign n72505 = n72502 & n72504;
  assign n72506 = n72458 & ~n72463;
  assign n72507 = n72466 & n72506;
  assign n72508 = n72479 & n72507;
  assign n72509 = n72505 & n72508;
  assign n72510 = n69980 & ~n72509;
  assign n72511 = ~n72442 & ~n72443;
  assign n13421 = n72510 | ~n72511;
  assign n72513 = P2_P2_INSTADDRPOINTER_REG_28_ & n69979;
  assign n72514 = P2_P2_REIP_REG_28_ & n70124;
  assign n72515 = P2_P2_INSTADDRPOINTER_REG_27_ & P2_P2_INSTADDRPOINTER_REG_28_;
  assign n72516 = ~n72446 & n72515;
  assign n72517 = n70915 & ~n72516;
  assign n72518 = P2_P2_INSTADDRPOINTER_REG_28_ & ~n70915;
  assign n72519 = ~P2_P2_INSTADDRPOINTER_REG_27_ & ~n72337;
  assign n72520 = ~n72369 & n72519;
  assign n72521 = ~n72445 & n72520;
  assign n72522 = ~n72517 & ~n72518;
  assign n72523 = ~n72521 & n72522;
  assign n72524 = P2_P2_INSTADDRPOINTER_REG_28_ & n72521;
  assign n72525 = ~n70915 & ~n72524;
  assign n72526 = P2_P2_INSTADDRPOINTER_REG_28_ & n70915;
  assign n72527 = P2_P2_INSTADDRPOINTER_REG_27_ & ~n72446;
  assign n72528 = ~n72525 & ~n72526;
  assign n72529 = ~n72527 & n72528;
  assign n72530 = ~n72523 & ~n72529;
  assign n72531 = n70085 & n72530;
  assign n72532 = P2_P2_INSTADDRPOINTER_REG_27_ & n72384;
  assign n72533 = ~P2_P2_INSTADDRPOINTER_REG_28_ & ~n72532;
  assign n72534 = n72384 & n72515;
  assign n72535 = ~n72533 & ~n72534;
  assign n72536 = n70087 & n72535;
  assign n72537 = ~n72531 & ~n72536;
  assign n72538 = P2_P2_INSTADDRPOINTER_REG_27_ & n72459;
  assign n72539 = ~P2_P2_INSTADDRPOINTER_REG_28_ & n72538;
  assign n72540 = P2_P2_INSTADDRPOINTER_REG_28_ & ~n72538;
  assign n72541 = ~n72539 & ~n72540;
  assign n72542 = ~n68102 & ~n72541;
  assign n72543 = n68212 & ~n72541;
  assign n72544 = n68055 & ~n72541;
  assign n72545 = ~n72543 & ~n72544;
  assign n72546 = P2_P2_INSTADDRPOINTER_REG_27_ & n72467;
  assign n72547 = ~P2_P2_INSTADDRPOINTER_REG_28_ & n72546;
  assign n72548 = P2_P2_INSTADDRPOINTER_REG_28_ & ~n72546;
  assign n72549 = ~n72547 & ~n72548;
  assign n72550 = n68173 & ~n72549;
  assign n72551 = n68174 & ~n72549;
  assign n72552 = n69988 & ~n72541;
  assign n72553 = n67989 & ~n72549;
  assign n72554 = n69991 & ~n72541;
  assign n72555 = ~n72553 & ~n72554;
  assign n72556 = ~n72550 & ~n72551;
  assign n72557 = ~n72552 & n72556;
  assign n72558 = n72555 & n72557;
  assign n72559 = P2_P2_INSTADDRPOINTER_REG_27_ & n72480;
  assign n72560 = ~P2_P2_INSTADDRPOINTER_REG_28_ & n72559;
  assign n72561 = P2_P2_INSTADDRPOINTER_REG_28_ & ~n72559;
  assign n72562 = ~n72560 & ~n72561;
  assign n72563 = n68013 & ~n72562;
  assign n72564 = n68005 & ~n72562;
  assign n72565 = ~n72563 & ~n72564;
  assign n72566 = n67915 & ~n72549;
  assign n72567 = n67993 & ~n72549;
  assign n72568 = n67997 & ~n72549;
  assign n72569 = ~n72566 & ~n72567;
  assign n72570 = ~n72568 & n72569;
  assign n72571 = P2_P2_INSTADDRPOINTER_REG_27_ & n72422;
  assign n72572 = ~P2_P2_INSTADDRPOINTER_REG_28_ & ~n72571;
  assign n72573 = n72422 & n72515;
  assign n72574 = ~n72572 & ~n72573;
  assign n72575 = n68016 & n72574;
  assign n72576 = n70104 & ~n72541;
  assign n72577 = ~n72575 & ~n72576;
  assign n72578 = n70093 & ~n72541;
  assign n72579 = n70097 & ~n72541;
  assign n72580 = n68059 & ~n72541;
  assign n72581 = ~n72578 & ~n72579;
  assign n72582 = ~n72580 & n72581;
  assign n72583 = n72565 & n72570;
  assign n72584 = n72577 & n72583;
  assign n72585 = n72582 & n72584;
  assign n72586 = n72537 & ~n72542;
  assign n72587 = n72545 & n72586;
  assign n72588 = n72558 & n72587;
  assign n72589 = n72585 & n72588;
  assign n72590 = n69980 & ~n72589;
  assign n72591 = ~n72513 & ~n72514;
  assign n13426 = n72590 | ~n72591;
  assign n72593 = P2_P2_INSTADDRPOINTER_REG_29_ & n69979;
  assign n72594 = P2_P2_REIP_REG_29_ & n70124;
  assign n72595 = ~n70915 & ~n72521;
  assign n72596 = ~n72518 & ~n72595;
  assign n72597 = ~n72516 & n72596;
  assign n72598 = ~P2_P2_INSTADDRPOINTER_REG_29_ & ~n70915;
  assign n72599 = P2_P2_INSTADDRPOINTER_REG_29_ & n70915;
  assign n72600 = ~n72598 & ~n72599;
  assign n72601 = n72597 & ~n72600;
  assign n72602 = ~n72597 & n72600;
  assign n72603 = ~n72601 & ~n72602;
  assign n72604 = n70085 & ~n72603;
  assign n72605 = ~P2_P2_INSTADDRPOINTER_REG_29_ & ~n72534;
  assign n72606 = P2_P2_INSTADDRPOINTER_REG_29_ & n72534;
  assign n72607 = ~n72605 & ~n72606;
  assign n72608 = n70087 & n72607;
  assign n72609 = ~n72604 & ~n72608;
  assign n72610 = P2_P2_INSTADDRPOINTER_REG_28_ & n72538;
  assign n72611 = ~P2_P2_INSTADDRPOINTER_REG_29_ & n72610;
  assign n72612 = P2_P2_INSTADDRPOINTER_REG_29_ & ~n72610;
  assign n72613 = ~n72611 & ~n72612;
  assign n72614 = ~n68102 & ~n72613;
  assign n72615 = n68212 & ~n72613;
  assign n72616 = n68055 & ~n72613;
  assign n72617 = ~n72615 & ~n72616;
  assign n72618 = P2_P2_INSTADDRPOINTER_REG_28_ & n72546;
  assign n72619 = ~P2_P2_INSTADDRPOINTER_REG_29_ & n72618;
  assign n72620 = P2_P2_INSTADDRPOINTER_REG_29_ & ~n72618;
  assign n72621 = ~n72619 & ~n72620;
  assign n72622 = n68173 & ~n72621;
  assign n72623 = n68174 & ~n72621;
  assign n72624 = n69988 & ~n72613;
  assign n72625 = n67989 & ~n72621;
  assign n72626 = n69991 & ~n72613;
  assign n72627 = ~n72625 & ~n72626;
  assign n72628 = ~n72622 & ~n72623;
  assign n72629 = ~n72624 & n72628;
  assign n72630 = n72627 & n72629;
  assign n72631 = P2_P2_INSTADDRPOINTER_REG_28_ & n72559;
  assign n72632 = ~P2_P2_INSTADDRPOINTER_REG_29_ & n72631;
  assign n72633 = P2_P2_INSTADDRPOINTER_REG_29_ & ~n72631;
  assign n72634 = ~n72632 & ~n72633;
  assign n72635 = n68013 & ~n72634;
  assign n72636 = n68005 & ~n72634;
  assign n72637 = ~n72635 & ~n72636;
  assign n72638 = n67915 & ~n72621;
  assign n72639 = n67993 & ~n72621;
  assign n72640 = n67997 & ~n72621;
  assign n72641 = ~n72638 & ~n72639;
  assign n72642 = ~n72640 & n72641;
  assign n72643 = ~P2_P2_INSTADDRPOINTER_REG_29_ & ~n72573;
  assign n72644 = P2_P2_INSTADDRPOINTER_REG_29_ & n72573;
  assign n72645 = ~n72643 & ~n72644;
  assign n72646 = n68016 & n72645;
  assign n72647 = n70104 & ~n72613;
  assign n72648 = ~n72646 & ~n72647;
  assign n72649 = n70093 & ~n72613;
  assign n72650 = n70097 & ~n72613;
  assign n72651 = n68059 & ~n72613;
  assign n72652 = ~n72649 & ~n72650;
  assign n72653 = ~n72651 & n72652;
  assign n72654 = n72637 & n72642;
  assign n72655 = n72648 & n72654;
  assign n72656 = n72653 & n72655;
  assign n72657 = n72609 & ~n72614;
  assign n72658 = n72617 & n72657;
  assign n72659 = n72630 & n72658;
  assign n72660 = n72656 & n72659;
  assign n72661 = n69980 & ~n72660;
  assign n72662 = ~n72593 & ~n72594;
  assign n13431 = n72661 | ~n72662;
  assign n72664 = P2_P2_INSTADDRPOINTER_REG_30_ & n69979;
  assign n72665 = P2_P2_REIP_REG_30_ & n70124;
  assign n72666 = ~P2_P2_INSTADDRPOINTER_REG_30_ & ~n70915;
  assign n72667 = P2_P2_INSTADDRPOINTER_REG_30_ & n70915;
  assign n72668 = ~n72666 & ~n72667;
  assign n72669 = P2_P2_INSTADDRPOINTER_REG_29_ & ~n70915;
  assign n72670 = ~P2_P2_INSTADDRPOINTER_REG_29_ & n70915;
  assign n72671 = ~n72597 & ~n72670;
  assign n72672 = ~n72669 & ~n72671;
  assign n72673 = ~n72668 & n72672;
  assign n72674 = n72668 & ~n72672;
  assign n72675 = ~n72673 & ~n72674;
  assign n72676 = n70085 & ~n72675;
  assign n72677 = ~P2_P2_INSTADDRPOINTER_REG_30_ & n72606;
  assign n72678 = P2_P2_INSTADDRPOINTER_REG_30_ & ~n72606;
  assign n72679 = ~n72677 & ~n72678;
  assign n72680 = n70087 & ~n72679;
  assign n72681 = ~n72676 & ~n72680;
  assign n72682 = P2_P2_INSTADDRPOINTER_REG_29_ & n72610;
  assign n72683 = ~P2_P2_INSTADDRPOINTER_REG_30_ & n72682;
  assign n72684 = P2_P2_INSTADDRPOINTER_REG_30_ & ~n72682;
  assign n72685 = ~n72683 & ~n72684;
  assign n72686 = ~n68102 & ~n72685;
  assign n72687 = n68212 & ~n72685;
  assign n72688 = n68055 & ~n72685;
  assign n72689 = ~n72687 & ~n72688;
  assign n72690 = P2_P2_INSTADDRPOINTER_REG_29_ & n72618;
  assign n72691 = ~P2_P2_INSTADDRPOINTER_REG_30_ & n72690;
  assign n72692 = P2_P2_INSTADDRPOINTER_REG_30_ & ~n72690;
  assign n72693 = ~n72691 & ~n72692;
  assign n72694 = n68173 & ~n72693;
  assign n72695 = n68174 & ~n72693;
  assign n72696 = n69988 & ~n72685;
  assign n72697 = n67989 & ~n72693;
  assign n72698 = n69991 & ~n72685;
  assign n72699 = ~n72697 & ~n72698;
  assign n72700 = ~n72694 & ~n72695;
  assign n72701 = ~n72696 & n72700;
  assign n72702 = n72699 & n72701;
  assign n72703 = P2_P2_INSTADDRPOINTER_REG_29_ & n72631;
  assign n72704 = ~P2_P2_INSTADDRPOINTER_REG_30_ & n72703;
  assign n72705 = P2_P2_INSTADDRPOINTER_REG_30_ & ~n72703;
  assign n72706 = ~n72704 & ~n72705;
  assign n72707 = n68013 & ~n72706;
  assign n72708 = n68005 & ~n72706;
  assign n72709 = ~n72707 & ~n72708;
  assign n72710 = n67915 & ~n72693;
  assign n72711 = n67993 & ~n72693;
  assign n72712 = n67997 & ~n72693;
  assign n72713 = ~n72710 & ~n72711;
  assign n72714 = ~n72712 & n72713;
  assign n72715 = ~P2_P2_INSTADDRPOINTER_REG_30_ & n72644;
  assign n72716 = P2_P2_INSTADDRPOINTER_REG_30_ & ~n72644;
  assign n72717 = ~n72715 & ~n72716;
  assign n72718 = n68016 & ~n72717;
  assign n72719 = n70104 & ~n72685;
  assign n72720 = ~n72718 & ~n72719;
  assign n72721 = n70093 & ~n72685;
  assign n72722 = n70097 & ~n72685;
  assign n72723 = n68059 & ~n72685;
  assign n72724 = ~n72721 & ~n72722;
  assign n72725 = ~n72723 & n72724;
  assign n72726 = n72709 & n72714;
  assign n72727 = n72720 & n72726;
  assign n72728 = n72725 & n72727;
  assign n72729 = n72681 & ~n72686;
  assign n72730 = n72689 & n72729;
  assign n72731 = n72702 & n72730;
  assign n72732 = n72728 & n72731;
  assign n72733 = n69980 & ~n72732;
  assign n72734 = ~n72664 & ~n72665;
  assign n13436 = n72733 | ~n72734;
  assign n72736 = P2_P2_INSTADDRPOINTER_REG_31_ & n69979;
  assign n72737 = P2_P2_REIP_REG_31_ & n70124;
  assign n72738 = P2_P2_INSTADDRPOINTER_REG_30_ & n72644;
  assign n72739 = ~P2_P2_INSTADDRPOINTER_REG_31_ & n72738;
  assign n72740 = P2_P2_INSTADDRPOINTER_REG_31_ & ~n72738;
  assign n72741 = ~n72739 & ~n72740;
  assign n72742 = n68016 & ~n72741;
  assign n72743 = P2_P2_INSTADDRPOINTER_REG_30_ & n72682;
  assign n72744 = ~P2_P2_INSTADDRPOINTER_REG_31_ & n72743;
  assign n72745 = P2_P2_INSTADDRPOINTER_REG_31_ & ~n72743;
  assign n72746 = ~n72744 & ~n72745;
  assign n72747 = n70104 & ~n72746;
  assign n72748 = n68059 & ~n72746;
  assign n72749 = ~n72747 & ~n72748;
  assign n72750 = P2_P2_INSTADDRPOINTER_REG_30_ & n72690;
  assign n72751 = ~P2_P2_INSTADDRPOINTER_REG_31_ & n72750;
  assign n72752 = P2_P2_INSTADDRPOINTER_REG_31_ & ~n72750;
  assign n72753 = ~n72751 & ~n72752;
  assign n72754 = n67997 & ~n72753;
  assign n72755 = n67915 & ~n72753;
  assign n72756 = P2_P2_INSTADDRPOINTER_REG_30_ & n72703;
  assign n72757 = ~P2_P2_INSTADDRPOINTER_REG_31_ & n72756;
  assign n72758 = P2_P2_INSTADDRPOINTER_REG_31_ & ~n72756;
  assign n72759 = ~n72757 & ~n72758;
  assign n72760 = n68005 & ~n72759;
  assign n72761 = ~n72754 & ~n72755;
  assign n72762 = ~n72760 & n72761;
  assign n72763 = n70093 & ~n72746;
  assign n72764 = n70097 & ~n72746;
  assign n72765 = n68013 & ~n72759;
  assign n72766 = ~n72764 & ~n72765;
  assign n72767 = n72762 & ~n72763;
  assign n72768 = n72766 & n72767;
  assign n72769 = ~n72736 & ~n72737;
  assign n72770 = ~n72742 & n72769;
  assign n72771 = n72749 & n72770;
  assign n72772 = n72768 & n72771;
  assign n72773 = P2_P2_INSTADDRPOINTER_REG_30_ & P2_P2_INSTADDRPOINTER_REG_31_;
  assign n72774 = ~n72672 & n72773;
  assign n72775 = n70915 & ~n72774;
  assign n72776 = P2_P2_INSTADDRPOINTER_REG_31_ & ~n70915;
  assign n72777 = ~P2_P2_INSTADDRPOINTER_REG_30_ & n72672;
  assign n72778 = ~n72775 & ~n72776;
  assign n72779 = ~n72777 & n72778;
  assign n72780 = ~P2_P2_INSTADDRPOINTER_REG_30_ & P2_P2_INSTADDRPOINTER_REG_31_;
  assign n72781 = ~n72669 & n72780;
  assign n72782 = ~n72671 & n72781;
  assign n72783 = ~n70915 & ~n72782;
  assign n72784 = P2_P2_INSTADDRPOINTER_REG_31_ & n70915;
  assign n72785 = P2_P2_INSTADDRPOINTER_REG_30_ & ~n72672;
  assign n72786 = ~n72783 & ~n72784;
  assign n72787 = ~n72785 & n72786;
  assign n72788 = ~n72779 & ~n72787;
  assign n72789 = n70085 & n72788;
  assign n72790 = P2_P2_INSTADDRPOINTER_REG_30_ & n72606;
  assign n72791 = ~P2_P2_INSTADDRPOINTER_REG_31_ & n72790;
  assign n72792 = P2_P2_INSTADDRPOINTER_REG_31_ & ~n72790;
  assign n72793 = ~n72791 & ~n72792;
  assign n72794 = n70087 & ~n72793;
  assign n72795 = ~n72789 & ~n72794;
  assign n72796 = ~n68102 & ~n72746;
  assign n72797 = n68212 & ~n72746;
  assign n72798 = n68055 & ~n72746;
  assign n72799 = ~n72797 & ~n72798;
  assign n72800 = n68174 & ~n72753;
  assign n72801 = n72799 & ~n72800;
  assign n72802 = n69988 & ~n72746;
  assign n72803 = n68173 & ~n72753;
  assign n72804 = n67993 & ~n72753;
  assign n72805 = n67989 & ~n72753;
  assign n72806 = n69991 & ~n72746;
  assign n72807 = ~n72804 & ~n72805;
  assign n72808 = ~n72806 & n72807;
  assign n72809 = ~n72802 & ~n72803;
  assign n72810 = n72808 & n72809;
  assign n72811 = n72795 & ~n72796;
  assign n72812 = n72801 & n72811;
  assign n72813 = n72810 & n72812;
  assign n72814 = n72772 & n72813;
  assign n72815 = ~n69980 & ~n72736;
  assign n72816 = ~n72737 & n72815;
  assign n13441 = ~n72814 & ~n72816;
  assign n72818 = P2_P2_STATE2_REG_0_ & ~n67882;
  assign n72819 = ~P2_P2_STATE2_REG_0_ & ~n69947;
  assign n72820 = n68016 & n68019;
  assign n72821 = n68021 & n68025;
  assign n72822 = ~n72820 & ~n72821;
  assign n72823 = n68268 & ~n72822;
  assign n72824 = ~n72819 & ~n72823;
  assign n72825 = n72818 & ~n72824;
  assign n72826 = ~n70084 & n72825;
  assign n72827 = ~n70053 & n72826;
  assign n72828 = n70084 & n72825;
  assign n72829 = ~n70053 & n72828;
  assign n72830 = P2_P2_STATE2_REG_1_ & ~n72824;
  assign n72831 = P2_P2_STATEBS16_REG & n72830;
  assign n72832 = P2_P2_PHYADDRPOINTER_REG_0_ & n72831;
  assign n72833 = ~P2_P2_STATEBS16_REG & n72830;
  assign n72834 = P2_P2_PHYADDRPOINTER_REG_0_ & n72833;
  assign n72835 = P2_P2_PHYADDRPOINTER_REG_0_ & n72824;
  assign n72836 = P2_P2_STATE2_REG_0_ & n67882;
  assign n72837 = ~n72824 & n72836;
  assign n72838 = ~n70101 & n72837;
  assign n72839 = P2_P2_STATE2_REG_2_ & ~P2_P2_STATE2_REG_0_;
  assign n72840 = ~n72824 & n72839;
  assign n72841 = P2_P2_PHYADDRPOINTER_REG_0_ & n72840;
  assign n72842 = n68284 & ~n72824;
  assign n72843 = P2_P2_REIP_REG_0_ & n72842;
  assign n72844 = ~n72835 & ~n72838;
  assign n72845 = ~n72841 & n72844;
  assign n72846 = ~n72843 & n72845;
  assign n72847 = ~n72827 & ~n72829;
  assign n72848 = ~n72832 & n72847;
  assign n72849 = ~n72834 & n72848;
  assign n13446 = ~n72846 | ~n72849;
  assign n72851 = ~n70225 & n72826;
  assign n72852 = ~n70175 & n72828;
  assign n72853 = P2_P2_PHYADDRPOINTER_REG_1_ & n72831;
  assign n72854 = ~P2_P2_PHYADDRPOINTER_REG_1_ & n72833;
  assign n72855 = P2_P2_PHYADDRPOINTER_REG_1_ & n72824;
  assign n72856 = ~n70205 & n72837;
  assign n72857 = ~P2_P2_PHYADDRPOINTER_REG_1_ & n72840;
  assign n72858 = P2_P2_REIP_REG_1_ & n72842;
  assign n72859 = ~n72855 & ~n72856;
  assign n72860 = ~n72857 & n72859;
  assign n72861 = ~n72858 & n72860;
  assign n72862 = ~n72851 & ~n72852;
  assign n72863 = ~n72853 & n72862;
  assign n72864 = ~n72854 & n72863;
  assign n13451 = ~n72861 | ~n72864;
  assign n72866 = ~n70310 & n72826;
  assign n72867 = ~n70297 & n72828;
  assign n72868 = ~P2_P2_PHYADDRPOINTER_REG_2_ & n72831;
  assign n72869 = P2_P2_PHYADDRPOINTER_REG_1_ & ~P2_P2_PHYADDRPOINTER_REG_2_;
  assign n72870 = ~P2_P2_PHYADDRPOINTER_REG_1_ & P2_P2_PHYADDRPOINTER_REG_2_;
  assign n72871 = ~n72869 & ~n72870;
  assign n72872 = n72833 & ~n72871;
  assign n72873 = n72840 & ~n72871;
  assign n72874 = P2_P2_REIP_REG_2_ & n72842;
  assign n72875 = P2_P2_PHYADDRPOINTER_REG_2_ & n72824;
  assign n72876 = ~n70347 & n72837;
  assign n72877 = ~n72873 & ~n72874;
  assign n72878 = ~n72875 & n72877;
  assign n72879 = ~n72876 & n72878;
  assign n72880 = ~n72866 & ~n72867;
  assign n72881 = ~n72868 & n72880;
  assign n72882 = ~n72872 & n72881;
  assign n13456 = ~n72879 | ~n72882;
  assign n72884 = ~n70425 & n72826;
  assign n72885 = n70440 & n72828;
  assign n72886 = P2_P2_PHYADDRPOINTER_REG_2_ & ~P2_P2_PHYADDRPOINTER_REG_3_;
  assign n72887 = ~P2_P2_PHYADDRPOINTER_REG_2_ & P2_P2_PHYADDRPOINTER_REG_3_;
  assign n72888 = ~n72886 & ~n72887;
  assign n72889 = n72831 & ~n72888;
  assign n72890 = P2_P2_PHYADDRPOINTER_REG_1_ & P2_P2_PHYADDRPOINTER_REG_2_;
  assign n72891 = ~P2_P2_PHYADDRPOINTER_REG_3_ & n72890;
  assign n72892 = P2_P2_PHYADDRPOINTER_REG_3_ & ~n72890;
  assign n72893 = ~n72891 & ~n72892;
  assign n72894 = n72833 & ~n72893;
  assign n72895 = n72840 & ~n72893;
  assign n72896 = P2_P2_REIP_REG_3_ & n72842;
  assign n72897 = P2_P2_PHYADDRPOINTER_REG_3_ & n72824;
  assign n72898 = n70478 & n72837;
  assign n72899 = ~n72895 & ~n72896;
  assign n72900 = ~n72897 & n72899;
  assign n72901 = ~n72898 & n72900;
  assign n72902 = ~n72884 & ~n72885;
  assign n72903 = ~n72889 & n72902;
  assign n72904 = ~n72894 & n72903;
  assign n13461 = ~n72901 | ~n72904;
  assign n72906 = P2_P2_PHYADDRPOINTER_REG_2_ & P2_P2_PHYADDRPOINTER_REG_3_;
  assign n72907 = ~P2_P2_PHYADDRPOINTER_REG_4_ & n72906;
  assign n72908 = P2_P2_PHYADDRPOINTER_REG_4_ & ~n72906;
  assign n72909 = ~n72907 & ~n72908;
  assign n72910 = n72831 & ~n72909;
  assign n72911 = P2_P2_PHYADDRPOINTER_REG_3_ & n72890;
  assign n72912 = ~P2_P2_PHYADDRPOINTER_REG_4_ & n72911;
  assign n72913 = P2_P2_PHYADDRPOINTER_REG_4_ & ~n72911;
  assign n72914 = ~n72912 & ~n72913;
  assign n72915 = n72833 & ~n72914;
  assign n72916 = n70553 & n72828;
  assign n72917 = ~n70575 & n72826;
  assign n72918 = n72840 & ~n72914;
  assign n72919 = P2_P2_REIP_REG_4_ & n72842;
  assign n72920 = P2_P2_PHYADDRPOINTER_REG_4_ & n72824;
  assign n72921 = ~n70614 & n72837;
  assign n72922 = ~n72918 & ~n72919;
  assign n72923 = ~n72920 & n72922;
  assign n72924 = ~n72921 & n72923;
  assign n72925 = ~n72910 & ~n72915;
  assign n72926 = ~n72916 & n72925;
  assign n72927 = ~n72917 & n72926;
  assign n13466 = ~n72924 | ~n72927;
  assign n72929 = P2_P2_PHYADDRPOINTER_REG_4_ & n72906;
  assign n72930 = ~P2_P2_PHYADDRPOINTER_REG_5_ & n72929;
  assign n72931 = P2_P2_PHYADDRPOINTER_REG_5_ & ~n72929;
  assign n72932 = ~n72930 & ~n72931;
  assign n72933 = n72831 & ~n72932;
  assign n72934 = P2_P2_PHYADDRPOINTER_REG_4_ & n72911;
  assign n72935 = ~P2_P2_PHYADDRPOINTER_REG_5_ & n72934;
  assign n72936 = P2_P2_PHYADDRPOINTER_REG_5_ & ~n72934;
  assign n72937 = ~n72935 & ~n72936;
  assign n72938 = n72833 & ~n72937;
  assign n72939 = ~n70690 & n72826;
  assign n72940 = ~n70708 & n72828;
  assign n72941 = n72840 & ~n72937;
  assign n72942 = P2_P2_REIP_REG_5_ & n72842;
  assign n72943 = P2_P2_PHYADDRPOINTER_REG_5_ & n72824;
  assign n72944 = n70747 & n72837;
  assign n72945 = ~n72941 & ~n72942;
  assign n72946 = ~n72943 & n72945;
  assign n72947 = ~n72944 & n72946;
  assign n72948 = ~n72933 & ~n72938;
  assign n72949 = ~n72939 & n72948;
  assign n72950 = ~n72940 & n72949;
  assign n13471 = ~n72947 | ~n72950;
  assign n72952 = P2_P2_PHYADDRPOINTER_REG_5_ & n72929;
  assign n72953 = ~P2_P2_PHYADDRPOINTER_REG_6_ & n72952;
  assign n72954 = P2_P2_PHYADDRPOINTER_REG_6_ & ~n72952;
  assign n72955 = ~n72953 & ~n72954;
  assign n72956 = n72831 & ~n72955;
  assign n72957 = P2_P2_PHYADDRPOINTER_REG_5_ & n72934;
  assign n72958 = ~P2_P2_PHYADDRPOINTER_REG_6_ & n72957;
  assign n72959 = P2_P2_PHYADDRPOINTER_REG_6_ & ~n72957;
  assign n72960 = ~n72958 & ~n72959;
  assign n72961 = n72833 & ~n72960;
  assign n72962 = ~n70821 & n72826;
  assign n72963 = ~n70840 & n72828;
  assign n72964 = n72840 & ~n72960;
  assign n72965 = P2_P2_REIP_REG_6_ & n72842;
  assign n72966 = P2_P2_PHYADDRPOINTER_REG_6_ & n72824;
  assign n72967 = ~n70878 & n72837;
  assign n72968 = ~n72964 & ~n72965;
  assign n72969 = ~n72966 & n72968;
  assign n72970 = ~n72967 & n72969;
  assign n72971 = ~n72956 & ~n72961;
  assign n72972 = ~n72962 & n72971;
  assign n72973 = ~n72963 & n72972;
  assign n13476 = ~n72970 | ~n72973;
  assign n72975 = P2_P2_PHYADDRPOINTER_REG_6_ & n72952;
  assign n72976 = ~P2_P2_PHYADDRPOINTER_REG_7_ & n72975;
  assign n72977 = P2_P2_PHYADDRPOINTER_REG_7_ & ~n72975;
  assign n72978 = ~n72976 & ~n72977;
  assign n72979 = n72831 & ~n72978;
  assign n72980 = P2_P2_PHYADDRPOINTER_REG_6_ & n72957;
  assign n72981 = ~P2_P2_PHYADDRPOINTER_REG_7_ & n72980;
  assign n72982 = P2_P2_PHYADDRPOINTER_REG_7_ & ~n72980;
  assign n72983 = ~n72981 & ~n72982;
  assign n72984 = n72833 & ~n72983;
  assign n72985 = ~n70922 & n72826;
  assign n72986 = ~n70940 & n72828;
  assign n72987 = n72840 & ~n72983;
  assign n72988 = P2_P2_REIP_REG_7_ & n72842;
  assign n72989 = P2_P2_PHYADDRPOINTER_REG_7_ & n72824;
  assign n72990 = ~n70976 & n72837;
  assign n72991 = ~n72987 & ~n72988;
  assign n72992 = ~n72989 & n72991;
  assign n72993 = ~n72990 & n72992;
  assign n72994 = ~n72979 & ~n72984;
  assign n72995 = ~n72985 & n72994;
  assign n72996 = ~n72986 & n72995;
  assign n13481 = ~n72993 | ~n72996;
  assign n72998 = P2_P2_PHYADDRPOINTER_REG_7_ & n72975;
  assign n72999 = ~P2_P2_PHYADDRPOINTER_REG_8_ & n72998;
  assign n73000 = P2_P2_PHYADDRPOINTER_REG_8_ & ~n72998;
  assign n73001 = ~n72999 & ~n73000;
  assign n73002 = n72831 & ~n73001;
  assign n73003 = P2_P2_PHYADDRPOINTER_REG_7_ & n72980;
  assign n73004 = ~P2_P2_PHYADDRPOINTER_REG_8_ & n73003;
  assign n73005 = P2_P2_PHYADDRPOINTER_REG_8_ & ~n73003;
  assign n73006 = ~n73004 & ~n73005;
  assign n73007 = n72833 & ~n73006;
  assign n73008 = ~n71016 & n72826;
  assign n73009 = ~n71032 & n72828;
  assign n73010 = n72840 & ~n73006;
  assign n73011 = P2_P2_REIP_REG_8_ & n72842;
  assign n73012 = P2_P2_PHYADDRPOINTER_REG_8_ & n72824;
  assign n73013 = ~n71066 & n72837;
  assign n73014 = ~n73010 & ~n73011;
  assign n73015 = ~n73012 & n73014;
  assign n73016 = ~n73013 & n73015;
  assign n73017 = ~n73002 & ~n73007;
  assign n73018 = ~n73008 & n73017;
  assign n73019 = ~n73009 & n73018;
  assign n13486 = ~n73016 | ~n73019;
  assign n73021 = P2_P2_PHYADDRPOINTER_REG_8_ & n72998;
  assign n73022 = ~P2_P2_PHYADDRPOINTER_REG_9_ & n73021;
  assign n73023 = P2_P2_PHYADDRPOINTER_REG_9_ & ~n73021;
  assign n73024 = ~n73022 & ~n73023;
  assign n73025 = n72831 & ~n73024;
  assign n73026 = P2_P2_PHYADDRPOINTER_REG_8_ & n73003;
  assign n73027 = ~P2_P2_PHYADDRPOINTER_REG_9_ & n73026;
  assign n73028 = P2_P2_PHYADDRPOINTER_REG_9_ & ~n73026;
  assign n73029 = ~n73027 & ~n73028;
  assign n73030 = n72833 & ~n73029;
  assign n73031 = ~n71109 & n72826;
  assign n73032 = n71120 & n72828;
  assign n73033 = n72840 & ~n73029;
  assign n73034 = P2_P2_REIP_REG_9_ & n72842;
  assign n73035 = P2_P2_PHYADDRPOINTER_REG_9_ & n72824;
  assign n73036 = n71149 & n72837;
  assign n73037 = ~n73033 & ~n73034;
  assign n73038 = ~n73035 & n73037;
  assign n73039 = ~n73036 & n73038;
  assign n73040 = ~n73025 & ~n73030;
  assign n73041 = ~n73031 & n73040;
  assign n73042 = ~n73032 & n73041;
  assign n13491 = ~n73039 | ~n73042;
  assign n73044 = P2_P2_PHYADDRPOINTER_REG_9_ & n73021;
  assign n73045 = ~P2_P2_PHYADDRPOINTER_REG_10_ & n73044;
  assign n73046 = P2_P2_PHYADDRPOINTER_REG_10_ & ~n73044;
  assign n73047 = ~n73045 & ~n73046;
  assign n73048 = n72831 & ~n73047;
  assign n73049 = P2_P2_PHYADDRPOINTER_REG_9_ & n73026;
  assign n73050 = ~P2_P2_PHYADDRPOINTER_REG_10_ & n73049;
  assign n73051 = P2_P2_PHYADDRPOINTER_REG_10_ & ~n73049;
  assign n73052 = ~n73050 & ~n73051;
  assign n73053 = n72833 & ~n73052;
  assign n73054 = ~n71192 & n72826;
  assign n73055 = n71200 & n72828;
  assign n73056 = n72840 & ~n73052;
  assign n73057 = P2_P2_REIP_REG_10_ & n72842;
  assign n73058 = P2_P2_PHYADDRPOINTER_REG_10_ & n72824;
  assign n73059 = n71225 & n72837;
  assign n73060 = ~n73056 & ~n73057;
  assign n73061 = ~n73058 & n73060;
  assign n73062 = ~n73059 & n73061;
  assign n73063 = ~n73048 & ~n73053;
  assign n73064 = ~n73054 & n73063;
  assign n73065 = ~n73055 & n73064;
  assign n13496 = ~n73062 | ~n73065;
  assign n73067 = P2_P2_PHYADDRPOINTER_REG_10_ & n73044;
  assign n73068 = ~P2_P2_PHYADDRPOINTER_REG_11_ & n73067;
  assign n73069 = P2_P2_PHYADDRPOINTER_REG_11_ & ~n73067;
  assign n73070 = ~n73068 & ~n73069;
  assign n73071 = n72831 & ~n73070;
  assign n73072 = P2_P2_PHYADDRPOINTER_REG_10_ & n73049;
  assign n73073 = ~P2_P2_PHYADDRPOINTER_REG_11_ & n73072;
  assign n73074 = P2_P2_PHYADDRPOINTER_REG_11_ & ~n73072;
  assign n73075 = ~n73073 & ~n73074;
  assign n73076 = n72833 & ~n73075;
  assign n73077 = ~n71286 & n72826;
  assign n73078 = ~n71299 & n72828;
  assign n73079 = n72840 & ~n73075;
  assign n73080 = P2_P2_REIP_REG_11_ & n72842;
  assign n73081 = P2_P2_PHYADDRPOINTER_REG_11_ & n72824;
  assign n73082 = ~n71269 & n72837;
  assign n73083 = ~n73079 & ~n73080;
  assign n73084 = ~n73081 & n73083;
  assign n73085 = ~n73082 & n73084;
  assign n73086 = ~n73071 & ~n73076;
  assign n73087 = ~n73077 & n73086;
  assign n73088 = ~n73078 & n73087;
  assign n13501 = ~n73085 | ~n73088;
  assign n73090 = P2_P2_PHYADDRPOINTER_REG_11_ & n73067;
  assign n73091 = ~P2_P2_PHYADDRPOINTER_REG_12_ & n73090;
  assign n73092 = P2_P2_PHYADDRPOINTER_REG_12_ & ~n73090;
  assign n73093 = ~n73091 & ~n73092;
  assign n73094 = n72831 & ~n73093;
  assign n73095 = P2_P2_PHYADDRPOINTER_REG_11_ & n73072;
  assign n73096 = ~P2_P2_PHYADDRPOINTER_REG_12_ & n73095;
  assign n73097 = P2_P2_PHYADDRPOINTER_REG_12_ & ~n73095;
  assign n73098 = ~n73096 & ~n73097;
  assign n73099 = n72833 & ~n73098;
  assign n73100 = ~n71340 & n72826;
  assign n73101 = n71349 & n72828;
  assign n73102 = P2_P2_PHYADDRPOINTER_REG_12_ & n72824;
  assign n73103 = P2_P2_REIP_REG_12_ & n72842;
  assign n73104 = n72840 & ~n73098;
  assign n73105 = n71375 & n72837;
  assign n73106 = ~n73102 & ~n73103;
  assign n73107 = ~n73104 & n73106;
  assign n73108 = ~n73105 & n73107;
  assign n73109 = ~n73094 & ~n73099;
  assign n73110 = ~n73100 & n73109;
  assign n73111 = ~n73101 & n73110;
  assign n13506 = ~n73108 | ~n73111;
  assign n73113 = P2_P2_PHYADDRPOINTER_REG_12_ & n73090;
  assign n73114 = ~P2_P2_PHYADDRPOINTER_REG_13_ & n73113;
  assign n73115 = P2_P2_PHYADDRPOINTER_REG_13_ & ~n73113;
  assign n73116 = ~n73114 & ~n73115;
  assign n73117 = n72831 & ~n73116;
  assign n73118 = P2_P2_PHYADDRPOINTER_REG_12_ & n73095;
  assign n73119 = ~P2_P2_PHYADDRPOINTER_REG_13_ & n73118;
  assign n73120 = P2_P2_PHYADDRPOINTER_REG_13_ & ~n73118;
  assign n73121 = ~n73119 & ~n73120;
  assign n73122 = n72833 & ~n73121;
  assign n73123 = n71418 & n72826;
  assign n73124 = n71425 & n72828;
  assign n73125 = P2_P2_PHYADDRPOINTER_REG_13_ & n72824;
  assign n73126 = P2_P2_REIP_REG_13_ & n72842;
  assign n73127 = n72840 & ~n73121;
  assign n73128 = n71450 & n72837;
  assign n73129 = ~n73125 & ~n73126;
  assign n73130 = ~n73127 & n73129;
  assign n73131 = ~n73128 & n73130;
  assign n73132 = ~n73117 & ~n73122;
  assign n73133 = ~n73123 & n73132;
  assign n73134 = ~n73124 & n73133;
  assign n13511 = ~n73131 | ~n73134;
  assign n73136 = P2_P2_PHYADDRPOINTER_REG_13_ & n73113;
  assign n73137 = ~P2_P2_PHYADDRPOINTER_REG_14_ & n73136;
  assign n73138 = P2_P2_PHYADDRPOINTER_REG_14_ & ~n73136;
  assign n73139 = ~n73137 & ~n73138;
  assign n73140 = n72831 & ~n73139;
  assign n73141 = P2_P2_PHYADDRPOINTER_REG_13_ & n73118;
  assign n73142 = ~P2_P2_PHYADDRPOINTER_REG_14_ & n73141;
  assign n73143 = P2_P2_PHYADDRPOINTER_REG_14_ & ~n73141;
  assign n73144 = ~n73142 & ~n73143;
  assign n73145 = n72833 & ~n73144;
  assign n73146 = ~n71521 & n72826;
  assign n73147 = ~n71525 & n72828;
  assign n73148 = P2_P2_PHYADDRPOINTER_REG_14_ & n72824;
  assign n73149 = P2_P2_REIP_REG_14_ & n72842;
  assign n73150 = n72840 & ~n73144;
  assign n73151 = ~n71494 & n72837;
  assign n73152 = ~n73148 & ~n73149;
  assign n73153 = ~n73150 & n73152;
  assign n73154 = ~n73151 & n73153;
  assign n73155 = ~n73140 & ~n73145;
  assign n73156 = ~n73146 & n73155;
  assign n73157 = ~n73147 & n73156;
  assign n13516 = ~n73154 | ~n73157;
  assign n73159 = P2_P2_PHYADDRPOINTER_REG_14_ & n73136;
  assign n73160 = ~P2_P2_PHYADDRPOINTER_REG_15_ & n73159;
  assign n73161 = P2_P2_PHYADDRPOINTER_REG_15_ & ~n73159;
  assign n73162 = ~n73160 & ~n73161;
  assign n73163 = n72831 & ~n73162;
  assign n73164 = P2_P2_PHYADDRPOINTER_REG_14_ & n73141;
  assign n73165 = ~P2_P2_PHYADDRPOINTER_REG_15_ & n73164;
  assign n73166 = P2_P2_PHYADDRPOINTER_REG_15_ & ~n73164;
  assign n73167 = ~n73165 & ~n73166;
  assign n73168 = n72833 & ~n73167;
  assign n73169 = ~n71598 & n72826;
  assign n73170 = n71603 & n72828;
  assign n73171 = P2_P2_PHYADDRPOINTER_REG_15_ & n72824;
  assign n73172 = P2_P2_REIP_REG_15_ & n72842;
  assign n73173 = n72840 & ~n73167;
  assign n73174 = n71570 & n72837;
  assign n73175 = ~n73171 & ~n73172;
  assign n73176 = ~n73173 & n73175;
  assign n73177 = ~n73174 & n73176;
  assign n73178 = ~n73163 & ~n73168;
  assign n73179 = ~n73169 & n73178;
  assign n73180 = ~n73170 & n73179;
  assign n13521 = ~n73177 | ~n73180;
  assign n73182 = P2_P2_PHYADDRPOINTER_REG_15_ & n73159;
  assign n73183 = ~P2_P2_PHYADDRPOINTER_REG_16_ & n73182;
  assign n73184 = P2_P2_PHYADDRPOINTER_REG_16_ & ~n73182;
  assign n73185 = ~n73183 & ~n73184;
  assign n73186 = n72831 & ~n73185;
  assign n73187 = P2_P2_PHYADDRPOINTER_REG_15_ & n73164;
  assign n73188 = ~P2_P2_PHYADDRPOINTER_REG_16_ & n73187;
  assign n73189 = P2_P2_PHYADDRPOINTER_REG_16_ & ~n73187;
  assign n73190 = ~n73188 & ~n73189;
  assign n73191 = n72833 & ~n73190;
  assign n73192 = ~n71662 & n72826;
  assign n73193 = ~n71675 & n72828;
  assign n73194 = P2_P2_PHYADDRPOINTER_REG_16_ & n72824;
  assign n73195 = P2_P2_REIP_REG_16_ & n72842;
  assign n73196 = n72840 & ~n73190;
  assign n73197 = ~n71645 & n72837;
  assign n73198 = ~n73194 & ~n73195;
  assign n73199 = ~n73196 & n73198;
  assign n73200 = ~n73197 & n73199;
  assign n73201 = ~n73186 & ~n73191;
  assign n73202 = ~n73192 & n73201;
  assign n73203 = ~n73193 & n73202;
  assign n13526 = ~n73200 | ~n73203;
  assign n73205 = P2_P2_PHYADDRPOINTER_REG_16_ & n73182;
  assign n73206 = ~P2_P2_PHYADDRPOINTER_REG_17_ & n73205;
  assign n73207 = P2_P2_PHYADDRPOINTER_REG_17_ & ~n73205;
  assign n73208 = ~n73206 & ~n73207;
  assign n73209 = n72831 & ~n73208;
  assign n73210 = P2_P2_PHYADDRPOINTER_REG_16_ & n73187;
  assign n73211 = ~P2_P2_PHYADDRPOINTER_REG_17_ & n73210;
  assign n73212 = P2_P2_PHYADDRPOINTER_REG_17_ & ~n73210;
  assign n73213 = ~n73211 & ~n73212;
  assign n73214 = n72833 & ~n73213;
  assign n73215 = n71718 & n72826;
  assign n73216 = n71726 & n72828;
  assign n73217 = P2_P2_PHYADDRPOINTER_REG_17_ & n72824;
  assign n73218 = P2_P2_REIP_REG_17_ & n72842;
  assign n73219 = n72840 & ~n73213;
  assign n73220 = n71752 & n72837;
  assign n73221 = ~n73217 & ~n73218;
  assign n73222 = ~n73219 & n73221;
  assign n73223 = ~n73220 & n73222;
  assign n73224 = ~n73209 & ~n73214;
  assign n73225 = ~n73215 & n73224;
  assign n73226 = ~n73216 & n73225;
  assign n13531 = ~n73223 | ~n73226;
  assign n73228 = P2_P2_PHYADDRPOINTER_REG_17_ & n73205;
  assign n73229 = ~P2_P2_PHYADDRPOINTER_REG_18_ & n73228;
  assign n73230 = P2_P2_PHYADDRPOINTER_REG_18_ & ~n73228;
  assign n73231 = ~n73229 & ~n73230;
  assign n73232 = n72831 & ~n73231;
  assign n73233 = P2_P2_PHYADDRPOINTER_REG_17_ & n73210;
  assign n73234 = ~P2_P2_PHYADDRPOINTER_REG_18_ & n73233;
  assign n73235 = P2_P2_PHYADDRPOINTER_REG_18_ & ~n73233;
  assign n73236 = ~n73234 & ~n73235;
  assign n73237 = n72833 & ~n73236;
  assign n73238 = ~n71812 & n72826;
  assign n73239 = ~n71825 & n72828;
  assign n73240 = P2_P2_PHYADDRPOINTER_REG_18_ & n72824;
  assign n73241 = P2_P2_REIP_REG_18_ & n72842;
  assign n73242 = n72840 & ~n73236;
  assign n73243 = ~n71796 & n72837;
  assign n73244 = ~n73240 & ~n73241;
  assign n73245 = ~n73242 & n73244;
  assign n73246 = ~n73243 & n73245;
  assign n73247 = ~n73232 & ~n73237;
  assign n73248 = ~n73238 & n73247;
  assign n73249 = ~n73239 & n73248;
  assign n13536 = ~n73246 | ~n73249;
  assign n73251 = P2_P2_PHYADDRPOINTER_REG_18_ & n73228;
  assign n73252 = ~P2_P2_PHYADDRPOINTER_REG_19_ & n73251;
  assign n73253 = P2_P2_PHYADDRPOINTER_REG_19_ & ~n73251;
  assign n73254 = ~n73252 & ~n73253;
  assign n73255 = n72831 & ~n73254;
  assign n73256 = P2_P2_PHYADDRPOINTER_REG_18_ & n73233;
  assign n73257 = ~P2_P2_PHYADDRPOINTER_REG_19_ & n73256;
  assign n73258 = P2_P2_PHYADDRPOINTER_REG_19_ & ~n73256;
  assign n73259 = ~n73257 & ~n73258;
  assign n73260 = n72833 & ~n73259;
  assign n73261 = ~n71866 & n72826;
  assign n73262 = n71875 & n72828;
  assign n73263 = P2_P2_PHYADDRPOINTER_REG_19_ & n72824;
  assign n73264 = P2_P2_REIP_REG_19_ & n72842;
  assign n73265 = n72840 & ~n73259;
  assign n73266 = n71901 & n72837;
  assign n73267 = ~n73263 & ~n73264;
  assign n73268 = ~n73265 & n73267;
  assign n73269 = ~n73266 & n73268;
  assign n73270 = ~n73255 & ~n73260;
  assign n73271 = ~n73261 & n73270;
  assign n73272 = ~n73262 & n73271;
  assign n13541 = ~n73269 | ~n73272;
  assign n73274 = P2_P2_PHYADDRPOINTER_REG_19_ & n73251;
  assign n73275 = ~P2_P2_PHYADDRPOINTER_REG_20_ & n73274;
  assign n73276 = P2_P2_PHYADDRPOINTER_REG_20_ & ~n73274;
  assign n73277 = ~n73275 & ~n73276;
  assign n73278 = n72831 & ~n73277;
  assign n73279 = P2_P2_PHYADDRPOINTER_REG_19_ & n73256;
  assign n73280 = ~P2_P2_PHYADDRPOINTER_REG_20_ & n73279;
  assign n73281 = P2_P2_PHYADDRPOINTER_REG_20_ & ~n73279;
  assign n73282 = ~n73280 & ~n73281;
  assign n73283 = n72833 & ~n73282;
  assign n73284 = n71953 & n72828;
  assign n73285 = P2_P2_PHYADDRPOINTER_REG_20_ & n72824;
  assign n73286 = P2_P2_REIP_REG_20_ & n72842;
  assign n73287 = n72840 & ~n73282;
  assign n73288 = n71977 & n72837;
  assign n73289 = ~n73285 & ~n73286;
  assign n73290 = ~n73287 & n73289;
  assign n73291 = ~n73288 & n73290;
  assign n73292 = n71928 & n72826;
  assign n73293 = ~n73278 & ~n73283;
  assign n73294 = ~n73284 & n73293;
  assign n73295 = n73291 & n73294;
  assign n13546 = n73292 | ~n73295;
  assign n73297 = P2_P2_PHYADDRPOINTER_REG_20_ & n73274;
  assign n73298 = ~P2_P2_PHYADDRPOINTER_REG_21_ & n73297;
  assign n73299 = P2_P2_PHYADDRPOINTER_REG_21_ & ~n73297;
  assign n73300 = ~n73298 & ~n73299;
  assign n73301 = n72831 & ~n73300;
  assign n73302 = P2_P2_PHYADDRPOINTER_REG_20_ & n73279;
  assign n73303 = ~P2_P2_PHYADDRPOINTER_REG_21_ & n73302;
  assign n73304 = P2_P2_PHYADDRPOINTER_REG_21_ & ~n73302;
  assign n73305 = ~n73303 & ~n73304;
  assign n73306 = n72833 & ~n73305;
  assign n73307 = n72010 & n72828;
  assign n73308 = P2_P2_PHYADDRPOINTER_REG_21_ & n72824;
  assign n73309 = P2_P2_REIP_REG_21_ & n72842;
  assign n73310 = n72840 & ~n73305;
  assign n73311 = n72035 & n72837;
  assign n73312 = ~n73308 & ~n73309;
  assign n73313 = ~n73310 & n73312;
  assign n73314 = ~n73311 & n73313;
  assign n73315 = ~n72051 & n72826;
  assign n73316 = ~n73301 & ~n73306;
  assign n73317 = ~n73307 & n73316;
  assign n73318 = n73314 & n73317;
  assign n13551 = n73315 | ~n73318;
  assign n73320 = P2_P2_PHYADDRPOINTER_REG_21_ & n73297;
  assign n73321 = ~P2_P2_PHYADDRPOINTER_REG_22_ & n73320;
  assign n73322 = P2_P2_PHYADDRPOINTER_REG_22_ & ~n73320;
  assign n73323 = ~n73321 & ~n73322;
  assign n73324 = n72831 & ~n73323;
  assign n73325 = ~n72112 & n72826;
  assign n73326 = P2_P2_PHYADDRPOINTER_REG_21_ & n73302;
  assign n73327 = ~P2_P2_PHYADDRPOINTER_REG_22_ & n73326;
  assign n73328 = P2_P2_PHYADDRPOINTER_REG_22_ & ~n73326;
  assign n73329 = ~n73327 & ~n73328;
  assign n73330 = n72833 & ~n73329;
  assign n73331 = ~n72129 & n72828;
  assign n73332 = P2_P2_PHYADDRPOINTER_REG_22_ & n72824;
  assign n73333 = P2_P2_REIP_REG_22_ & n72842;
  assign n73334 = n72840 & ~n73329;
  assign n73335 = ~n72091 & n72837;
  assign n73336 = ~n73332 & ~n73333;
  assign n73337 = ~n73334 & n73336;
  assign n73338 = ~n73335 & n73337;
  assign n73339 = ~n73324 & ~n73325;
  assign n73340 = ~n73330 & n73339;
  assign n73341 = ~n73331 & n73340;
  assign n13556 = ~n73338 | ~n73341;
  assign n73343 = P2_P2_PHYADDRPOINTER_REG_22_ & n73320;
  assign n73344 = ~P2_P2_PHYADDRPOINTER_REG_23_ & n73343;
  assign n73345 = P2_P2_PHYADDRPOINTER_REG_23_ & ~n73343;
  assign n73346 = ~n73344 & ~n73345;
  assign n73347 = n72831 & ~n73346;
  assign n73348 = ~n72188 & n72826;
  assign n73349 = P2_P2_PHYADDRPOINTER_REG_22_ & n73326;
  assign n73350 = ~P2_P2_PHYADDRPOINTER_REG_23_ & n73349;
  assign n73351 = P2_P2_PHYADDRPOINTER_REG_23_ & ~n73349;
  assign n73352 = ~n73350 & ~n73351;
  assign n73353 = n72833 & ~n73352;
  assign n73354 = n72206 & n72828;
  assign n73355 = P2_P2_PHYADDRPOINTER_REG_23_ & n72824;
  assign n73356 = P2_P2_REIP_REG_23_ & n72842;
  assign n73357 = n72840 & ~n73352;
  assign n73358 = n72170 & n72837;
  assign n73359 = ~n73355 & ~n73356;
  assign n73360 = ~n73357 & n73359;
  assign n73361 = ~n73358 & n73360;
  assign n73362 = ~n73347 & ~n73348;
  assign n73363 = ~n73353 & n73362;
  assign n73364 = ~n73354 & n73363;
  assign n13561 = ~n73361 | ~n73364;
  assign n73366 = P2_P2_PHYADDRPOINTER_REG_23_ & n73343;
  assign n73367 = ~P2_P2_PHYADDRPOINTER_REG_24_ & n73366;
  assign n73368 = P2_P2_PHYADDRPOINTER_REG_24_ & ~n73366;
  assign n73369 = ~n73367 & ~n73368;
  assign n73370 = n72831 & ~n73369;
  assign n73371 = ~n72263 & n72826;
  assign n73372 = P2_P2_PHYADDRPOINTER_REG_23_ & n73349;
  assign n73373 = ~P2_P2_PHYADDRPOINTER_REG_24_ & n73372;
  assign n73374 = P2_P2_PHYADDRPOINTER_REG_24_ & ~n73372;
  assign n73375 = ~n73373 & ~n73374;
  assign n73376 = n72833 & ~n73375;
  assign n73377 = ~n72271 & n72828;
  assign n73378 = P2_P2_PHYADDRPOINTER_REG_24_ & n72824;
  assign n73379 = P2_P2_REIP_REG_24_ & n72842;
  assign n73380 = n72840 & ~n73375;
  assign n73381 = ~n72236 & n72837;
  assign n73382 = ~n73378 & ~n73379;
  assign n73383 = ~n73380 & n73382;
  assign n73384 = ~n73381 & n73383;
  assign n73385 = ~n73370 & ~n73371;
  assign n73386 = ~n73376 & n73385;
  assign n73387 = ~n73377 & n73386;
  assign n13566 = ~n73384 | ~n73387;
  assign n73389 = P2_P2_PHYADDRPOINTER_REG_24_ & n73366;
  assign n73390 = ~P2_P2_PHYADDRPOINTER_REG_25_ & n73389;
  assign n73391 = P2_P2_PHYADDRPOINTER_REG_25_ & ~n73389;
  assign n73392 = ~n73390 & ~n73391;
  assign n73393 = n72831 & ~n73392;
  assign n73394 = ~n72340 & n72826;
  assign n73395 = P2_P2_PHYADDRPOINTER_REG_24_ & n73372;
  assign n73396 = ~P2_P2_PHYADDRPOINTER_REG_25_ & n73395;
  assign n73397 = P2_P2_PHYADDRPOINTER_REG_25_ & ~n73395;
  assign n73398 = ~n73396 & ~n73397;
  assign n73399 = n72833 & ~n73398;
  assign n73400 = n72346 & n72828;
  assign n73401 = P2_P2_PHYADDRPOINTER_REG_25_ & n72824;
  assign n73402 = P2_P2_REIP_REG_25_ & n72842;
  assign n73403 = n72840 & ~n73398;
  assign n73404 = n72312 & n72837;
  assign n73405 = ~n73401 & ~n73402;
  assign n73406 = ~n73403 & n73405;
  assign n73407 = ~n73404 & n73406;
  assign n73408 = ~n73393 & ~n73394;
  assign n73409 = ~n73399 & n73408;
  assign n73410 = ~n73400 & n73409;
  assign n13571 = ~n73407 | ~n73410;
  assign n73412 = P2_P2_PHYADDRPOINTER_REG_25_ & n73389;
  assign n73413 = ~P2_P2_PHYADDRPOINTER_REG_26_ & n73412;
  assign n73414 = P2_P2_PHYADDRPOINTER_REG_26_ & ~n73412;
  assign n73415 = ~n73413 & ~n73414;
  assign n73416 = n72831 & ~n73415;
  assign n73417 = n72381 & n72826;
  assign n73418 = P2_P2_PHYADDRPOINTER_REG_25_ & n73395;
  assign n73419 = ~P2_P2_PHYADDRPOINTER_REG_26_ & n73418;
  assign n73420 = P2_P2_PHYADDRPOINTER_REG_26_ & ~n73418;
  assign n73421 = ~n73419 & ~n73420;
  assign n73422 = n72833 & ~n73421;
  assign n73423 = n72385 & n72828;
  assign n73424 = P2_P2_PHYADDRPOINTER_REG_26_ & n72824;
  assign n73425 = n72423 & n72837;
  assign n73426 = n72840 & ~n73421;
  assign n73427 = P2_P2_REIP_REG_26_ & n72842;
  assign n73428 = ~n73424 & ~n73425;
  assign n73429 = ~n73426 & n73428;
  assign n73430 = ~n73427 & n73429;
  assign n73431 = ~n73416 & ~n73417;
  assign n73432 = ~n73422 & n73431;
  assign n73433 = ~n73423 & n73432;
  assign n13576 = ~n73430 | ~n73433;
  assign n73435 = P2_P2_PHYADDRPOINTER_REG_26_ & n73412;
  assign n73436 = ~P2_P2_PHYADDRPOINTER_REG_27_ & n73435;
  assign n73437 = P2_P2_PHYADDRPOINTER_REG_27_ & ~n73435;
  assign n73438 = ~n73436 & ~n73437;
  assign n73439 = n72831 & ~n73438;
  assign n73440 = ~n72452 & n72826;
  assign n73441 = P2_P2_PHYADDRPOINTER_REG_26_ & n73418;
  assign n73442 = ~P2_P2_PHYADDRPOINTER_REG_27_ & n73441;
  assign n73443 = P2_P2_PHYADDRPOINTER_REG_27_ & ~n73441;
  assign n73444 = ~n73442 & ~n73443;
  assign n73445 = n72833 & ~n73444;
  assign n73446 = ~n72456 & n72828;
  assign n73447 = P2_P2_PHYADDRPOINTER_REG_27_ & n72824;
  assign n73448 = ~n72494 & n72837;
  assign n73449 = n72840 & ~n73444;
  assign n73450 = P2_P2_REIP_REG_27_ & n72842;
  assign n73451 = ~n73447 & ~n73448;
  assign n73452 = ~n73449 & n73451;
  assign n73453 = ~n73450 & n73452;
  assign n73454 = ~n73439 & ~n73440;
  assign n73455 = ~n73445 & n73454;
  assign n73456 = ~n73446 & n73455;
  assign n13581 = ~n73453 | ~n73456;
  assign n73458 = n72530 & n72826;
  assign n73459 = n72535 & n72828;
  assign n73460 = P2_P2_PHYADDRPOINTER_REG_27_ & n73435;
  assign n73461 = ~P2_P2_PHYADDRPOINTER_REG_28_ & n73460;
  assign n73462 = P2_P2_PHYADDRPOINTER_REG_28_ & ~n73460;
  assign n73463 = ~n73461 & ~n73462;
  assign n73464 = n72831 & ~n73463;
  assign n73465 = P2_P2_PHYADDRPOINTER_REG_27_ & n73441;
  assign n73466 = ~P2_P2_PHYADDRPOINTER_REG_28_ & n73465;
  assign n73467 = P2_P2_PHYADDRPOINTER_REG_28_ & ~n73465;
  assign n73468 = ~n73466 & ~n73467;
  assign n73469 = n72833 & ~n73468;
  assign n73470 = P2_P2_PHYADDRPOINTER_REG_28_ & n72824;
  assign n73471 = n72574 & n72837;
  assign n73472 = n72840 & ~n73468;
  assign n73473 = P2_P2_REIP_REG_28_ & n72842;
  assign n73474 = ~n73470 & ~n73471;
  assign n73475 = ~n73472 & n73474;
  assign n73476 = ~n73473 & n73475;
  assign n73477 = ~n73458 & ~n73459;
  assign n73478 = ~n73464 & n73477;
  assign n73479 = ~n73469 & n73478;
  assign n13586 = ~n73476 | ~n73479;
  assign n73481 = ~n72603 & n72826;
  assign n73482 = n72607 & n72828;
  assign n73483 = P2_P2_PHYADDRPOINTER_REG_28_ & n73460;
  assign n73484 = ~P2_P2_PHYADDRPOINTER_REG_29_ & n73483;
  assign n73485 = P2_P2_PHYADDRPOINTER_REG_29_ & ~n73483;
  assign n73486 = ~n73484 & ~n73485;
  assign n73487 = n72831 & ~n73486;
  assign n73488 = P2_P2_PHYADDRPOINTER_REG_28_ & n73465;
  assign n73489 = ~P2_P2_PHYADDRPOINTER_REG_29_ & n73488;
  assign n73490 = P2_P2_PHYADDRPOINTER_REG_29_ & ~n73488;
  assign n73491 = ~n73489 & ~n73490;
  assign n73492 = n72833 & ~n73491;
  assign n73493 = P2_P2_PHYADDRPOINTER_REG_29_ & n72824;
  assign n73494 = P2_P2_REIP_REG_29_ & n72842;
  assign n73495 = n72645 & n72837;
  assign n73496 = n72840 & ~n73491;
  assign n73497 = ~n73493 & ~n73494;
  assign n73498 = ~n73495 & n73497;
  assign n73499 = ~n73496 & n73498;
  assign n73500 = ~n73481 & ~n73482;
  assign n73501 = ~n73487 & n73500;
  assign n73502 = ~n73492 & n73501;
  assign n13591 = ~n73499 | ~n73502;
  assign n73504 = ~n72675 & n72826;
  assign n73505 = ~n72679 & n72828;
  assign n73506 = P2_P2_PHYADDRPOINTER_REG_29_ & n73483;
  assign n73507 = ~P2_P2_PHYADDRPOINTER_REG_30_ & n73506;
  assign n73508 = P2_P2_PHYADDRPOINTER_REG_30_ & ~n73506;
  assign n73509 = ~n73507 & ~n73508;
  assign n73510 = n72831 & ~n73509;
  assign n73511 = P2_P2_PHYADDRPOINTER_REG_29_ & n73488;
  assign n73512 = ~P2_P2_PHYADDRPOINTER_REG_30_ & n73511;
  assign n73513 = P2_P2_PHYADDRPOINTER_REG_30_ & ~n73511;
  assign n73514 = ~n73512 & ~n73513;
  assign n73515 = n72833 & ~n73514;
  assign n73516 = P2_P2_PHYADDRPOINTER_REG_30_ & n72824;
  assign n73517 = P2_P2_REIP_REG_30_ & n72842;
  assign n73518 = ~n72717 & n72837;
  assign n73519 = n72840 & ~n73514;
  assign n73520 = ~n73516 & ~n73517;
  assign n73521 = ~n73518 & n73520;
  assign n73522 = ~n73519 & n73521;
  assign n73523 = ~n73504 & ~n73505;
  assign n73524 = ~n73510 & n73523;
  assign n73525 = ~n73515 & n73524;
  assign n13596 = ~n73522 | ~n73525;
  assign n73527 = n72788 & n72826;
  assign n73528 = P2_P2_PHYADDRPOINTER_REG_30_ & n73506;
  assign n73529 = ~P2_P2_PHYADDRPOINTER_REG_31_ & n73528;
  assign n73530 = P2_P2_PHYADDRPOINTER_REG_31_ & ~n73528;
  assign n73531 = ~n73529 & ~n73530;
  assign n73532 = n72831 & ~n73531;
  assign n73533 = ~n72793 & n72828;
  assign n73534 = P2_P2_PHYADDRPOINTER_REG_30_ & n73511;
  assign n73535 = ~P2_P2_PHYADDRPOINTER_REG_31_ & n73534;
  assign n73536 = P2_P2_PHYADDRPOINTER_REG_31_ & ~n73534;
  assign n73537 = ~n73535 & ~n73536;
  assign n73538 = n72833 & ~n73537;
  assign n73539 = P2_P2_PHYADDRPOINTER_REG_31_ & n72824;
  assign n73540 = P2_P2_REIP_REG_31_ & n72842;
  assign n73541 = ~n72741 & n72837;
  assign n73542 = n72840 & ~n73537;
  assign n73543 = ~n73539 & ~n73540;
  assign n73544 = ~n73541 & n73543;
  assign n73545 = ~n73542 & n73544;
  assign n73546 = ~n73527 & ~n73532;
  assign n73547 = ~n73533 & n73546;
  assign n73548 = ~n73538 & n73547;
  assign n13601 = ~n73545 | ~n73548;
  assign n73550 = P2_BUF1_REG_15_ & n12836_1;
  assign n73551 = P2_BUF2_REG_15_ & ~n12836_1;
  assign n73552 = ~n73550 & ~n73551;
  assign n73553 = ~n67541 & n67997;
  assign n73554 = n67966 & n73553;
  assign n73555 = ~n68153 & ~n73554;
  assign n73556 = n68268 & ~n73555;
  assign n73557 = ~n67882 & n73556;
  assign n73558 = ~n73552 & n73557;
  assign n73559 = n67882 & n73556;
  assign n73560 = P2_P2_EAX_REG_15_ & n73559;
  assign n73561 = P2_P2_LWORD_REG_15_ & ~n73556;
  assign n73562 = ~n73558 & ~n73560;
  assign n13606 = n73561 | ~n73562;
  assign n73564 = P2_BUF1_REG_14_ & n12836_1;
  assign n73565 = P2_BUF2_REG_14_ & ~n12836_1;
  assign n73566 = ~n73564 & ~n73565;
  assign n73567 = n73557 & ~n73566;
  assign n73568 = P2_P2_EAX_REG_14_ & n73559;
  assign n73569 = P2_P2_LWORD_REG_14_ & ~n73556;
  assign n73570 = ~n73567 & ~n73568;
  assign n13611 = n73569 | ~n73570;
  assign n73572 = P2_BUF1_REG_13_ & n12836_1;
  assign n73573 = P2_BUF2_REG_13_ & ~n12836_1;
  assign n73574 = ~n73572 & ~n73573;
  assign n73575 = n73557 & ~n73574;
  assign n73576 = P2_P2_EAX_REG_13_ & n73559;
  assign n73577 = P2_P2_LWORD_REG_13_ & ~n73556;
  assign n73578 = ~n73575 & ~n73576;
  assign n13616 = n73577 | ~n73578;
  assign n73580 = P2_BUF1_REG_12_ & n12836_1;
  assign n73581 = P2_BUF2_REG_12_ & ~n12836_1;
  assign n73582 = ~n73580 & ~n73581;
  assign n73583 = n73557 & ~n73582;
  assign n73584 = P2_P2_EAX_REG_12_ & n73559;
  assign n73585 = P2_P2_LWORD_REG_12_ & ~n73556;
  assign n73586 = ~n73583 & ~n73584;
  assign n13621 = n73585 | ~n73586;
  assign n73588 = P2_BUF1_REG_11_ & n12836_1;
  assign n73589 = P2_BUF2_REG_11_ & ~n12836_1;
  assign n73590 = ~n73588 & ~n73589;
  assign n73591 = n73557 & ~n73590;
  assign n73592 = P2_P2_EAX_REG_11_ & n73559;
  assign n73593 = P2_P2_LWORD_REG_11_ & ~n73556;
  assign n73594 = ~n73591 & ~n73592;
  assign n13626 = n73593 | ~n73594;
  assign n73596 = P2_BUF1_REG_10_ & n12836_1;
  assign n73597 = P2_BUF2_REG_10_ & ~n12836_1;
  assign n73598 = ~n73596 & ~n73597;
  assign n73599 = n73557 & ~n73598;
  assign n73600 = P2_P2_EAX_REG_10_ & n73559;
  assign n73601 = P2_P2_LWORD_REG_10_ & ~n73556;
  assign n73602 = ~n73599 & ~n73600;
  assign n13631 = n73601 | ~n73602;
  assign n73604 = P2_BUF1_REG_9_ & n12836_1;
  assign n73605 = P2_BUF2_REG_9_ & ~n12836_1;
  assign n73606 = ~n73604 & ~n73605;
  assign n73607 = n73557 & ~n73606;
  assign n73608 = P2_P2_EAX_REG_9_ & n73559;
  assign n73609 = P2_P2_LWORD_REG_9_ & ~n73556;
  assign n73610 = ~n73607 & ~n73608;
  assign n13636 = n73609 | ~n73610;
  assign n73612 = P2_BUF1_REG_8_ & n12836_1;
  assign n73613 = P2_BUF2_REG_8_ & ~n12836_1;
  assign n73614 = ~n73612 & ~n73613;
  assign n73615 = n73557 & ~n73614;
  assign n73616 = P2_P2_EAX_REG_8_ & n73559;
  assign n73617 = P2_P2_LWORD_REG_8_ & ~n73556;
  assign n73618 = ~n73615 & ~n73616;
  assign n13641 = n73617 | ~n73618;
  assign n73620 = ~n68405 & n73557;
  assign n73621 = P2_P2_EAX_REG_7_ & n73559;
  assign n73622 = P2_P2_LWORD_REG_7_ & ~n73556;
  assign n73623 = ~n73620 & ~n73621;
  assign n13646 = n73622 | ~n73623;
  assign n73625 = ~n68427 & n73557;
  assign n73626 = P2_P2_EAX_REG_6_ & n73559;
  assign n73627 = P2_P2_LWORD_REG_6_ & ~n73556;
  assign n73628 = ~n73625 & ~n73626;
  assign n13651 = n73627 | ~n73628;
  assign n73630 = ~n68449 & n73557;
  assign n73631 = P2_P2_EAX_REG_5_ & n73559;
  assign n73632 = P2_P2_LWORD_REG_5_ & ~n73556;
  assign n73633 = ~n73630 & ~n73631;
  assign n13656 = n73632 | ~n73633;
  assign n73635 = ~n68471 & n73557;
  assign n73636 = P2_P2_EAX_REG_4_ & n73559;
  assign n73637 = P2_P2_LWORD_REG_4_ & ~n73556;
  assign n73638 = ~n73635 & ~n73636;
  assign n13661 = n73637 | ~n73638;
  assign n73640 = ~n68493 & n73557;
  assign n73641 = P2_P2_EAX_REG_3_ & n73559;
  assign n73642 = P2_P2_LWORD_REG_3_ & ~n73556;
  assign n73643 = ~n73640 & ~n73641;
  assign n13666 = n73642 | ~n73643;
  assign n73645 = ~n68515 & n73557;
  assign n73646 = P2_P2_EAX_REG_2_ & n73559;
  assign n73647 = P2_P2_LWORD_REG_2_ & ~n73556;
  assign n73648 = ~n73645 & ~n73646;
  assign n13671 = n73647 | ~n73648;
  assign n73650 = ~n68537 & n73557;
  assign n73651 = P2_P2_EAX_REG_1_ & n73559;
  assign n73652 = P2_P2_LWORD_REG_1_ & ~n73556;
  assign n73653 = ~n73650 & ~n73651;
  assign n13676 = n73652 | ~n73653;
  assign n73655 = ~n68559 & n73557;
  assign n73656 = P2_P2_EAX_REG_0_ & n73559;
  assign n73657 = P2_P2_LWORD_REG_0_ & ~n73556;
  assign n73658 = ~n73655 & ~n73656;
  assign n13681 = n73657 | ~n73658;
  assign n73660 = P2_P2_EAX_REG_30_ & n73559;
  assign n73661 = P2_P2_UWORD_REG_14_ & ~n73556;
  assign n73662 = ~n73567 & ~n73660;
  assign n13686 = n73661 | ~n73662;
  assign n73664 = P2_P2_EAX_REG_29_ & n73559;
  assign n73665 = P2_P2_UWORD_REG_13_ & ~n73556;
  assign n73666 = ~n73575 & ~n73664;
  assign n13691 = n73665 | ~n73666;
  assign n73668 = P2_P2_EAX_REG_28_ & n73559;
  assign n73669 = P2_P2_UWORD_REG_12_ & ~n73556;
  assign n73670 = ~n73583 & ~n73668;
  assign n13696 = n73669 | ~n73670;
  assign n73672 = P2_P2_EAX_REG_27_ & n73559;
  assign n73673 = P2_P2_UWORD_REG_11_ & ~n73556;
  assign n73674 = ~n73591 & ~n73672;
  assign n13701 = n73673 | ~n73674;
  assign n73676 = P2_P2_EAX_REG_26_ & n73559;
  assign n73677 = P2_P2_UWORD_REG_10_ & ~n73556;
  assign n73678 = ~n73599 & ~n73676;
  assign n13706 = n73677 | ~n73678;
  assign n73680 = P2_P2_EAX_REG_25_ & n73559;
  assign n73681 = P2_P2_UWORD_REG_9_ & ~n73556;
  assign n73682 = ~n73607 & ~n73680;
  assign n13711 = n73681 | ~n73682;
  assign n73684 = P2_P2_EAX_REG_24_ & n73559;
  assign n73685 = P2_P2_UWORD_REG_8_ & ~n73556;
  assign n73686 = ~n73615 & ~n73684;
  assign n13716 = n73685 | ~n73686;
  assign n73688 = P2_P2_EAX_REG_23_ & n73559;
  assign n73689 = P2_P2_UWORD_REG_7_ & ~n73556;
  assign n73690 = ~n73620 & ~n73688;
  assign n13721 = n73689 | ~n73690;
  assign n73692 = P2_P2_EAX_REG_22_ & n73559;
  assign n73693 = P2_P2_UWORD_REG_6_ & ~n73556;
  assign n73694 = ~n73625 & ~n73692;
  assign n13726 = n73693 | ~n73694;
  assign n73696 = P2_P2_EAX_REG_21_ & n73559;
  assign n73697 = P2_P2_UWORD_REG_5_ & ~n73556;
  assign n73698 = ~n73630 & ~n73696;
  assign n13731 = n73697 | ~n73698;
  assign n73700 = P2_P2_EAX_REG_20_ & n73559;
  assign n73701 = P2_P2_UWORD_REG_4_ & ~n73556;
  assign n73702 = ~n73635 & ~n73700;
  assign n13736 = n73701 | ~n73702;
  assign n73704 = P2_P2_EAX_REG_19_ & n73559;
  assign n73705 = P2_P2_UWORD_REG_3_ & ~n73556;
  assign n73706 = ~n73640 & ~n73704;
  assign n13741 = n73705 | ~n73706;
  assign n73708 = P2_P2_EAX_REG_18_ & n73559;
  assign n73709 = P2_P2_UWORD_REG_2_ & ~n73556;
  assign n73710 = ~n73645 & ~n73708;
  assign n13746 = n73709 | ~n73710;
  assign n73712 = P2_P2_EAX_REG_17_ & n73559;
  assign n73713 = P2_P2_UWORD_REG_1_ & ~n73556;
  assign n73714 = ~n73650 & ~n73712;
  assign n13751 = n73713 | ~n73714;
  assign n73716 = P2_P2_EAX_REG_16_ & n73559;
  assign n73717 = P2_P2_UWORD_REG_0_ & ~n73556;
  assign n73718 = ~n73655 & ~n73716;
  assign n13756 = n73717 | ~n73718;
  assign n73720 = ~P2_P2_STATE2_REG_0_ & n67626;
  assign n73721 = n67632 & n68268;
  assign n73722 = ~n68154 & n73721;
  assign n73723 = ~n73720 & ~n73722;
  assign n73724 = P2_P2_STATE2_REG_0_ & ~n73723;
  assign n73725 = P2_P2_EAX_REG_0_ & n73724;
  assign n73726 = ~P2_P2_STATE2_REG_0_ & ~n73723;
  assign n73727 = P2_P2_LWORD_REG_0_ & n73726;
  assign n73728 = P2_P2_DATAO_REG_0_ & n73723;
  assign n73729 = ~n73725 & ~n73727;
  assign n13761 = n73728 | ~n73729;
  assign n73731 = P2_P2_EAX_REG_1_ & n73724;
  assign n73732 = P2_P2_LWORD_REG_1_ & n73726;
  assign n73733 = P2_P2_DATAO_REG_1_ & n73723;
  assign n73734 = ~n73731 & ~n73732;
  assign n13766 = n73733 | ~n73734;
  assign n73736 = P2_P2_EAX_REG_2_ & n73724;
  assign n73737 = P2_P2_LWORD_REG_2_ & n73726;
  assign n73738 = P2_P2_DATAO_REG_2_ & n73723;
  assign n73739 = ~n73736 & ~n73737;
  assign n13771 = n73738 | ~n73739;
  assign n73741 = P2_P2_EAX_REG_3_ & n73724;
  assign n73742 = P2_P2_LWORD_REG_3_ & n73726;
  assign n73743 = P2_P2_DATAO_REG_3_ & n73723;
  assign n73744 = ~n73741 & ~n73742;
  assign n13776 = n73743 | ~n73744;
  assign n73746 = P2_P2_EAX_REG_4_ & n73724;
  assign n73747 = P2_P2_LWORD_REG_4_ & n73726;
  assign n73748 = P2_P2_DATAO_REG_4_ & n73723;
  assign n73749 = ~n73746 & ~n73747;
  assign n13781 = n73748 | ~n73749;
  assign n73751 = P2_P2_EAX_REG_5_ & n73724;
  assign n73752 = P2_P2_LWORD_REG_5_ & n73726;
  assign n73753 = P2_P2_DATAO_REG_5_ & n73723;
  assign n73754 = ~n73751 & ~n73752;
  assign n13786 = n73753 | ~n73754;
  assign n73756 = P2_P2_EAX_REG_6_ & n73724;
  assign n73757 = P2_P2_LWORD_REG_6_ & n73726;
  assign n73758 = P2_P2_DATAO_REG_6_ & n73723;
  assign n73759 = ~n73756 & ~n73757;
  assign n13791 = n73758 | ~n73759;
  assign n73761 = P2_P2_EAX_REG_7_ & n73724;
  assign n73762 = P2_P2_LWORD_REG_7_ & n73726;
  assign n73763 = P2_P2_DATAO_REG_7_ & n73723;
  assign n73764 = ~n73761 & ~n73762;
  assign n13796 = n73763 | ~n73764;
  assign n73766 = P2_P2_EAX_REG_8_ & n73724;
  assign n73767 = P2_P2_LWORD_REG_8_ & n73726;
  assign n73768 = P2_P2_DATAO_REG_8_ & n73723;
  assign n73769 = ~n73766 & ~n73767;
  assign n13801 = n73768 | ~n73769;
  assign n73771 = P2_P2_EAX_REG_9_ & n73724;
  assign n73772 = P2_P2_LWORD_REG_9_ & n73726;
  assign n73773 = P2_P2_DATAO_REG_9_ & n73723;
  assign n73774 = ~n73771 & ~n73772;
  assign n13806 = n73773 | ~n73774;
  assign n73776 = P2_P2_EAX_REG_10_ & n73724;
  assign n73777 = P2_P2_LWORD_REG_10_ & n73726;
  assign n73778 = P2_P2_DATAO_REG_10_ & n73723;
  assign n73779 = ~n73776 & ~n73777;
  assign n13811 = n73778 | ~n73779;
  assign n73781 = P2_P2_EAX_REG_11_ & n73724;
  assign n73782 = P2_P2_LWORD_REG_11_ & n73726;
  assign n73783 = P2_P2_DATAO_REG_11_ & n73723;
  assign n73784 = ~n73781 & ~n73782;
  assign n13816 = n73783 | ~n73784;
  assign n73786 = P2_P2_EAX_REG_12_ & n73724;
  assign n73787 = P2_P2_LWORD_REG_12_ & n73726;
  assign n73788 = P2_P2_DATAO_REG_12_ & n73723;
  assign n73789 = ~n73786 & ~n73787;
  assign n13821 = n73788 | ~n73789;
  assign n73791 = P2_P2_EAX_REG_13_ & n73724;
  assign n73792 = P2_P2_LWORD_REG_13_ & n73726;
  assign n73793 = P2_P2_DATAO_REG_13_ & n73723;
  assign n73794 = ~n73791 & ~n73792;
  assign n13826 = n73793 | ~n73794;
  assign n73796 = P2_P2_EAX_REG_14_ & n73724;
  assign n73797 = P2_P2_LWORD_REG_14_ & n73726;
  assign n73798 = P2_P2_DATAO_REG_14_ & n73723;
  assign n73799 = ~n73796 & ~n73797;
  assign n13831 = n73798 | ~n73799;
  assign n73801 = P2_P2_EAX_REG_15_ & n73724;
  assign n73802 = P2_P2_LWORD_REG_15_ & n73726;
  assign n73803 = P2_P2_DATAO_REG_15_ & n73723;
  assign n73804 = ~n73801 & ~n73802;
  assign n13836 = n73803 | ~n73804;
  assign n73806 = P2_P2_UWORD_REG_0_ & n73726;
  assign n73807 = P2_P2_DATAO_REG_16_ & n73723;
  assign n73808 = ~n73806 & ~n73807;
  assign n73809 = ~n67913 & n73724;
  assign n73810 = P2_P2_EAX_REG_16_ & n73809;
  assign n13841 = ~n73808 | n73810;
  assign n73812 = P2_P2_UWORD_REG_1_ & n73726;
  assign n73813 = P2_P2_DATAO_REG_17_ & n73723;
  assign n73814 = ~n73812 & ~n73813;
  assign n73815 = P2_P2_EAX_REG_17_ & n73809;
  assign n13846 = ~n73814 | n73815;
  assign n73817 = P2_P2_UWORD_REG_2_ & n73726;
  assign n73818 = P2_P2_DATAO_REG_18_ & n73723;
  assign n73819 = ~n73817 & ~n73818;
  assign n73820 = P2_P2_EAX_REG_18_ & n73809;
  assign n13851 = ~n73819 | n73820;
  assign n73822 = P2_P2_UWORD_REG_3_ & n73726;
  assign n73823 = P2_P2_DATAO_REG_19_ & n73723;
  assign n73824 = ~n73822 & ~n73823;
  assign n73825 = P2_P2_EAX_REG_19_ & n73809;
  assign n13856 = ~n73824 | n73825;
  assign n73827 = P2_P2_UWORD_REG_4_ & n73726;
  assign n73828 = P2_P2_DATAO_REG_20_ & n73723;
  assign n73829 = ~n73827 & ~n73828;
  assign n73830 = P2_P2_EAX_REG_20_ & n73809;
  assign n13861 = ~n73829 | n73830;
  assign n73832 = P2_P2_UWORD_REG_5_ & n73726;
  assign n73833 = P2_P2_DATAO_REG_21_ & n73723;
  assign n73834 = ~n73832 & ~n73833;
  assign n73835 = P2_P2_EAX_REG_21_ & n73809;
  assign n13866 = ~n73834 | n73835;
  assign n73837 = P2_P2_UWORD_REG_6_ & n73726;
  assign n73838 = P2_P2_DATAO_REG_22_ & n73723;
  assign n73839 = ~n73837 & ~n73838;
  assign n73840 = P2_P2_EAX_REG_22_ & n73809;
  assign n13871 = ~n73839 | n73840;
  assign n73842 = P2_P2_UWORD_REG_7_ & n73726;
  assign n73843 = P2_P2_DATAO_REG_23_ & n73723;
  assign n73844 = ~n73842 & ~n73843;
  assign n73845 = P2_P2_EAX_REG_23_ & n73809;
  assign n13876 = ~n73844 | n73845;
  assign n73847 = P2_P2_UWORD_REG_8_ & n73726;
  assign n73848 = P2_P2_DATAO_REG_24_ & n73723;
  assign n73849 = ~n73847 & ~n73848;
  assign n73850 = P2_P2_EAX_REG_24_ & n73809;
  assign n13881 = ~n73849 | n73850;
  assign n73852 = P2_P2_UWORD_REG_9_ & n73726;
  assign n73853 = P2_P2_DATAO_REG_25_ & n73723;
  assign n73854 = ~n73852 & ~n73853;
  assign n73855 = P2_P2_EAX_REG_25_ & n73809;
  assign n13886 = ~n73854 | n73855;
  assign n73857 = P2_P2_UWORD_REG_10_ & n73726;
  assign n73858 = P2_P2_DATAO_REG_26_ & n73723;
  assign n73859 = ~n73857 & ~n73858;
  assign n73860 = P2_P2_EAX_REG_26_ & n73809;
  assign n13891 = ~n73859 | n73860;
  assign n73862 = P2_P2_UWORD_REG_11_ & n73726;
  assign n73863 = P2_P2_DATAO_REG_27_ & n73723;
  assign n73864 = ~n73862 & ~n73863;
  assign n73865 = P2_P2_EAX_REG_27_ & n73809;
  assign n13896 = ~n73864 | n73865;
  assign n73867 = P2_P2_UWORD_REG_12_ & n73726;
  assign n73868 = P2_P2_DATAO_REG_28_ & n73723;
  assign n73869 = ~n73867 & ~n73868;
  assign n73870 = P2_P2_EAX_REG_28_ & n73809;
  assign n13901 = ~n73869 | n73870;
  assign n73872 = P2_P2_UWORD_REG_13_ & n73726;
  assign n73873 = P2_P2_DATAO_REG_29_ & n73723;
  assign n73874 = ~n73872 & ~n73873;
  assign n73875 = P2_P2_EAX_REG_29_ & n73809;
  assign n13906 = ~n73874 | n73875;
  assign n73877 = P2_P2_UWORD_REG_14_ & n73726;
  assign n73878 = P2_P2_DATAO_REG_30_ & n73723;
  assign n73879 = ~n73877 & ~n73878;
  assign n73880 = P2_P2_EAX_REG_30_ & n73809;
  assign n13911 = ~n73879 | n73880;
  assign n13916 = P2_P2_DATAO_REG_31_ & n73723;
  assign n73883 = n68148 & ~n68212;
  assign n73884 = n68268 & ~n73883;
  assign n73885 = n68002 & n73884;
  assign n73886 = ~n70050 & n73885;
  assign n73887 = ~n67785 & n73884;
  assign n73888 = ~n68002 & n73887;
  assign n73889 = ~n68559 & n73888;
  assign n73890 = P2_P2_EAX_REG_0_ & ~n73884;
  assign n73891 = n67785 & n73884;
  assign n73892 = ~P2_P2_EAX_REG_0_ & n73891;
  assign n73893 = ~n73890 & ~n73892;
  assign n73894 = ~n73886 & ~n73889;
  assign n13921 = ~n73893 | ~n73894;
  assign n73896 = ~n70168 & n73885;
  assign n73897 = ~n68537 & n73888;
  assign n73898 = P2_P2_EAX_REG_1_ & ~n73884;
  assign n73899 = ~P2_P2_EAX_REG_0_ & P2_P2_EAX_REG_1_;
  assign n73900 = P2_P2_EAX_REG_0_ & ~P2_P2_EAX_REG_1_;
  assign n73901 = ~n73899 & ~n73900;
  assign n73902 = n73891 & ~n73901;
  assign n73903 = ~n73898 & ~n73902;
  assign n73904 = ~n73896 & ~n73897;
  assign n13926 = ~n73903 | ~n73904;
  assign n73906 = ~n70288 & n73885;
  assign n73907 = ~n68515 & n73888;
  assign n73908 = P2_P2_EAX_REG_2_ & ~n73884;
  assign n73909 = P2_P2_EAX_REG_0_ & P2_P2_EAX_REG_1_;
  assign n73910 = ~P2_P2_EAX_REG_2_ & n73909;
  assign n73911 = P2_P2_EAX_REG_2_ & ~n73909;
  assign n73912 = ~n73910 & ~n73911;
  assign n73913 = n73891 & ~n73912;
  assign n73914 = ~n73908 & ~n73913;
  assign n73915 = ~n73906 & ~n73907;
  assign n13931 = ~n73914 | ~n73915;
  assign n73917 = ~n70412 & n73885;
  assign n73918 = ~n68493 & n73888;
  assign n73919 = P2_P2_EAX_REG_3_ & ~n73884;
  assign n73920 = P2_P2_EAX_REG_0_ & P2_P2_EAX_REG_2_;
  assign n73921 = P2_P2_EAX_REG_1_ & n73920;
  assign n73922 = P2_P2_EAX_REG_3_ & ~n73921;
  assign n73923 = ~P2_P2_EAX_REG_3_ & n73921;
  assign n73924 = ~n73922 & ~n73923;
  assign n73925 = n73891 & ~n73924;
  assign n73926 = ~n73919 & ~n73925;
  assign n73927 = ~n73917 & ~n73918;
  assign n13936 = ~n73926 | ~n73927;
  assign n73929 = ~n70539 & n73885;
  assign n73930 = ~n68471 & n73888;
  assign n73931 = P2_P2_EAX_REG_4_ & ~n73884;
  assign n73932 = P2_P2_EAX_REG_3_ & n73921;
  assign n73933 = ~P2_P2_EAX_REG_4_ & n73932;
  assign n73934 = P2_P2_EAX_REG_4_ & ~n73932;
  assign n73935 = ~n73933 & ~n73934;
  assign n73936 = n73891 & ~n73935;
  assign n73937 = ~n73931 & ~n73936;
  assign n73938 = ~n73929 & ~n73930;
  assign n13941 = ~n73937 | ~n73938;
  assign n73940 = ~n70680 & n73885;
  assign n73941 = ~n68449 & n73888;
  assign n73942 = P2_P2_EAX_REG_5_ & ~n73884;
  assign n73943 = P2_P2_EAX_REG_3_ & P2_P2_EAX_REG_4_;
  assign n73944 = n73921 & n73943;
  assign n73945 = P2_P2_EAX_REG_5_ & ~n73944;
  assign n73946 = ~P2_P2_EAX_REG_5_ & n73944;
  assign n73947 = ~n73945 & ~n73946;
  assign n73948 = n73891 & ~n73947;
  assign n73949 = ~n73942 & ~n73948;
  assign n73950 = ~n73940 & ~n73941;
  assign n13946 = ~n73949 | ~n73950;
  assign n73952 = ~n70812 & n73885;
  assign n73953 = ~n68427 & n73888;
  assign n73954 = P2_P2_EAX_REG_6_ & ~n73884;
  assign n73955 = P2_P2_EAX_REG_5_ & n73944;
  assign n73956 = ~P2_P2_EAX_REG_6_ & n73955;
  assign n73957 = P2_P2_EAX_REG_6_ & ~n73955;
  assign n73958 = ~n73956 & ~n73957;
  assign n73959 = n73891 & ~n73958;
  assign n73960 = ~n73954 & ~n73959;
  assign n73961 = ~n73952 & ~n73953;
  assign n13951 = ~n73960 | ~n73961;
  assign n73963 = ~n70084 & n73885;
  assign n73964 = ~n68405 & n73888;
  assign n73965 = P2_P2_EAX_REG_7_ & ~n73884;
  assign n73966 = P2_P2_EAX_REG_5_ & P2_P2_EAX_REG_6_;
  assign n73967 = n73944 & n73966;
  assign n73968 = P2_P2_EAX_REG_7_ & ~n73967;
  assign n73969 = ~P2_P2_EAX_REG_7_ & n73967;
  assign n73970 = ~n73968 & ~n73969;
  assign n73971 = n73891 & ~n73970;
  assign n73972 = ~n73965 & ~n73971;
  assign n73973 = ~n73963 & ~n73964;
  assign n13956 = ~n73972 | ~n73973;
  assign n73975 = ~n68162 & ~n68169;
  assign n73976 = ~n68113 & ~n73975;
  assign n73977 = n67643 & n73976;
  assign n73978 = P2_P2_INSTQUEUE_REG_15__0_ & n73977;
  assign n73979 = n67647 & n73976;
  assign n73980 = P2_P2_INSTQUEUE_REG_14__0_ & n73979;
  assign n73981 = n67634 & n73976;
  assign n73982 = P2_P2_INSTQUEUE_REG_13__0_ & n73981;
  assign n73983 = n67638 & n73976;
  assign n73984 = P2_P2_INSTQUEUE_REG_12__0_ & n73983;
  assign n73985 = ~n73978 & ~n73980;
  assign n73986 = ~n73982 & n73985;
  assign n73987 = ~n73984 & n73986;
  assign n73988 = n68113 & ~n73975;
  assign n73989 = n67643 & n73988;
  assign n73990 = P2_P2_INSTQUEUE_REG_11__0_ & n73989;
  assign n73991 = n67647 & n73988;
  assign n73992 = P2_P2_INSTQUEUE_REG_10__0_ & n73991;
  assign n73993 = n67634 & n73988;
  assign n73994 = P2_P2_INSTQUEUE_REG_9__0_ & n73993;
  assign n73995 = n67638 & n73988;
  assign n73996 = P2_P2_INSTQUEUE_REG_8__0_ & n73995;
  assign n73997 = ~n73990 & ~n73992;
  assign n73998 = ~n73994 & n73997;
  assign n73999 = ~n73996 & n73998;
  assign n74000 = ~n68113 & n73975;
  assign n74001 = n67643 & n74000;
  assign n74002 = P2_P2_INSTQUEUE_REG_7__0_ & n74001;
  assign n74003 = n67647 & n74000;
  assign n74004 = P2_P2_INSTQUEUE_REG_6__0_ & n74003;
  assign n74005 = n67634 & n74000;
  assign n74006 = P2_P2_INSTQUEUE_REG_5__0_ & n74005;
  assign n74007 = n67638 & n74000;
  assign n74008 = P2_P2_INSTQUEUE_REG_4__0_ & n74007;
  assign n74009 = ~n74002 & ~n74004;
  assign n74010 = ~n74006 & n74009;
  assign n74011 = ~n74008 & n74010;
  assign n74012 = n68113 & n73975;
  assign n74013 = n67643 & n74012;
  assign n74014 = P2_P2_INSTQUEUE_REG_3__0_ & n74013;
  assign n74015 = n67647 & n74012;
  assign n74016 = P2_P2_INSTQUEUE_REG_2__0_ & n74015;
  assign n74017 = n67634 & n74012;
  assign n74018 = P2_P2_INSTQUEUE_REG_1__0_ & n74017;
  assign n74019 = n67638 & n74012;
  assign n74020 = P2_P2_INSTQUEUE_REG_0__0_ & n74019;
  assign n74021 = ~n74014 & ~n74016;
  assign n74022 = ~n74018 & n74021;
  assign n74023 = ~n74020 & n74022;
  assign n74024 = n73987 & n73999;
  assign n74025 = n74011 & n74024;
  assign n74026 = n74023 & n74025;
  assign n74027 = n73885 & ~n74026;
  assign n74028 = ~n73614 & n73888;
  assign n74029 = P2_P2_EAX_REG_8_ & ~n73884;
  assign n74030 = P2_P2_EAX_REG_7_ & n73967;
  assign n74031 = ~P2_P2_EAX_REG_8_ & n74030;
  assign n74032 = P2_P2_EAX_REG_8_ & ~n74030;
  assign n74033 = ~n74031 & ~n74032;
  assign n74034 = n73891 & ~n74033;
  assign n74035 = ~n74029 & ~n74034;
  assign n74036 = ~n74027 & ~n74028;
  assign n13961 = ~n74035 | ~n74036;
  assign n74038 = P2_P2_INSTQUEUE_REG_15__1_ & n73977;
  assign n74039 = P2_P2_INSTQUEUE_REG_14__1_ & n73979;
  assign n74040 = P2_P2_INSTQUEUE_REG_13__1_ & n73981;
  assign n74041 = P2_P2_INSTQUEUE_REG_12__1_ & n73983;
  assign n74042 = ~n74038 & ~n74039;
  assign n74043 = ~n74040 & n74042;
  assign n74044 = ~n74041 & n74043;
  assign n74045 = P2_P2_INSTQUEUE_REG_11__1_ & n73989;
  assign n74046 = P2_P2_INSTQUEUE_REG_10__1_ & n73991;
  assign n74047 = P2_P2_INSTQUEUE_REG_9__1_ & n73993;
  assign n74048 = P2_P2_INSTQUEUE_REG_8__1_ & n73995;
  assign n74049 = ~n74045 & ~n74046;
  assign n74050 = ~n74047 & n74049;
  assign n74051 = ~n74048 & n74050;
  assign n74052 = P2_P2_INSTQUEUE_REG_7__1_ & n74001;
  assign n74053 = P2_P2_INSTQUEUE_REG_6__1_ & n74003;
  assign n74054 = P2_P2_INSTQUEUE_REG_5__1_ & n74005;
  assign n74055 = P2_P2_INSTQUEUE_REG_4__1_ & n74007;
  assign n74056 = ~n74052 & ~n74053;
  assign n74057 = ~n74054 & n74056;
  assign n74058 = ~n74055 & n74057;
  assign n74059 = P2_P2_INSTQUEUE_REG_3__1_ & n74013;
  assign n74060 = P2_P2_INSTQUEUE_REG_2__1_ & n74015;
  assign n74061 = P2_P2_INSTQUEUE_REG_1__1_ & n74017;
  assign n74062 = P2_P2_INSTQUEUE_REG_0__1_ & n74019;
  assign n74063 = ~n74059 & ~n74060;
  assign n74064 = ~n74061 & n74063;
  assign n74065 = ~n74062 & n74064;
  assign n74066 = n74044 & n74051;
  assign n74067 = n74058 & n74066;
  assign n74068 = n74065 & n74067;
  assign n74069 = n73885 & ~n74068;
  assign n74070 = ~n73606 & n73888;
  assign n74071 = P2_P2_EAX_REG_9_ & ~n73884;
  assign n74072 = P2_P2_EAX_REG_7_ & P2_P2_EAX_REG_8_;
  assign n74073 = n73967 & n74072;
  assign n74074 = P2_P2_EAX_REG_9_ & ~n74073;
  assign n74075 = ~P2_P2_EAX_REG_9_ & n74073;
  assign n74076 = ~n74074 & ~n74075;
  assign n74077 = n73891 & ~n74076;
  assign n74078 = ~n74071 & ~n74077;
  assign n74079 = ~n74069 & ~n74070;
  assign n13966 = ~n74078 | ~n74079;
  assign n74081 = P2_P2_INSTQUEUE_REG_15__2_ & n73977;
  assign n74082 = P2_P2_INSTQUEUE_REG_14__2_ & n73979;
  assign n74083 = P2_P2_INSTQUEUE_REG_13__2_ & n73981;
  assign n74084 = P2_P2_INSTQUEUE_REG_12__2_ & n73983;
  assign n74085 = ~n74081 & ~n74082;
  assign n74086 = ~n74083 & n74085;
  assign n74087 = ~n74084 & n74086;
  assign n74088 = P2_P2_INSTQUEUE_REG_11__2_ & n73989;
  assign n74089 = P2_P2_INSTQUEUE_REG_10__2_ & n73991;
  assign n74090 = P2_P2_INSTQUEUE_REG_9__2_ & n73993;
  assign n74091 = P2_P2_INSTQUEUE_REG_8__2_ & n73995;
  assign n74092 = ~n74088 & ~n74089;
  assign n74093 = ~n74090 & n74092;
  assign n74094 = ~n74091 & n74093;
  assign n74095 = P2_P2_INSTQUEUE_REG_7__2_ & n74001;
  assign n74096 = P2_P2_INSTQUEUE_REG_6__2_ & n74003;
  assign n74097 = P2_P2_INSTQUEUE_REG_5__2_ & n74005;
  assign n74098 = P2_P2_INSTQUEUE_REG_4__2_ & n74007;
  assign n74099 = ~n74095 & ~n74096;
  assign n74100 = ~n74097 & n74099;
  assign n74101 = ~n74098 & n74100;
  assign n74102 = P2_P2_INSTQUEUE_REG_3__2_ & n74013;
  assign n74103 = P2_P2_INSTQUEUE_REG_2__2_ & n74015;
  assign n74104 = P2_P2_INSTQUEUE_REG_1__2_ & n74017;
  assign n74105 = P2_P2_INSTQUEUE_REG_0__2_ & n74019;
  assign n74106 = ~n74102 & ~n74103;
  assign n74107 = ~n74104 & n74106;
  assign n74108 = ~n74105 & n74107;
  assign n74109 = n74087 & n74094;
  assign n74110 = n74101 & n74109;
  assign n74111 = n74108 & n74110;
  assign n74112 = n73885 & ~n74111;
  assign n74113 = ~n73598 & n73888;
  assign n74114 = P2_P2_EAX_REG_10_ & ~n73884;
  assign n74115 = P2_P2_EAX_REG_9_ & n74073;
  assign n74116 = ~P2_P2_EAX_REG_10_ & n74115;
  assign n74117 = P2_P2_EAX_REG_10_ & ~n74115;
  assign n74118 = ~n74116 & ~n74117;
  assign n74119 = n73891 & ~n74118;
  assign n74120 = ~n74114 & ~n74119;
  assign n74121 = ~n74112 & ~n74113;
  assign n13971 = ~n74120 | ~n74121;
  assign n74123 = P2_P2_INSTQUEUE_REG_15__3_ & n73977;
  assign n74124 = P2_P2_INSTQUEUE_REG_14__3_ & n73979;
  assign n74125 = P2_P2_INSTQUEUE_REG_13__3_ & n73981;
  assign n74126 = P2_P2_INSTQUEUE_REG_12__3_ & n73983;
  assign n74127 = ~n74123 & ~n74124;
  assign n74128 = ~n74125 & n74127;
  assign n74129 = ~n74126 & n74128;
  assign n74130 = P2_P2_INSTQUEUE_REG_11__3_ & n73989;
  assign n74131 = P2_P2_INSTQUEUE_REG_10__3_ & n73991;
  assign n74132 = P2_P2_INSTQUEUE_REG_9__3_ & n73993;
  assign n74133 = P2_P2_INSTQUEUE_REG_8__3_ & n73995;
  assign n74134 = ~n74130 & ~n74131;
  assign n74135 = ~n74132 & n74134;
  assign n74136 = ~n74133 & n74135;
  assign n74137 = P2_P2_INSTQUEUE_REG_7__3_ & n74001;
  assign n74138 = P2_P2_INSTQUEUE_REG_6__3_ & n74003;
  assign n74139 = P2_P2_INSTQUEUE_REG_5__3_ & n74005;
  assign n74140 = P2_P2_INSTQUEUE_REG_4__3_ & n74007;
  assign n74141 = ~n74137 & ~n74138;
  assign n74142 = ~n74139 & n74141;
  assign n74143 = ~n74140 & n74142;
  assign n74144 = P2_P2_INSTQUEUE_REG_3__3_ & n74013;
  assign n74145 = P2_P2_INSTQUEUE_REG_2__3_ & n74015;
  assign n74146 = P2_P2_INSTQUEUE_REG_1__3_ & n74017;
  assign n74147 = P2_P2_INSTQUEUE_REG_0__3_ & n74019;
  assign n74148 = ~n74144 & ~n74145;
  assign n74149 = ~n74146 & n74148;
  assign n74150 = ~n74147 & n74149;
  assign n74151 = n74129 & n74136;
  assign n74152 = n74143 & n74151;
  assign n74153 = n74150 & n74152;
  assign n74154 = n73885 & ~n74153;
  assign n74155 = ~n73590 & n73888;
  assign n74156 = P2_P2_EAX_REG_11_ & ~n73884;
  assign n74157 = P2_P2_EAX_REG_9_ & P2_P2_EAX_REG_10_;
  assign n74158 = n74073 & n74157;
  assign n74159 = P2_P2_EAX_REG_11_ & ~n74158;
  assign n74160 = ~P2_P2_EAX_REG_11_ & n74158;
  assign n74161 = ~n74159 & ~n74160;
  assign n74162 = n73891 & ~n74161;
  assign n74163 = ~n74156 & ~n74162;
  assign n74164 = ~n74154 & ~n74155;
  assign n13976 = ~n74163 | ~n74164;
  assign n74166 = P2_P2_INSTQUEUE_REG_15__4_ & n73977;
  assign n74167 = P2_P2_INSTQUEUE_REG_14__4_ & n73979;
  assign n74168 = P2_P2_INSTQUEUE_REG_13__4_ & n73981;
  assign n74169 = P2_P2_INSTQUEUE_REG_12__4_ & n73983;
  assign n74170 = ~n74166 & ~n74167;
  assign n74171 = ~n74168 & n74170;
  assign n74172 = ~n74169 & n74171;
  assign n74173 = P2_P2_INSTQUEUE_REG_11__4_ & n73989;
  assign n74174 = P2_P2_INSTQUEUE_REG_10__4_ & n73991;
  assign n74175 = P2_P2_INSTQUEUE_REG_9__4_ & n73993;
  assign n74176 = P2_P2_INSTQUEUE_REG_8__4_ & n73995;
  assign n74177 = ~n74173 & ~n74174;
  assign n74178 = ~n74175 & n74177;
  assign n74179 = ~n74176 & n74178;
  assign n74180 = P2_P2_INSTQUEUE_REG_7__4_ & n74001;
  assign n74181 = P2_P2_INSTQUEUE_REG_6__4_ & n74003;
  assign n74182 = P2_P2_INSTQUEUE_REG_5__4_ & n74005;
  assign n74183 = P2_P2_INSTQUEUE_REG_4__4_ & n74007;
  assign n74184 = ~n74180 & ~n74181;
  assign n74185 = ~n74182 & n74184;
  assign n74186 = ~n74183 & n74185;
  assign n74187 = P2_P2_INSTQUEUE_REG_3__4_ & n74013;
  assign n74188 = P2_P2_INSTQUEUE_REG_2__4_ & n74015;
  assign n74189 = P2_P2_INSTQUEUE_REG_1__4_ & n74017;
  assign n74190 = P2_P2_INSTQUEUE_REG_0__4_ & n74019;
  assign n74191 = ~n74187 & ~n74188;
  assign n74192 = ~n74189 & n74191;
  assign n74193 = ~n74190 & n74192;
  assign n74194 = n74172 & n74179;
  assign n74195 = n74186 & n74194;
  assign n74196 = n74193 & n74195;
  assign n74197 = n73885 & ~n74196;
  assign n74198 = ~n73582 & n73888;
  assign n74199 = P2_P2_EAX_REG_12_ & ~n73884;
  assign n74200 = P2_P2_EAX_REG_11_ & n74158;
  assign n74201 = ~P2_P2_EAX_REG_12_ & n74200;
  assign n74202 = P2_P2_EAX_REG_12_ & ~n74200;
  assign n74203 = ~n74201 & ~n74202;
  assign n74204 = n73891 & ~n74203;
  assign n74205 = ~n74199 & ~n74204;
  assign n74206 = ~n74197 & ~n74198;
  assign n13981 = ~n74205 | ~n74206;
  assign n74208 = ~n73574 & n73888;
  assign n74209 = P2_P2_INSTQUEUE_REG_15__5_ & n73977;
  assign n74210 = P2_P2_INSTQUEUE_REG_14__5_ & n73979;
  assign n74211 = P2_P2_INSTQUEUE_REG_13__5_ & n73981;
  assign n74212 = P2_P2_INSTQUEUE_REG_12__5_ & n73983;
  assign n74213 = ~n74209 & ~n74210;
  assign n74214 = ~n74211 & n74213;
  assign n74215 = ~n74212 & n74214;
  assign n74216 = P2_P2_INSTQUEUE_REG_11__5_ & n73989;
  assign n74217 = P2_P2_INSTQUEUE_REG_10__5_ & n73991;
  assign n74218 = P2_P2_INSTQUEUE_REG_9__5_ & n73993;
  assign n74219 = P2_P2_INSTQUEUE_REG_8__5_ & n73995;
  assign n74220 = ~n74216 & ~n74217;
  assign n74221 = ~n74218 & n74220;
  assign n74222 = ~n74219 & n74221;
  assign n74223 = P2_P2_INSTQUEUE_REG_7__5_ & n74001;
  assign n74224 = P2_P2_INSTQUEUE_REG_6__5_ & n74003;
  assign n74225 = P2_P2_INSTQUEUE_REG_5__5_ & n74005;
  assign n74226 = P2_P2_INSTQUEUE_REG_4__5_ & n74007;
  assign n74227 = ~n74223 & ~n74224;
  assign n74228 = ~n74225 & n74227;
  assign n74229 = ~n74226 & n74228;
  assign n74230 = P2_P2_INSTQUEUE_REG_3__5_ & n74013;
  assign n74231 = P2_P2_INSTQUEUE_REG_2__5_ & n74015;
  assign n74232 = P2_P2_INSTQUEUE_REG_1__5_ & n74017;
  assign n74233 = P2_P2_INSTQUEUE_REG_0__5_ & n74019;
  assign n74234 = ~n74230 & ~n74231;
  assign n74235 = ~n74232 & n74234;
  assign n74236 = ~n74233 & n74235;
  assign n74237 = n74215 & n74222;
  assign n74238 = n74229 & n74237;
  assign n74239 = n74236 & n74238;
  assign n74240 = n73885 & ~n74239;
  assign n74241 = P2_P2_EAX_REG_13_ & ~n73884;
  assign n74242 = ~n74240 & ~n74241;
  assign n74243 = P2_P2_EAX_REG_11_ & P2_P2_EAX_REG_12_;
  assign n74244 = n74158 & n74243;
  assign n74245 = P2_P2_EAX_REG_13_ & ~n74244;
  assign n74246 = ~P2_P2_EAX_REG_13_ & n74244;
  assign n74247 = ~n74245 & ~n74246;
  assign n74248 = n73891 & ~n74247;
  assign n74249 = ~n74208 & n74242;
  assign n13986 = n74248 | ~n74249;
  assign n74251 = ~n73566 & n73888;
  assign n74252 = P2_P2_INSTQUEUE_REG_15__6_ & n73977;
  assign n74253 = P2_P2_INSTQUEUE_REG_14__6_ & n73979;
  assign n74254 = P2_P2_INSTQUEUE_REG_13__6_ & n73981;
  assign n74255 = P2_P2_INSTQUEUE_REG_12__6_ & n73983;
  assign n74256 = ~n74252 & ~n74253;
  assign n74257 = ~n74254 & n74256;
  assign n74258 = ~n74255 & n74257;
  assign n74259 = P2_P2_INSTQUEUE_REG_11__6_ & n73989;
  assign n74260 = P2_P2_INSTQUEUE_REG_10__6_ & n73991;
  assign n74261 = P2_P2_INSTQUEUE_REG_9__6_ & n73993;
  assign n74262 = P2_P2_INSTQUEUE_REG_8__6_ & n73995;
  assign n74263 = ~n74259 & ~n74260;
  assign n74264 = ~n74261 & n74263;
  assign n74265 = ~n74262 & n74264;
  assign n74266 = P2_P2_INSTQUEUE_REG_7__6_ & n74001;
  assign n74267 = P2_P2_INSTQUEUE_REG_6__6_ & n74003;
  assign n74268 = P2_P2_INSTQUEUE_REG_5__6_ & n74005;
  assign n74269 = P2_P2_INSTQUEUE_REG_4__6_ & n74007;
  assign n74270 = ~n74266 & ~n74267;
  assign n74271 = ~n74268 & n74270;
  assign n74272 = ~n74269 & n74271;
  assign n74273 = P2_P2_INSTQUEUE_REG_3__6_ & n74013;
  assign n74274 = P2_P2_INSTQUEUE_REG_2__6_ & n74015;
  assign n74275 = P2_P2_INSTQUEUE_REG_1__6_ & n74017;
  assign n74276 = P2_P2_INSTQUEUE_REG_0__6_ & n74019;
  assign n74277 = ~n74273 & ~n74274;
  assign n74278 = ~n74275 & n74277;
  assign n74279 = ~n74276 & n74278;
  assign n74280 = n74258 & n74265;
  assign n74281 = n74272 & n74280;
  assign n74282 = n74279 & n74281;
  assign n74283 = n73885 & ~n74282;
  assign n74284 = P2_P2_EAX_REG_14_ & ~n73884;
  assign n74285 = ~n74283 & ~n74284;
  assign n74286 = P2_P2_EAX_REG_13_ & n74244;
  assign n74287 = ~P2_P2_EAX_REG_14_ & n74286;
  assign n74288 = P2_P2_EAX_REG_14_ & ~n74286;
  assign n74289 = ~n74287 & ~n74288;
  assign n74290 = n73891 & ~n74289;
  assign n74291 = ~n74251 & n74285;
  assign n13991 = n74290 | ~n74291;
  assign n74293 = ~n73552 & n73888;
  assign n74294 = P2_P2_INSTQUEUE_REG_15__7_ & n73977;
  assign n74295 = P2_P2_INSTQUEUE_REG_14__7_ & n73979;
  assign n74296 = P2_P2_INSTQUEUE_REG_13__7_ & n73981;
  assign n74297 = P2_P2_INSTQUEUE_REG_12__7_ & n73983;
  assign n74298 = ~n74294 & ~n74295;
  assign n74299 = ~n74296 & n74298;
  assign n74300 = ~n74297 & n74299;
  assign n74301 = P2_P2_INSTQUEUE_REG_11__7_ & n73989;
  assign n74302 = P2_P2_INSTQUEUE_REG_10__7_ & n73991;
  assign n74303 = P2_P2_INSTQUEUE_REG_9__7_ & n73993;
  assign n74304 = P2_P2_INSTQUEUE_REG_8__7_ & n73995;
  assign n74305 = ~n74301 & ~n74302;
  assign n74306 = ~n74303 & n74305;
  assign n74307 = ~n74304 & n74306;
  assign n74308 = P2_P2_INSTQUEUE_REG_7__7_ & n74001;
  assign n74309 = P2_P2_INSTQUEUE_REG_6__7_ & n74003;
  assign n74310 = P2_P2_INSTQUEUE_REG_5__7_ & n74005;
  assign n74311 = P2_P2_INSTQUEUE_REG_4__7_ & n74007;
  assign n74312 = ~n74308 & ~n74309;
  assign n74313 = ~n74310 & n74312;
  assign n74314 = ~n74311 & n74313;
  assign n74315 = P2_P2_INSTQUEUE_REG_3__7_ & n74013;
  assign n74316 = P2_P2_INSTQUEUE_REG_2__7_ & n74015;
  assign n74317 = P2_P2_INSTQUEUE_REG_1__7_ & n74017;
  assign n74318 = P2_P2_INSTQUEUE_REG_0__7_ & n74019;
  assign n74319 = ~n74315 & ~n74316;
  assign n74320 = ~n74317 & n74319;
  assign n74321 = ~n74318 & n74320;
  assign n74322 = n74300 & n74307;
  assign n74323 = n74314 & n74322;
  assign n74324 = n74321 & n74323;
  assign n74325 = n73885 & ~n74324;
  assign n74326 = P2_P2_EAX_REG_15_ & ~n73884;
  assign n74327 = ~n74325 & ~n74326;
  assign n74328 = P2_P2_EAX_REG_13_ & P2_P2_EAX_REG_14_;
  assign n74329 = n74244 & n74328;
  assign n74330 = P2_P2_EAX_REG_15_ & ~n74329;
  assign n74331 = ~P2_P2_EAX_REG_15_ & n74329;
  assign n74332 = ~n74330 & ~n74331;
  assign n74333 = n73891 & ~n74332;
  assign n74334 = ~n74293 & n74327;
  assign n13996 = n74333 | ~n74334;
  assign n74336 = ~n67722 & n73887;
  assign n74337 = ~n68545 & n74336;
  assign n74338 = n67691 & n73887;
  assign n74339 = ~n68559 & n74338;
  assign n74340 = P2_P2_EAX_REG_16_ & ~n73884;
  assign n74341 = P2_P2_INSTQUEUERD_ADDR_REG_2_ & ~n67647;
  assign n74342 = ~P2_P2_INSTQUEUERD_ADDR_REG_3_ & n74341;
  assign n74343 = P2_P2_INSTQUEUERD_ADDR_REG_3_ & ~n74341;
  assign n74344 = ~n74342 & ~n74343;
  assign n74345 = ~n67648 & ~n74341;
  assign n74346 = n74344 & n74345;
  assign n74347 = n70000 & n74346;
  assign n74348 = P2_P2_INSTQUEUE_REG_7__0_ & n74347;
  assign n74349 = n69997 & n74346;
  assign n74350 = P2_P2_INSTQUEUE_REG_6__0_ & n74349;
  assign n74351 = n70006 & n74346;
  assign n74352 = P2_P2_INSTQUEUE_REG_5__0_ & n74351;
  assign n74353 = n70003 & n74346;
  assign n74354 = P2_P2_INSTQUEUE_REG_4__0_ & n74353;
  assign n74355 = ~n74348 & ~n74350;
  assign n74356 = ~n74352 & n74355;
  assign n74357 = ~n74354 & n74356;
  assign n74358 = n74344 & ~n74345;
  assign n74359 = n70000 & n74358;
  assign n74360 = P2_P2_INSTQUEUE_REG_3__0_ & n74359;
  assign n74361 = n69997 & n74358;
  assign n74362 = P2_P2_INSTQUEUE_REG_2__0_ & n74361;
  assign n74363 = n70006 & n74358;
  assign n74364 = P2_P2_INSTQUEUE_REG_1__0_ & n74363;
  assign n74365 = n70003 & n74358;
  assign n74366 = P2_P2_INSTQUEUE_REG_0__0_ & n74365;
  assign n74367 = ~n74360 & ~n74362;
  assign n74368 = ~n74364 & n74367;
  assign n74369 = ~n74366 & n74368;
  assign n74370 = ~n74344 & n74345;
  assign n74371 = n70000 & n74370;
  assign n74372 = P2_P2_INSTQUEUE_REG_15__0_ & n74371;
  assign n74373 = n69997 & n74370;
  assign n74374 = P2_P2_INSTQUEUE_REG_14__0_ & n74373;
  assign n74375 = n70006 & n74370;
  assign n74376 = P2_P2_INSTQUEUE_REG_13__0_ & n74375;
  assign n74377 = n70003 & n74370;
  assign n74378 = P2_P2_INSTQUEUE_REG_12__0_ & n74377;
  assign n74379 = ~n74372 & ~n74374;
  assign n74380 = ~n74376 & n74379;
  assign n74381 = ~n74378 & n74380;
  assign n74382 = ~n74344 & ~n74345;
  assign n74383 = n70000 & n74382;
  assign n74384 = P2_P2_INSTQUEUE_REG_11__0_ & n74383;
  assign n74385 = n69997 & n74382;
  assign n74386 = P2_P2_INSTQUEUE_REG_10__0_ & n74385;
  assign n74387 = n70006 & n74382;
  assign n74388 = P2_P2_INSTQUEUE_REG_9__0_ & n74387;
  assign n74389 = n70003 & n74382;
  assign n74390 = P2_P2_INSTQUEUE_REG_8__0_ & n74389;
  assign n74391 = ~n74384 & ~n74386;
  assign n74392 = ~n74388 & n74391;
  assign n74393 = ~n74390 & n74392;
  assign n74394 = n74357 & n74369;
  assign n74395 = n74381 & n74394;
  assign n74396 = n74393 & n74395;
  assign n74397 = n73885 & ~n74396;
  assign n74398 = ~n74340 & ~n74397;
  assign n74399 = P2_P2_EAX_REG_15_ & n74329;
  assign n74400 = ~P2_P2_EAX_REG_16_ & n74399;
  assign n74401 = P2_P2_EAX_REG_16_ & ~n74399;
  assign n74402 = ~n74400 & ~n74401;
  assign n74403 = n73891 & ~n74402;
  assign n74404 = ~n74337 & ~n74339;
  assign n74405 = n74398 & n74404;
  assign n14001 = n74403 | ~n74405;
  assign n74407 = ~n68523 & n74336;
  assign n74408 = ~n68537 & n74338;
  assign n74409 = P2_P2_EAX_REG_17_ & ~n73884;
  assign n74410 = P2_P2_INSTQUEUE_REG_7__1_ & n74347;
  assign n74411 = P2_P2_INSTQUEUE_REG_6__1_ & n74349;
  assign n74412 = P2_P2_INSTQUEUE_REG_5__1_ & n74351;
  assign n74413 = P2_P2_INSTQUEUE_REG_4__1_ & n74353;
  assign n74414 = ~n74410 & ~n74411;
  assign n74415 = ~n74412 & n74414;
  assign n74416 = ~n74413 & n74415;
  assign n74417 = P2_P2_INSTQUEUE_REG_3__1_ & n74359;
  assign n74418 = P2_P2_INSTQUEUE_REG_2__1_ & n74361;
  assign n74419 = P2_P2_INSTQUEUE_REG_1__1_ & n74363;
  assign n74420 = P2_P2_INSTQUEUE_REG_0__1_ & n74365;
  assign n74421 = ~n74417 & ~n74418;
  assign n74422 = ~n74419 & n74421;
  assign n74423 = ~n74420 & n74422;
  assign n74424 = P2_P2_INSTQUEUE_REG_15__1_ & n74371;
  assign n74425 = P2_P2_INSTQUEUE_REG_14__1_ & n74373;
  assign n74426 = P2_P2_INSTQUEUE_REG_13__1_ & n74375;
  assign n74427 = P2_P2_INSTQUEUE_REG_12__1_ & n74377;
  assign n74428 = ~n74424 & ~n74425;
  assign n74429 = ~n74426 & n74428;
  assign n74430 = ~n74427 & n74429;
  assign n74431 = P2_P2_INSTQUEUE_REG_11__1_ & n74383;
  assign n74432 = P2_P2_INSTQUEUE_REG_10__1_ & n74385;
  assign n74433 = P2_P2_INSTQUEUE_REG_9__1_ & n74387;
  assign n74434 = P2_P2_INSTQUEUE_REG_8__1_ & n74389;
  assign n74435 = ~n74431 & ~n74432;
  assign n74436 = ~n74433 & n74435;
  assign n74437 = ~n74434 & n74436;
  assign n74438 = n74416 & n74423;
  assign n74439 = n74430 & n74438;
  assign n74440 = n74437 & n74439;
  assign n74441 = n73885 & ~n74440;
  assign n74442 = ~n74409 & ~n74441;
  assign n74443 = P2_P2_EAX_REG_15_ & P2_P2_EAX_REG_16_;
  assign n74444 = n74329 & n74443;
  assign n74445 = P2_P2_EAX_REG_17_ & ~n74444;
  assign n74446 = ~P2_P2_EAX_REG_17_ & n74444;
  assign n74447 = ~n74445 & ~n74446;
  assign n74448 = n73891 & ~n74447;
  assign n74449 = ~n74407 & ~n74408;
  assign n74450 = n74442 & n74449;
  assign n14006 = n74448 | ~n74450;
  assign n74452 = ~n68501 & n74336;
  assign n74453 = ~n68515 & n74338;
  assign n74454 = P2_P2_EAX_REG_18_ & ~n73884;
  assign n74455 = P2_P2_INSTQUEUE_REG_7__2_ & n74347;
  assign n74456 = P2_P2_INSTQUEUE_REG_6__2_ & n74349;
  assign n74457 = P2_P2_INSTQUEUE_REG_5__2_ & n74351;
  assign n74458 = P2_P2_INSTQUEUE_REG_4__2_ & n74353;
  assign n74459 = ~n74455 & ~n74456;
  assign n74460 = ~n74457 & n74459;
  assign n74461 = ~n74458 & n74460;
  assign n74462 = P2_P2_INSTQUEUE_REG_3__2_ & n74359;
  assign n74463 = P2_P2_INSTQUEUE_REG_2__2_ & n74361;
  assign n74464 = P2_P2_INSTQUEUE_REG_1__2_ & n74363;
  assign n74465 = P2_P2_INSTQUEUE_REG_0__2_ & n74365;
  assign n74466 = ~n74462 & ~n74463;
  assign n74467 = ~n74464 & n74466;
  assign n74468 = ~n74465 & n74467;
  assign n74469 = P2_P2_INSTQUEUE_REG_15__2_ & n74371;
  assign n74470 = P2_P2_INSTQUEUE_REG_14__2_ & n74373;
  assign n74471 = P2_P2_INSTQUEUE_REG_13__2_ & n74375;
  assign n74472 = P2_P2_INSTQUEUE_REG_12__2_ & n74377;
  assign n74473 = ~n74469 & ~n74470;
  assign n74474 = ~n74471 & n74473;
  assign n74475 = ~n74472 & n74474;
  assign n74476 = P2_P2_INSTQUEUE_REG_11__2_ & n74383;
  assign n74477 = P2_P2_INSTQUEUE_REG_10__2_ & n74385;
  assign n74478 = P2_P2_INSTQUEUE_REG_9__2_ & n74387;
  assign n74479 = P2_P2_INSTQUEUE_REG_8__2_ & n74389;
  assign n74480 = ~n74476 & ~n74477;
  assign n74481 = ~n74478 & n74480;
  assign n74482 = ~n74479 & n74481;
  assign n74483 = n74461 & n74468;
  assign n74484 = n74475 & n74483;
  assign n74485 = n74482 & n74484;
  assign n74486 = n73885 & ~n74485;
  assign n74487 = ~n74454 & ~n74486;
  assign n74488 = P2_P2_EAX_REG_17_ & n74444;
  assign n74489 = ~P2_P2_EAX_REG_18_ & n74488;
  assign n74490 = P2_P2_EAX_REG_18_ & ~n74488;
  assign n74491 = ~n74489 & ~n74490;
  assign n74492 = n73891 & ~n74491;
  assign n74493 = ~n74452 & ~n74453;
  assign n74494 = n74487 & n74493;
  assign n14011 = n74492 | ~n74494;
  assign n74496 = ~n68479 & n74336;
  assign n74497 = ~n68493 & n74338;
  assign n74498 = P2_P2_EAX_REG_19_ & ~n73884;
  assign n74499 = P2_P2_INSTQUEUE_REG_7__3_ & n74347;
  assign n74500 = P2_P2_INSTQUEUE_REG_6__3_ & n74349;
  assign n74501 = P2_P2_INSTQUEUE_REG_5__3_ & n74351;
  assign n74502 = P2_P2_INSTQUEUE_REG_4__3_ & n74353;
  assign n74503 = ~n74499 & ~n74500;
  assign n74504 = ~n74501 & n74503;
  assign n74505 = ~n74502 & n74504;
  assign n74506 = P2_P2_INSTQUEUE_REG_3__3_ & n74359;
  assign n74507 = P2_P2_INSTQUEUE_REG_2__3_ & n74361;
  assign n74508 = P2_P2_INSTQUEUE_REG_1__3_ & n74363;
  assign n74509 = P2_P2_INSTQUEUE_REG_0__3_ & n74365;
  assign n74510 = ~n74506 & ~n74507;
  assign n74511 = ~n74508 & n74510;
  assign n74512 = ~n74509 & n74511;
  assign n74513 = P2_P2_INSTQUEUE_REG_15__3_ & n74371;
  assign n74514 = P2_P2_INSTQUEUE_REG_14__3_ & n74373;
  assign n74515 = P2_P2_INSTQUEUE_REG_13__3_ & n74375;
  assign n74516 = P2_P2_INSTQUEUE_REG_12__3_ & n74377;
  assign n74517 = ~n74513 & ~n74514;
  assign n74518 = ~n74515 & n74517;
  assign n74519 = ~n74516 & n74518;
  assign n74520 = P2_P2_INSTQUEUE_REG_11__3_ & n74383;
  assign n74521 = P2_P2_INSTQUEUE_REG_10__3_ & n74385;
  assign n74522 = P2_P2_INSTQUEUE_REG_9__3_ & n74387;
  assign n74523 = P2_P2_INSTQUEUE_REG_8__3_ & n74389;
  assign n74524 = ~n74520 & ~n74521;
  assign n74525 = ~n74522 & n74524;
  assign n74526 = ~n74523 & n74525;
  assign n74527 = n74505 & n74512;
  assign n74528 = n74519 & n74527;
  assign n74529 = n74526 & n74528;
  assign n74530 = n73885 & ~n74529;
  assign n74531 = ~n74498 & ~n74530;
  assign n74532 = P2_P2_EAX_REG_17_ & P2_P2_EAX_REG_18_;
  assign n74533 = n74444 & n74532;
  assign n74534 = P2_P2_EAX_REG_19_ & ~n74533;
  assign n74535 = ~P2_P2_EAX_REG_19_ & n74533;
  assign n74536 = ~n74534 & ~n74535;
  assign n74537 = n73891 & ~n74536;
  assign n74538 = ~n74496 & ~n74497;
  assign n74539 = n74531 & n74538;
  assign n14016 = n74537 | ~n74539;
  assign n74541 = ~n68457 & n74336;
  assign n74542 = ~n68471 & n74338;
  assign n74543 = P2_P2_EAX_REG_20_ & ~n73884;
  assign n74544 = P2_P2_INSTQUEUE_REG_7__4_ & n74347;
  assign n74545 = P2_P2_INSTQUEUE_REG_6__4_ & n74349;
  assign n74546 = P2_P2_INSTQUEUE_REG_5__4_ & n74351;
  assign n74547 = P2_P2_INSTQUEUE_REG_4__4_ & n74353;
  assign n74548 = ~n74544 & ~n74545;
  assign n74549 = ~n74546 & n74548;
  assign n74550 = ~n74547 & n74549;
  assign n74551 = P2_P2_INSTQUEUE_REG_3__4_ & n74359;
  assign n74552 = P2_P2_INSTQUEUE_REG_2__4_ & n74361;
  assign n74553 = P2_P2_INSTQUEUE_REG_1__4_ & n74363;
  assign n74554 = P2_P2_INSTQUEUE_REG_0__4_ & n74365;
  assign n74555 = ~n74551 & ~n74552;
  assign n74556 = ~n74553 & n74555;
  assign n74557 = ~n74554 & n74556;
  assign n74558 = P2_P2_INSTQUEUE_REG_15__4_ & n74371;
  assign n74559 = P2_P2_INSTQUEUE_REG_14__4_ & n74373;
  assign n74560 = P2_P2_INSTQUEUE_REG_13__4_ & n74375;
  assign n74561 = P2_P2_INSTQUEUE_REG_12__4_ & n74377;
  assign n74562 = ~n74558 & ~n74559;
  assign n74563 = ~n74560 & n74562;
  assign n74564 = ~n74561 & n74563;
  assign n74565 = P2_P2_INSTQUEUE_REG_11__4_ & n74383;
  assign n74566 = P2_P2_INSTQUEUE_REG_10__4_ & n74385;
  assign n74567 = P2_P2_INSTQUEUE_REG_9__4_ & n74387;
  assign n74568 = P2_P2_INSTQUEUE_REG_8__4_ & n74389;
  assign n74569 = ~n74565 & ~n74566;
  assign n74570 = ~n74567 & n74569;
  assign n74571 = ~n74568 & n74570;
  assign n74572 = n74550 & n74557;
  assign n74573 = n74564 & n74572;
  assign n74574 = n74571 & n74573;
  assign n74575 = n73885 & ~n74574;
  assign n74576 = ~n74543 & ~n74575;
  assign n74577 = P2_P2_EAX_REG_19_ & n74533;
  assign n74578 = ~P2_P2_EAX_REG_20_ & n74577;
  assign n74579 = P2_P2_EAX_REG_20_ & ~n74577;
  assign n74580 = ~n74578 & ~n74579;
  assign n74581 = n73891 & ~n74580;
  assign n74582 = ~n74541 & ~n74542;
  assign n74583 = n74576 & n74582;
  assign n14021 = n74581 | ~n74583;
  assign n74585 = ~n68435 & n74336;
  assign n74586 = ~n68449 & n74338;
  assign n74587 = P2_P2_EAX_REG_21_ & ~n73884;
  assign n74588 = P2_P2_INSTQUEUE_REG_7__5_ & n74347;
  assign n74589 = P2_P2_INSTQUEUE_REG_6__5_ & n74349;
  assign n74590 = P2_P2_INSTQUEUE_REG_5__5_ & n74351;
  assign n74591 = P2_P2_INSTQUEUE_REG_4__5_ & n74353;
  assign n74592 = ~n74588 & ~n74589;
  assign n74593 = ~n74590 & n74592;
  assign n74594 = ~n74591 & n74593;
  assign n74595 = P2_P2_INSTQUEUE_REG_3__5_ & n74359;
  assign n74596 = P2_P2_INSTQUEUE_REG_2__5_ & n74361;
  assign n74597 = P2_P2_INSTQUEUE_REG_1__5_ & n74363;
  assign n74598 = P2_P2_INSTQUEUE_REG_0__5_ & n74365;
  assign n74599 = ~n74595 & ~n74596;
  assign n74600 = ~n74597 & n74599;
  assign n74601 = ~n74598 & n74600;
  assign n74602 = P2_P2_INSTQUEUE_REG_15__5_ & n74371;
  assign n74603 = P2_P2_INSTQUEUE_REG_14__5_ & n74373;
  assign n74604 = P2_P2_INSTQUEUE_REG_13__5_ & n74375;
  assign n74605 = P2_P2_INSTQUEUE_REG_12__5_ & n74377;
  assign n74606 = ~n74602 & ~n74603;
  assign n74607 = ~n74604 & n74606;
  assign n74608 = ~n74605 & n74607;
  assign n74609 = P2_P2_INSTQUEUE_REG_11__5_ & n74383;
  assign n74610 = P2_P2_INSTQUEUE_REG_10__5_ & n74385;
  assign n74611 = P2_P2_INSTQUEUE_REG_9__5_ & n74387;
  assign n74612 = P2_P2_INSTQUEUE_REG_8__5_ & n74389;
  assign n74613 = ~n74609 & ~n74610;
  assign n74614 = ~n74611 & n74613;
  assign n74615 = ~n74612 & n74614;
  assign n74616 = n74594 & n74601;
  assign n74617 = n74608 & n74616;
  assign n74618 = n74615 & n74617;
  assign n74619 = n73885 & ~n74618;
  assign n74620 = ~n74587 & ~n74619;
  assign n74621 = P2_P2_EAX_REG_19_ & P2_P2_EAX_REG_20_;
  assign n74622 = n74533 & n74621;
  assign n74623 = P2_P2_EAX_REG_21_ & ~n74622;
  assign n74624 = ~P2_P2_EAX_REG_21_ & n74622;
  assign n74625 = ~n74623 & ~n74624;
  assign n74626 = n73891 & ~n74625;
  assign n74627 = ~n74585 & ~n74586;
  assign n74628 = n74620 & n74627;
  assign n14026 = n74626 | ~n74628;
  assign n74630 = ~n68413 & n74336;
  assign n74631 = ~n68427 & n74338;
  assign n74632 = P2_P2_EAX_REG_22_ & ~n73884;
  assign n74633 = P2_P2_INSTQUEUE_REG_7__6_ & n74347;
  assign n74634 = P2_P2_INSTQUEUE_REG_6__6_ & n74349;
  assign n74635 = P2_P2_INSTQUEUE_REG_5__6_ & n74351;
  assign n74636 = P2_P2_INSTQUEUE_REG_4__6_ & n74353;
  assign n74637 = ~n74633 & ~n74634;
  assign n74638 = ~n74635 & n74637;
  assign n74639 = ~n74636 & n74638;
  assign n74640 = P2_P2_INSTQUEUE_REG_3__6_ & n74359;
  assign n74641 = P2_P2_INSTQUEUE_REG_2__6_ & n74361;
  assign n74642 = P2_P2_INSTQUEUE_REG_1__6_ & n74363;
  assign n74643 = P2_P2_INSTQUEUE_REG_0__6_ & n74365;
  assign n74644 = ~n74640 & ~n74641;
  assign n74645 = ~n74642 & n74644;
  assign n74646 = ~n74643 & n74645;
  assign n74647 = P2_P2_INSTQUEUE_REG_15__6_ & n74371;
  assign n74648 = P2_P2_INSTQUEUE_REG_14__6_ & n74373;
  assign n74649 = P2_P2_INSTQUEUE_REG_13__6_ & n74375;
  assign n74650 = P2_P2_INSTQUEUE_REG_12__6_ & n74377;
  assign n74651 = ~n74647 & ~n74648;
  assign n74652 = ~n74649 & n74651;
  assign n74653 = ~n74650 & n74652;
  assign n74654 = P2_P2_INSTQUEUE_REG_11__6_ & n74383;
  assign n74655 = P2_P2_INSTQUEUE_REG_10__6_ & n74385;
  assign n74656 = P2_P2_INSTQUEUE_REG_9__6_ & n74387;
  assign n74657 = P2_P2_INSTQUEUE_REG_8__6_ & n74389;
  assign n74658 = ~n74654 & ~n74655;
  assign n74659 = ~n74656 & n74658;
  assign n74660 = ~n74657 & n74659;
  assign n74661 = n74639 & n74646;
  assign n74662 = n74653 & n74661;
  assign n74663 = n74660 & n74662;
  assign n74664 = n73885 & ~n74663;
  assign n74665 = ~n74632 & ~n74664;
  assign n74666 = P2_P2_EAX_REG_21_ & n74622;
  assign n74667 = ~P2_P2_EAX_REG_22_ & n74666;
  assign n74668 = P2_P2_EAX_REG_22_ & ~n74666;
  assign n74669 = ~n74667 & ~n74668;
  assign n74670 = n73891 & ~n74669;
  assign n74671 = ~n74630 & ~n74631;
  assign n74672 = n74665 & n74671;
  assign n14031 = n74670 | ~n74672;
  assign n74674 = ~n68385 & n74336;
  assign n74675 = ~n68405 & n74338;
  assign n74676 = P2_P2_EAX_REG_23_ & ~n73884;
  assign n74677 = P2_P2_INSTQUEUERD_ADDR_REG_3_ & ~P2_P2_INSTQUEUERD_ADDR_REG_2_;
  assign n74678 = ~n67664 & ~n74677;
  assign n74679 = n67635 & n74678;
  assign n74680 = P2_P2_INSTQUEUE_REG_7__0_ & n74679;
  assign n74681 = n67639 & n74678;
  assign n74682 = P2_P2_INSTQUEUE_REG_6__0_ & n74681;
  assign n74683 = n67644 & n74678;
  assign n74684 = P2_P2_INSTQUEUE_REG_5__0_ & n74683;
  assign n74685 = n67648 & n74678;
  assign n74686 = P2_P2_INSTQUEUE_REG_4__0_ & n74685;
  assign n74687 = ~n74680 & ~n74682;
  assign n74688 = ~n74684 & n74687;
  assign n74689 = ~n74686 & n74688;
  assign n74690 = P2_P2_INSTQUEUERD_ADDR_REG_2_ & n74678;
  assign n74691 = n67634 & n74690;
  assign n74692 = P2_P2_INSTQUEUE_REG_3__0_ & n74691;
  assign n74693 = n67638 & n74690;
  assign n74694 = P2_P2_INSTQUEUE_REG_2__0_ & n74693;
  assign n74695 = n67643 & n74690;
  assign n74696 = P2_P2_INSTQUEUE_REG_1__0_ & n74695;
  assign n74697 = n67647 & n74690;
  assign n74698 = P2_P2_INSTQUEUE_REG_0__0_ & n74697;
  assign n74699 = ~n74692 & ~n74694;
  assign n74700 = ~n74696 & n74699;
  assign n74701 = ~n74698 & n74700;
  assign n74702 = n67635 & ~n74678;
  assign n74703 = P2_P2_INSTQUEUE_REG_15__0_ & n74702;
  assign n74704 = n67639 & ~n74678;
  assign n74705 = P2_P2_INSTQUEUE_REG_14__0_ & n74704;
  assign n74706 = n67644 & ~n74678;
  assign n74707 = P2_P2_INSTQUEUE_REG_13__0_ & n74706;
  assign n74708 = n67648 & ~n74678;
  assign n74709 = P2_P2_INSTQUEUE_REG_12__0_ & n74708;
  assign n74710 = ~n74703 & ~n74705;
  assign n74711 = ~n74707 & n74710;
  assign n74712 = ~n74709 & n74711;
  assign n74713 = P2_P2_INSTQUEUERD_ADDR_REG_2_ & ~n74678;
  assign n74714 = n67634 & n74713;
  assign n74715 = P2_P2_INSTQUEUE_REG_11__0_ & n74714;
  assign n74716 = n67638 & n74713;
  assign n74717 = P2_P2_INSTQUEUE_REG_10__0_ & n74716;
  assign n74718 = n67643 & n74713;
  assign n74719 = P2_P2_INSTQUEUE_REG_9__0_ & n74718;
  assign n74720 = n67647 & n74713;
  assign n74721 = P2_P2_INSTQUEUE_REG_8__0_ & n74720;
  assign n74722 = ~n74715 & ~n74717;
  assign n74723 = ~n74719 & n74722;
  assign n74724 = ~n74721 & n74723;
  assign n74725 = n74689 & n74701;
  assign n74726 = n74712 & n74725;
  assign n74727 = n74724 & n74726;
  assign n74728 = P2_P2_INSTQUEUE_REG_7__7_ & n74347;
  assign n74729 = P2_P2_INSTQUEUE_REG_6__7_ & n74349;
  assign n74730 = P2_P2_INSTQUEUE_REG_5__7_ & n74351;
  assign n74731 = P2_P2_INSTQUEUE_REG_4__7_ & n74353;
  assign n74732 = ~n74728 & ~n74729;
  assign n74733 = ~n74730 & n74732;
  assign n74734 = ~n74731 & n74733;
  assign n74735 = P2_P2_INSTQUEUE_REG_3__7_ & n74359;
  assign n74736 = P2_P2_INSTQUEUE_REG_2__7_ & n74361;
  assign n74737 = P2_P2_INSTQUEUE_REG_1__7_ & n74363;
  assign n74738 = P2_P2_INSTQUEUE_REG_0__7_ & n74365;
  assign n74739 = ~n74735 & ~n74736;
  assign n74740 = ~n74737 & n74739;
  assign n74741 = ~n74738 & n74740;
  assign n74742 = P2_P2_INSTQUEUE_REG_15__7_ & n74371;
  assign n74743 = P2_P2_INSTQUEUE_REG_14__7_ & n74373;
  assign n74744 = P2_P2_INSTQUEUE_REG_13__7_ & n74375;
  assign n74745 = P2_P2_INSTQUEUE_REG_12__7_ & n74377;
  assign n74746 = ~n74742 & ~n74743;
  assign n74747 = ~n74744 & n74746;
  assign n74748 = ~n74745 & n74747;
  assign n74749 = P2_P2_INSTQUEUE_REG_11__7_ & n74383;
  assign n74750 = P2_P2_INSTQUEUE_REG_10__7_ & n74385;
  assign n74751 = P2_P2_INSTQUEUE_REG_9__7_ & n74387;
  assign n74752 = P2_P2_INSTQUEUE_REG_8__7_ & n74389;
  assign n74753 = ~n74749 & ~n74750;
  assign n74754 = ~n74751 & n74753;
  assign n74755 = ~n74752 & n74754;
  assign n74756 = n74734 & n74741;
  assign n74757 = n74748 & n74756;
  assign n74758 = n74755 & n74757;
  assign n74759 = ~n74727 & n74758;
  assign n74760 = n74727 & ~n74758;
  assign n74761 = ~n74759 & ~n74760;
  assign n74762 = n73885 & ~n74761;
  assign n74763 = ~n74676 & ~n74762;
  assign n74764 = P2_P2_EAX_REG_21_ & P2_P2_EAX_REG_22_;
  assign n74765 = n74622 & n74764;
  assign n74766 = P2_P2_EAX_REG_23_ & ~n74765;
  assign n74767 = ~P2_P2_EAX_REG_23_ & n74765;
  assign n74768 = ~n74766 & ~n74767;
  assign n74769 = n73891 & ~n74768;
  assign n74770 = ~n74674 & ~n74675;
  assign n74771 = n74763 & n74770;
  assign n14036 = n74769 | ~n74771;
  assign n74773 = ~n68553 & n74336;
  assign n74774 = ~n73614 & n74338;
  assign n74775 = P2_P2_EAX_REG_24_ & ~n73884;
  assign n74776 = ~n74727 & ~n74758;
  assign n74777 = P2_P2_INSTQUEUE_REG_7__1_ & n74679;
  assign n74778 = P2_P2_INSTQUEUE_REG_6__1_ & n74681;
  assign n74779 = P2_P2_INSTQUEUE_REG_5__1_ & n74683;
  assign n74780 = P2_P2_INSTQUEUE_REG_4__1_ & n74685;
  assign n74781 = ~n74777 & ~n74778;
  assign n74782 = ~n74779 & n74781;
  assign n74783 = ~n74780 & n74782;
  assign n74784 = P2_P2_INSTQUEUE_REG_3__1_ & n74691;
  assign n74785 = P2_P2_INSTQUEUE_REG_2__1_ & n74693;
  assign n74786 = P2_P2_INSTQUEUE_REG_1__1_ & n74695;
  assign n74787 = P2_P2_INSTQUEUE_REG_0__1_ & n74697;
  assign n74788 = ~n74784 & ~n74785;
  assign n74789 = ~n74786 & n74788;
  assign n74790 = ~n74787 & n74789;
  assign n74791 = P2_P2_INSTQUEUE_REG_15__1_ & n74702;
  assign n74792 = P2_P2_INSTQUEUE_REG_14__1_ & n74704;
  assign n74793 = P2_P2_INSTQUEUE_REG_13__1_ & n74706;
  assign n74794 = P2_P2_INSTQUEUE_REG_12__1_ & n74708;
  assign n74795 = ~n74791 & ~n74792;
  assign n74796 = ~n74793 & n74795;
  assign n74797 = ~n74794 & n74796;
  assign n74798 = P2_P2_INSTQUEUE_REG_11__1_ & n74714;
  assign n74799 = P2_P2_INSTQUEUE_REG_10__1_ & n74716;
  assign n74800 = P2_P2_INSTQUEUE_REG_9__1_ & n74718;
  assign n74801 = P2_P2_INSTQUEUE_REG_8__1_ & n74720;
  assign n74802 = ~n74798 & ~n74799;
  assign n74803 = ~n74800 & n74802;
  assign n74804 = ~n74801 & n74803;
  assign n74805 = n74783 & n74790;
  assign n74806 = n74797 & n74805;
  assign n74807 = n74804 & n74806;
  assign n74808 = n74776 & n74807;
  assign n74809 = ~n74776 & ~n74807;
  assign n74810 = ~n74808 & ~n74809;
  assign n74811 = n73885 & ~n74810;
  assign n74812 = ~n74775 & ~n74811;
  assign n74813 = P2_P2_EAX_REG_23_ & n74765;
  assign n74814 = ~P2_P2_EAX_REG_24_ & n74813;
  assign n74815 = P2_P2_EAX_REG_24_ & ~n74813;
  assign n74816 = ~n74814 & ~n74815;
  assign n74817 = n73891 & ~n74816;
  assign n74818 = ~n74773 & ~n74774;
  assign n74819 = n74812 & n74818;
  assign n14041 = n74817 | ~n74819;
  assign n74821 = ~n68531 & n74336;
  assign n74822 = ~n73606 & n74338;
  assign n74823 = P2_P2_EAX_REG_25_ & ~n73884;
  assign n74824 = n74776 & ~n74807;
  assign n74825 = P2_P2_INSTQUEUE_REG_7__2_ & n74679;
  assign n74826 = P2_P2_INSTQUEUE_REG_6__2_ & n74681;
  assign n74827 = P2_P2_INSTQUEUE_REG_5__2_ & n74683;
  assign n74828 = P2_P2_INSTQUEUE_REG_4__2_ & n74685;
  assign n74829 = ~n74825 & ~n74826;
  assign n74830 = ~n74827 & n74829;
  assign n74831 = ~n74828 & n74830;
  assign n74832 = P2_P2_INSTQUEUE_REG_3__2_ & n74691;
  assign n74833 = P2_P2_INSTQUEUE_REG_2__2_ & n74693;
  assign n74834 = P2_P2_INSTQUEUE_REG_1__2_ & n74695;
  assign n74835 = P2_P2_INSTQUEUE_REG_0__2_ & n74697;
  assign n74836 = ~n74832 & ~n74833;
  assign n74837 = ~n74834 & n74836;
  assign n74838 = ~n74835 & n74837;
  assign n74839 = P2_P2_INSTQUEUE_REG_15__2_ & n74702;
  assign n74840 = P2_P2_INSTQUEUE_REG_14__2_ & n74704;
  assign n74841 = P2_P2_INSTQUEUE_REG_13__2_ & n74706;
  assign n74842 = P2_P2_INSTQUEUE_REG_12__2_ & n74708;
  assign n74843 = ~n74839 & ~n74840;
  assign n74844 = ~n74841 & n74843;
  assign n74845 = ~n74842 & n74844;
  assign n74846 = P2_P2_INSTQUEUE_REG_11__2_ & n74714;
  assign n74847 = P2_P2_INSTQUEUE_REG_10__2_ & n74716;
  assign n74848 = P2_P2_INSTQUEUE_REG_9__2_ & n74718;
  assign n74849 = P2_P2_INSTQUEUE_REG_8__2_ & n74720;
  assign n74850 = ~n74846 & ~n74847;
  assign n74851 = ~n74848 & n74850;
  assign n74852 = ~n74849 & n74851;
  assign n74853 = n74831 & n74838;
  assign n74854 = n74845 & n74853;
  assign n74855 = n74852 & n74854;
  assign n74856 = n74824 & n74855;
  assign n74857 = ~n74824 & ~n74855;
  assign n74858 = ~n74856 & ~n74857;
  assign n74859 = n73885 & ~n74858;
  assign n74860 = ~n74823 & ~n74859;
  assign n74861 = P2_P2_EAX_REG_23_ & P2_P2_EAX_REG_24_;
  assign n74862 = n74765 & n74861;
  assign n74863 = P2_P2_EAX_REG_25_ & ~n74862;
  assign n74864 = ~P2_P2_EAX_REG_25_ & n74862;
  assign n74865 = ~n74863 & ~n74864;
  assign n74866 = n73891 & ~n74865;
  assign n74867 = ~n74821 & ~n74822;
  assign n74868 = n74860 & n74867;
  assign n14046 = n74866 | ~n74868;
  assign n74870 = ~n68509 & n74336;
  assign n74871 = ~n73598 & n74338;
  assign n74872 = P2_P2_EAX_REG_26_ & ~n73884;
  assign n74873 = n74824 & ~n74855;
  assign n74874 = P2_P2_INSTQUEUE_REG_7__3_ & n74679;
  assign n74875 = P2_P2_INSTQUEUE_REG_6__3_ & n74681;
  assign n74876 = P2_P2_INSTQUEUE_REG_5__3_ & n74683;
  assign n74877 = P2_P2_INSTQUEUE_REG_4__3_ & n74685;
  assign n74878 = ~n74874 & ~n74875;
  assign n74879 = ~n74876 & n74878;
  assign n74880 = ~n74877 & n74879;
  assign n74881 = P2_P2_INSTQUEUE_REG_3__3_ & n74691;
  assign n74882 = P2_P2_INSTQUEUE_REG_2__3_ & n74693;
  assign n74883 = P2_P2_INSTQUEUE_REG_1__3_ & n74695;
  assign n74884 = P2_P2_INSTQUEUE_REG_0__3_ & n74697;
  assign n74885 = ~n74881 & ~n74882;
  assign n74886 = ~n74883 & n74885;
  assign n74887 = ~n74884 & n74886;
  assign n74888 = P2_P2_INSTQUEUE_REG_15__3_ & n74702;
  assign n74889 = P2_P2_INSTQUEUE_REG_14__3_ & n74704;
  assign n74890 = P2_P2_INSTQUEUE_REG_13__3_ & n74706;
  assign n74891 = P2_P2_INSTQUEUE_REG_12__3_ & n74708;
  assign n74892 = ~n74888 & ~n74889;
  assign n74893 = ~n74890 & n74892;
  assign n74894 = ~n74891 & n74893;
  assign n74895 = P2_P2_INSTQUEUE_REG_11__3_ & n74714;
  assign n74896 = P2_P2_INSTQUEUE_REG_10__3_ & n74716;
  assign n74897 = P2_P2_INSTQUEUE_REG_9__3_ & n74718;
  assign n74898 = P2_P2_INSTQUEUE_REG_8__3_ & n74720;
  assign n74899 = ~n74895 & ~n74896;
  assign n74900 = ~n74897 & n74899;
  assign n74901 = ~n74898 & n74900;
  assign n74902 = n74880 & n74887;
  assign n74903 = n74894 & n74902;
  assign n74904 = n74901 & n74903;
  assign n74905 = n74873 & n74904;
  assign n74906 = ~n74873 & ~n74904;
  assign n74907 = ~n74905 & ~n74906;
  assign n74908 = n73885 & ~n74907;
  assign n74909 = ~n74872 & ~n74908;
  assign n74910 = P2_P2_EAX_REG_25_ & n74862;
  assign n74911 = ~P2_P2_EAX_REG_26_ & n74910;
  assign n74912 = P2_P2_EAX_REG_26_ & ~n74910;
  assign n74913 = ~n74911 & ~n74912;
  assign n74914 = n73891 & ~n74913;
  assign n74915 = ~n74870 & ~n74871;
  assign n74916 = n74909 & n74915;
  assign n14051 = n74914 | ~n74916;
  assign n74918 = ~n68487 & n74336;
  assign n74919 = ~n73590 & n74338;
  assign n74920 = P2_P2_EAX_REG_27_ & ~n73884;
  assign n74921 = n74873 & ~n74904;
  assign n74922 = P2_P2_INSTQUEUE_REG_7__4_ & n74679;
  assign n74923 = P2_P2_INSTQUEUE_REG_6__4_ & n74681;
  assign n74924 = P2_P2_INSTQUEUE_REG_5__4_ & n74683;
  assign n74925 = P2_P2_INSTQUEUE_REG_4__4_ & n74685;
  assign n74926 = ~n74922 & ~n74923;
  assign n74927 = ~n74924 & n74926;
  assign n74928 = ~n74925 & n74927;
  assign n74929 = P2_P2_INSTQUEUE_REG_3__4_ & n74691;
  assign n74930 = P2_P2_INSTQUEUE_REG_2__4_ & n74693;
  assign n74931 = P2_P2_INSTQUEUE_REG_1__4_ & n74695;
  assign n74932 = P2_P2_INSTQUEUE_REG_0__4_ & n74697;
  assign n74933 = ~n74929 & ~n74930;
  assign n74934 = ~n74931 & n74933;
  assign n74935 = ~n74932 & n74934;
  assign n74936 = P2_P2_INSTQUEUE_REG_15__4_ & n74702;
  assign n74937 = P2_P2_INSTQUEUE_REG_14__4_ & n74704;
  assign n74938 = P2_P2_INSTQUEUE_REG_13__4_ & n74706;
  assign n74939 = P2_P2_INSTQUEUE_REG_12__4_ & n74708;
  assign n74940 = ~n74936 & ~n74937;
  assign n74941 = ~n74938 & n74940;
  assign n74942 = ~n74939 & n74941;
  assign n74943 = P2_P2_INSTQUEUE_REG_11__4_ & n74714;
  assign n74944 = P2_P2_INSTQUEUE_REG_10__4_ & n74716;
  assign n74945 = P2_P2_INSTQUEUE_REG_9__4_ & n74718;
  assign n74946 = P2_P2_INSTQUEUE_REG_8__4_ & n74720;
  assign n74947 = ~n74943 & ~n74944;
  assign n74948 = ~n74945 & n74947;
  assign n74949 = ~n74946 & n74948;
  assign n74950 = n74928 & n74935;
  assign n74951 = n74942 & n74950;
  assign n74952 = n74949 & n74951;
  assign n74953 = n74921 & n74952;
  assign n74954 = ~n74921 & ~n74952;
  assign n74955 = ~n74953 & ~n74954;
  assign n74956 = n73885 & ~n74955;
  assign n74957 = ~n74920 & ~n74956;
  assign n74958 = P2_P2_EAX_REG_25_ & P2_P2_EAX_REG_26_;
  assign n74959 = n74862 & n74958;
  assign n74960 = P2_P2_EAX_REG_27_ & ~n74959;
  assign n74961 = ~P2_P2_EAX_REG_27_ & n74959;
  assign n74962 = ~n74960 & ~n74961;
  assign n74963 = n73891 & ~n74962;
  assign n74964 = ~n74918 & ~n74919;
  assign n74965 = n74957 & n74964;
  assign n14056 = n74963 | ~n74965;
  assign n74967 = ~n68465 & n74336;
  assign n74968 = ~n73582 & n74338;
  assign n74969 = P2_P2_EAX_REG_28_ & ~n73884;
  assign n74970 = n74921 & ~n74952;
  assign n74971 = P2_P2_INSTQUEUE_REG_7__5_ & n74679;
  assign n74972 = P2_P2_INSTQUEUE_REG_6__5_ & n74681;
  assign n74973 = P2_P2_INSTQUEUE_REG_5__5_ & n74683;
  assign n74974 = P2_P2_INSTQUEUE_REG_4__5_ & n74685;
  assign n74975 = ~n74971 & ~n74972;
  assign n74976 = ~n74973 & n74975;
  assign n74977 = ~n74974 & n74976;
  assign n74978 = P2_P2_INSTQUEUE_REG_3__5_ & n74691;
  assign n74979 = P2_P2_INSTQUEUE_REG_2__5_ & n74693;
  assign n74980 = P2_P2_INSTQUEUE_REG_1__5_ & n74695;
  assign n74981 = P2_P2_INSTQUEUE_REG_0__5_ & n74697;
  assign n74982 = ~n74978 & ~n74979;
  assign n74983 = ~n74980 & n74982;
  assign n74984 = ~n74981 & n74983;
  assign n74985 = P2_P2_INSTQUEUE_REG_15__5_ & n74702;
  assign n74986 = P2_P2_INSTQUEUE_REG_14__5_ & n74704;
  assign n74987 = P2_P2_INSTQUEUE_REG_13__5_ & n74706;
  assign n74988 = P2_P2_INSTQUEUE_REG_12__5_ & n74708;
  assign n74989 = ~n74985 & ~n74986;
  assign n74990 = ~n74987 & n74989;
  assign n74991 = ~n74988 & n74990;
  assign n74992 = P2_P2_INSTQUEUE_REG_11__5_ & n74714;
  assign n74993 = P2_P2_INSTQUEUE_REG_10__5_ & n74716;
  assign n74994 = P2_P2_INSTQUEUE_REG_9__5_ & n74718;
  assign n74995 = P2_P2_INSTQUEUE_REG_8__5_ & n74720;
  assign n74996 = ~n74992 & ~n74993;
  assign n74997 = ~n74994 & n74996;
  assign n74998 = ~n74995 & n74997;
  assign n74999 = n74977 & n74984;
  assign n75000 = n74991 & n74999;
  assign n75001 = n74998 & n75000;
  assign n75002 = n74970 & n75001;
  assign n75003 = ~n74970 & ~n75001;
  assign n75004 = ~n75002 & ~n75003;
  assign n75005 = n73885 & ~n75004;
  assign n75006 = P2_P2_EAX_REG_27_ & n74959;
  assign n75007 = ~P2_P2_EAX_REG_28_ & n75006;
  assign n75008 = P2_P2_EAX_REG_28_ & ~n75006;
  assign n75009 = ~n75007 & ~n75008;
  assign n75010 = n73891 & ~n75009;
  assign n75011 = ~n74967 & ~n74968;
  assign n75012 = ~n74969 & n75011;
  assign n75013 = ~n75005 & n75012;
  assign n14061 = n75010 | ~n75013;
  assign n75015 = ~n68443 & n74336;
  assign n75016 = ~n73574 & n74338;
  assign n75017 = P2_P2_EAX_REG_29_ & ~n73884;
  assign n75018 = n74970 & ~n75001;
  assign n75019 = P2_P2_INSTQUEUE_REG_7__6_ & n74679;
  assign n75020 = P2_P2_INSTQUEUE_REG_6__6_ & n74681;
  assign n75021 = P2_P2_INSTQUEUE_REG_5__6_ & n74683;
  assign n75022 = P2_P2_INSTQUEUE_REG_4__6_ & n74685;
  assign n75023 = ~n75019 & ~n75020;
  assign n75024 = ~n75021 & n75023;
  assign n75025 = ~n75022 & n75024;
  assign n75026 = P2_P2_INSTQUEUE_REG_3__6_ & n74691;
  assign n75027 = P2_P2_INSTQUEUE_REG_2__6_ & n74693;
  assign n75028 = P2_P2_INSTQUEUE_REG_1__6_ & n74695;
  assign n75029 = P2_P2_INSTQUEUE_REG_0__6_ & n74697;
  assign n75030 = ~n75026 & ~n75027;
  assign n75031 = ~n75028 & n75030;
  assign n75032 = ~n75029 & n75031;
  assign n75033 = P2_P2_INSTQUEUE_REG_15__6_ & n74702;
  assign n75034 = P2_P2_INSTQUEUE_REG_14__6_ & n74704;
  assign n75035 = P2_P2_INSTQUEUE_REG_13__6_ & n74706;
  assign n75036 = P2_P2_INSTQUEUE_REG_12__6_ & n74708;
  assign n75037 = ~n75033 & ~n75034;
  assign n75038 = ~n75035 & n75037;
  assign n75039 = ~n75036 & n75038;
  assign n75040 = P2_P2_INSTQUEUE_REG_11__6_ & n74714;
  assign n75041 = P2_P2_INSTQUEUE_REG_10__6_ & n74716;
  assign n75042 = P2_P2_INSTQUEUE_REG_9__6_ & n74718;
  assign n75043 = P2_P2_INSTQUEUE_REG_8__6_ & n74720;
  assign n75044 = ~n75040 & ~n75041;
  assign n75045 = ~n75042 & n75044;
  assign n75046 = ~n75043 & n75045;
  assign n75047 = n75025 & n75032;
  assign n75048 = n75039 & n75047;
  assign n75049 = n75046 & n75048;
  assign n75050 = n75018 & n75049;
  assign n75051 = ~n75018 & ~n75049;
  assign n75052 = ~n75050 & ~n75051;
  assign n75053 = n73885 & ~n75052;
  assign n75054 = P2_P2_EAX_REG_27_ & P2_P2_EAX_REG_28_;
  assign n75055 = n74959 & n75054;
  assign n75056 = P2_P2_EAX_REG_29_ & ~n75055;
  assign n75057 = ~P2_P2_EAX_REG_29_ & n75055;
  assign n75058 = ~n75056 & ~n75057;
  assign n75059 = n73891 & ~n75058;
  assign n75060 = ~n75015 & ~n75016;
  assign n75061 = ~n75017 & n75060;
  assign n75062 = ~n75053 & n75061;
  assign n14066 = n75059 | ~n75062;
  assign n75064 = ~n68421 & n74336;
  assign n75065 = ~n73566 & n74338;
  assign n75066 = P2_P2_EAX_REG_30_ & ~n73884;
  assign n75067 = n75018 & ~n75049;
  assign n75068 = P2_P2_INSTQUEUE_REG_7__7_ & n74679;
  assign n75069 = P2_P2_INSTQUEUE_REG_6__7_ & n74681;
  assign n75070 = P2_P2_INSTQUEUE_REG_5__7_ & n74683;
  assign n75071 = P2_P2_INSTQUEUE_REG_4__7_ & n74685;
  assign n75072 = ~n75068 & ~n75069;
  assign n75073 = ~n75070 & n75072;
  assign n75074 = ~n75071 & n75073;
  assign n75075 = P2_P2_INSTQUEUE_REG_3__7_ & n74691;
  assign n75076 = P2_P2_INSTQUEUE_REG_2__7_ & n74693;
  assign n75077 = P2_P2_INSTQUEUE_REG_1__7_ & n74695;
  assign n75078 = P2_P2_INSTQUEUE_REG_0__7_ & n74697;
  assign n75079 = ~n75075 & ~n75076;
  assign n75080 = ~n75077 & n75079;
  assign n75081 = ~n75078 & n75080;
  assign n75082 = P2_P2_INSTQUEUE_REG_15__7_ & n74702;
  assign n75083 = P2_P2_INSTQUEUE_REG_14__7_ & n74704;
  assign n75084 = P2_P2_INSTQUEUE_REG_13__7_ & n74706;
  assign n75085 = P2_P2_INSTQUEUE_REG_12__7_ & n74708;
  assign n75086 = ~n75082 & ~n75083;
  assign n75087 = ~n75084 & n75086;
  assign n75088 = ~n75085 & n75087;
  assign n75089 = P2_P2_INSTQUEUE_REG_11__7_ & n74714;
  assign n75090 = P2_P2_INSTQUEUE_REG_10__7_ & n74716;
  assign n75091 = P2_P2_INSTQUEUE_REG_9__7_ & n74718;
  assign n75092 = P2_P2_INSTQUEUE_REG_8__7_ & n74720;
  assign n75093 = ~n75089 & ~n75090;
  assign n75094 = ~n75091 & n75093;
  assign n75095 = ~n75092 & n75094;
  assign n75096 = n75074 & n75081;
  assign n75097 = n75088 & n75096;
  assign n75098 = n75095 & n75097;
  assign n75099 = n75067 & n75098;
  assign n75100 = ~n75067 & ~n75098;
  assign n75101 = ~n75099 & ~n75100;
  assign n75102 = n73885 & ~n75101;
  assign n75103 = P2_P2_EAX_REG_29_ & n75055;
  assign n75104 = ~P2_P2_EAX_REG_30_ & n75103;
  assign n75105 = P2_P2_EAX_REG_30_ & ~n75103;
  assign n75106 = ~n75104 & ~n75105;
  assign n75107 = n73891 & ~n75106;
  assign n75108 = ~n75064 & ~n75065;
  assign n75109 = ~n75066 & n75108;
  assign n75110 = ~n75102 & n75109;
  assign n14071 = n75107 | ~n75110;
  assign n75112 = P2_P2_EAX_REG_31_ & ~n73884;
  assign n75113 = ~n68396 & n74336;
  assign n75114 = P2_P2_EAX_REG_30_ & n75103;
  assign n75115 = ~P2_P2_EAX_REG_31_ & n75114;
  assign n75116 = P2_P2_EAX_REG_31_ & ~n75114;
  assign n75117 = ~n75115 & ~n75116;
  assign n75118 = n73891 & ~n75117;
  assign n75119 = ~n75112 & ~n75113;
  assign n14076 = n75118 | ~n75119;
  assign n75121 = ~n68055 & ~n68149;
  assign n75122 = n68268 & ~n75121;
  assign n75123 = n67785 & n75122;
  assign n75124 = ~P2_P2_EBX_REG_0_ & n75123;
  assign n75125 = ~n67785 & n75122;
  assign n75126 = P2_P2_INSTQUEUE_REG_0__0_ & n75125;
  assign n75127 = P2_P2_EBX_REG_0_ & ~n75122;
  assign n75128 = ~n75124 & ~n75126;
  assign n14081 = n75127 | ~n75128;
  assign n75130 = ~P2_P2_EBX_REG_0_ & P2_P2_EBX_REG_1_;
  assign n75131 = P2_P2_EBX_REG_0_ & ~P2_P2_EBX_REG_1_;
  assign n75132 = ~n75130 & ~n75131;
  assign n75133 = n75123 & ~n75132;
  assign n75134 = P2_P2_INSTQUEUE_REG_0__1_ & n75125;
  assign n75135 = P2_P2_EBX_REG_1_ & ~n75122;
  assign n75136 = ~n75133 & ~n75134;
  assign n14086 = n75135 | ~n75136;
  assign n75138 = P2_P2_EBX_REG_0_ & P2_P2_EBX_REG_1_;
  assign n75139 = ~P2_P2_EBX_REG_2_ & n75138;
  assign n75140 = P2_P2_EBX_REG_2_ & ~n75138;
  assign n75141 = ~n75139 & ~n75140;
  assign n75142 = n75123 & ~n75141;
  assign n75143 = P2_P2_INSTQUEUE_REG_0__2_ & n75125;
  assign n75144 = P2_P2_EBX_REG_2_ & ~n75122;
  assign n75145 = ~n75142 & ~n75143;
  assign n14091 = n75144 | ~n75145;
  assign n75147 = P2_P2_EBX_REG_0_ & P2_P2_EBX_REG_2_;
  assign n75148 = P2_P2_EBX_REG_1_ & n75147;
  assign n75149 = P2_P2_EBX_REG_3_ & ~n75148;
  assign n75150 = ~P2_P2_EBX_REG_3_ & n75148;
  assign n75151 = ~n75149 & ~n75150;
  assign n75152 = n75123 & ~n75151;
  assign n75153 = P2_P2_INSTQUEUE_REG_0__3_ & n75125;
  assign n75154 = P2_P2_EBX_REG_3_ & ~n75122;
  assign n75155 = ~n75152 & ~n75153;
  assign n14096 = n75154 | ~n75155;
  assign n75157 = P2_P2_EBX_REG_3_ & n75148;
  assign n75158 = ~P2_P2_EBX_REG_4_ & n75157;
  assign n75159 = P2_P2_EBX_REG_4_ & ~n75157;
  assign n75160 = ~n75158 & ~n75159;
  assign n75161 = n75123 & ~n75160;
  assign n75162 = P2_P2_INSTQUEUE_REG_0__4_ & n75125;
  assign n75163 = P2_P2_EBX_REG_4_ & ~n75122;
  assign n75164 = ~n75161 & ~n75162;
  assign n14101 = n75163 | ~n75164;
  assign n75166 = P2_P2_EBX_REG_3_ & P2_P2_EBX_REG_4_;
  assign n75167 = n75148 & n75166;
  assign n75168 = P2_P2_EBX_REG_5_ & ~n75167;
  assign n75169 = ~P2_P2_EBX_REG_5_ & n75167;
  assign n75170 = ~n75168 & ~n75169;
  assign n75171 = n75123 & ~n75170;
  assign n75172 = P2_P2_INSTQUEUE_REG_0__5_ & n75125;
  assign n75173 = P2_P2_EBX_REG_5_ & ~n75122;
  assign n75174 = ~n75171 & ~n75172;
  assign n14106 = n75173 | ~n75174;
  assign n75176 = P2_P2_EBX_REG_5_ & n75167;
  assign n75177 = ~P2_P2_EBX_REG_6_ & n75176;
  assign n75178 = P2_P2_EBX_REG_6_ & ~n75176;
  assign n75179 = ~n75177 & ~n75178;
  assign n75180 = n75123 & ~n75179;
  assign n75181 = P2_P2_INSTQUEUE_REG_0__6_ & n75125;
  assign n75182 = P2_P2_EBX_REG_6_ & ~n75122;
  assign n75183 = ~n75180 & ~n75181;
  assign n14111 = n75182 | ~n75183;
  assign n75185 = P2_P2_EBX_REG_5_ & P2_P2_EBX_REG_6_;
  assign n75186 = n75167 & n75185;
  assign n75187 = P2_P2_EBX_REG_7_ & ~n75186;
  assign n75188 = ~P2_P2_EBX_REG_7_ & n75186;
  assign n75189 = ~n75187 & ~n75188;
  assign n75190 = n75123 & ~n75189;
  assign n75191 = P2_P2_INSTQUEUE_REG_0__7_ & n75125;
  assign n75192 = P2_P2_EBX_REG_7_ & ~n75122;
  assign n75193 = ~n75190 & ~n75191;
  assign n14116 = n75192 | ~n75193;
  assign n75195 = P2_P2_EBX_REG_7_ & n75186;
  assign n75196 = ~P2_P2_EBX_REG_8_ & n75195;
  assign n75197 = P2_P2_EBX_REG_8_ & ~n75195;
  assign n75198 = ~n75196 & ~n75197;
  assign n75199 = n75123 & ~n75198;
  assign n75200 = ~n74026 & n75125;
  assign n75201 = P2_P2_EBX_REG_8_ & ~n75122;
  assign n75202 = ~n75199 & ~n75200;
  assign n14121 = n75201 | ~n75202;
  assign n75204 = P2_P2_EBX_REG_7_ & P2_P2_EBX_REG_8_;
  assign n75205 = n75186 & n75204;
  assign n75206 = P2_P2_EBX_REG_9_ & ~n75205;
  assign n75207 = ~P2_P2_EBX_REG_9_ & n75205;
  assign n75208 = ~n75206 & ~n75207;
  assign n75209 = n75123 & ~n75208;
  assign n75210 = ~n74068 & n75125;
  assign n75211 = P2_P2_EBX_REG_9_ & ~n75122;
  assign n75212 = ~n75209 & ~n75210;
  assign n14126 = n75211 | ~n75212;
  assign n75214 = P2_P2_EBX_REG_10_ & ~n75122;
  assign n75215 = ~n74111 & n75125;
  assign n75216 = P2_P2_EBX_REG_9_ & n75205;
  assign n75217 = ~P2_P2_EBX_REG_10_ & n75216;
  assign n75218 = P2_P2_EBX_REG_10_ & ~n75216;
  assign n75219 = ~n75217 & ~n75218;
  assign n75220 = n75123 & ~n75219;
  assign n75221 = ~n75214 & ~n75215;
  assign n14131 = n75220 | ~n75221;
  assign n75223 = P2_P2_EBX_REG_11_ & ~n75122;
  assign n75224 = ~n74153 & n75125;
  assign n75225 = P2_P2_EBX_REG_9_ & P2_P2_EBX_REG_10_;
  assign n75226 = n75205 & n75225;
  assign n75227 = P2_P2_EBX_REG_11_ & ~n75226;
  assign n75228 = ~P2_P2_EBX_REG_11_ & n75226;
  assign n75229 = ~n75227 & ~n75228;
  assign n75230 = n75123 & ~n75229;
  assign n75231 = ~n75223 & ~n75224;
  assign n14136 = n75230 | ~n75231;
  assign n75233 = P2_P2_EBX_REG_12_ & ~n75122;
  assign n75234 = ~n74196 & n75125;
  assign n75235 = P2_P2_EBX_REG_11_ & n75226;
  assign n75236 = ~P2_P2_EBX_REG_12_ & n75235;
  assign n75237 = P2_P2_EBX_REG_12_ & ~n75235;
  assign n75238 = ~n75236 & ~n75237;
  assign n75239 = n75123 & ~n75238;
  assign n75240 = ~n75233 & ~n75234;
  assign n14141 = n75239 | ~n75240;
  assign n75242 = P2_P2_EBX_REG_13_ & ~n75122;
  assign n75243 = ~n74239 & n75125;
  assign n75244 = P2_P2_EBX_REG_11_ & P2_P2_EBX_REG_12_;
  assign n75245 = n75226 & n75244;
  assign n75246 = P2_P2_EBX_REG_13_ & ~n75245;
  assign n75247 = ~P2_P2_EBX_REG_13_ & n75245;
  assign n75248 = ~n75246 & ~n75247;
  assign n75249 = n75123 & ~n75248;
  assign n75250 = ~n75242 & ~n75243;
  assign n14146 = n75249 | ~n75250;
  assign n75252 = P2_P2_EBX_REG_14_ & ~n75122;
  assign n75253 = ~n74282 & n75125;
  assign n75254 = P2_P2_EBX_REG_13_ & n75245;
  assign n75255 = ~P2_P2_EBX_REG_14_ & n75254;
  assign n75256 = P2_P2_EBX_REG_14_ & ~n75254;
  assign n75257 = ~n75255 & ~n75256;
  assign n75258 = n75123 & ~n75257;
  assign n75259 = ~n75252 & ~n75253;
  assign n14151 = n75258 | ~n75259;
  assign n75261 = P2_P2_EBX_REG_15_ & ~n75122;
  assign n75262 = ~n74324 & n75125;
  assign n75263 = P2_P2_EBX_REG_13_ & P2_P2_EBX_REG_14_;
  assign n75264 = n75245 & n75263;
  assign n75265 = P2_P2_EBX_REG_15_ & ~n75264;
  assign n75266 = ~P2_P2_EBX_REG_15_ & n75264;
  assign n75267 = ~n75265 & ~n75266;
  assign n75268 = n75123 & ~n75267;
  assign n75269 = ~n75261 & ~n75262;
  assign n14156 = n75268 | ~n75269;
  assign n75271 = P2_P2_EBX_REG_16_ & ~n75122;
  assign n75272 = ~n74396 & n75125;
  assign n75273 = P2_P2_EBX_REG_15_ & n75264;
  assign n75274 = ~P2_P2_EBX_REG_16_ & n75273;
  assign n75275 = P2_P2_EBX_REG_16_ & ~n75273;
  assign n75276 = ~n75274 & ~n75275;
  assign n75277 = n75123 & ~n75276;
  assign n75278 = ~n75271 & ~n75272;
  assign n14161 = n75277 | ~n75278;
  assign n75280 = P2_P2_EBX_REG_17_ & ~n75122;
  assign n75281 = ~n74440 & n75125;
  assign n75282 = P2_P2_EBX_REG_15_ & P2_P2_EBX_REG_16_;
  assign n75283 = n75264 & n75282;
  assign n75284 = P2_P2_EBX_REG_17_ & ~n75283;
  assign n75285 = ~P2_P2_EBX_REG_17_ & n75283;
  assign n75286 = ~n75284 & ~n75285;
  assign n75287 = n75123 & ~n75286;
  assign n75288 = ~n75280 & ~n75281;
  assign n14166 = n75287 | ~n75288;
  assign n75290 = P2_P2_EBX_REG_18_ & ~n75122;
  assign n75291 = ~n74485 & n75125;
  assign n75292 = P2_P2_EBX_REG_17_ & n75283;
  assign n75293 = ~P2_P2_EBX_REG_18_ & n75292;
  assign n75294 = P2_P2_EBX_REG_18_ & ~n75292;
  assign n75295 = ~n75293 & ~n75294;
  assign n75296 = n75123 & ~n75295;
  assign n75297 = ~n75290 & ~n75291;
  assign n14171 = n75296 | ~n75297;
  assign n75299 = P2_P2_EBX_REG_19_ & ~n75122;
  assign n75300 = ~n74529 & n75125;
  assign n75301 = P2_P2_EBX_REG_17_ & P2_P2_EBX_REG_18_;
  assign n75302 = n75283 & n75301;
  assign n75303 = P2_P2_EBX_REG_19_ & ~n75302;
  assign n75304 = ~P2_P2_EBX_REG_19_ & n75302;
  assign n75305 = ~n75303 & ~n75304;
  assign n75306 = n75123 & ~n75305;
  assign n75307 = ~n75299 & ~n75300;
  assign n14176 = n75306 | ~n75307;
  assign n75309 = P2_P2_EBX_REG_20_ & ~n75122;
  assign n75310 = ~n74574 & n75125;
  assign n75311 = P2_P2_EBX_REG_19_ & n75302;
  assign n75312 = ~P2_P2_EBX_REG_20_ & n75311;
  assign n75313 = P2_P2_EBX_REG_20_ & ~n75311;
  assign n75314 = ~n75312 & ~n75313;
  assign n75315 = n75123 & ~n75314;
  assign n75316 = ~n75309 & ~n75310;
  assign n14181 = n75315 | ~n75316;
  assign n75318 = P2_P2_EBX_REG_21_ & ~n75122;
  assign n75319 = ~n74618 & n75125;
  assign n75320 = P2_P2_EBX_REG_19_ & P2_P2_EBX_REG_20_;
  assign n75321 = n75302 & n75320;
  assign n75322 = P2_P2_EBX_REG_21_ & ~n75321;
  assign n75323 = ~P2_P2_EBX_REG_21_ & n75321;
  assign n75324 = ~n75322 & ~n75323;
  assign n75325 = n75123 & ~n75324;
  assign n75326 = ~n75318 & ~n75319;
  assign n14186 = n75325 | ~n75326;
  assign n75328 = P2_P2_EBX_REG_22_ & ~n75122;
  assign n75329 = ~n74663 & n75125;
  assign n75330 = P2_P2_EBX_REG_21_ & n75321;
  assign n75331 = ~P2_P2_EBX_REG_22_ & n75330;
  assign n75332 = P2_P2_EBX_REG_22_ & ~n75330;
  assign n75333 = ~n75331 & ~n75332;
  assign n75334 = n75123 & ~n75333;
  assign n75335 = ~n75328 & ~n75329;
  assign n14191 = n75334 | ~n75335;
  assign n75337 = P2_P2_EBX_REG_23_ & ~n75122;
  assign n75338 = ~n74761 & n75125;
  assign n75339 = P2_P2_EBX_REG_21_ & P2_P2_EBX_REG_22_;
  assign n75340 = n75321 & n75339;
  assign n75341 = P2_P2_EBX_REG_23_ & ~n75340;
  assign n75342 = ~P2_P2_EBX_REG_23_ & n75340;
  assign n75343 = ~n75341 & ~n75342;
  assign n75344 = n75123 & ~n75343;
  assign n75345 = ~n75337 & ~n75338;
  assign n14196 = n75344 | ~n75345;
  assign n75347 = P2_P2_EBX_REG_24_ & ~n75122;
  assign n75348 = ~n74810 & n75125;
  assign n75349 = P2_P2_EBX_REG_23_ & n75340;
  assign n75350 = ~P2_P2_EBX_REG_24_ & n75349;
  assign n75351 = P2_P2_EBX_REG_24_ & ~n75349;
  assign n75352 = ~n75350 & ~n75351;
  assign n75353 = n75123 & ~n75352;
  assign n75354 = ~n75347 & ~n75348;
  assign n14201 = n75353 | ~n75354;
  assign n75356 = P2_P2_EBX_REG_25_ & ~n75122;
  assign n75357 = ~n74858 & n75125;
  assign n75358 = P2_P2_EBX_REG_23_ & P2_P2_EBX_REG_24_;
  assign n75359 = n75340 & n75358;
  assign n75360 = P2_P2_EBX_REG_25_ & ~n75359;
  assign n75361 = ~P2_P2_EBX_REG_25_ & n75359;
  assign n75362 = ~n75360 & ~n75361;
  assign n75363 = n75123 & ~n75362;
  assign n75364 = ~n75356 & ~n75357;
  assign n14206 = n75363 | ~n75364;
  assign n75366 = P2_P2_EBX_REG_26_ & ~n75122;
  assign n75367 = ~n74907 & n75125;
  assign n75368 = P2_P2_EBX_REG_25_ & n75359;
  assign n75369 = ~P2_P2_EBX_REG_26_ & n75368;
  assign n75370 = P2_P2_EBX_REG_26_ & ~n75368;
  assign n75371 = ~n75369 & ~n75370;
  assign n75372 = n75123 & ~n75371;
  assign n75373 = ~n75366 & ~n75367;
  assign n14211 = n75372 | ~n75373;
  assign n75375 = P2_P2_EBX_REG_27_ & ~n75122;
  assign n75376 = ~n74955 & n75125;
  assign n75377 = P2_P2_EBX_REG_25_ & P2_P2_EBX_REG_26_;
  assign n75378 = n75359 & n75377;
  assign n75379 = P2_P2_EBX_REG_27_ & ~n75378;
  assign n75380 = ~P2_P2_EBX_REG_27_ & n75378;
  assign n75381 = ~n75379 & ~n75380;
  assign n75382 = n75123 & ~n75381;
  assign n75383 = ~n75375 & ~n75376;
  assign n14216 = n75382 | ~n75383;
  assign n75385 = P2_P2_EBX_REG_28_ & ~n75122;
  assign n75386 = ~n75004 & n75125;
  assign n75387 = P2_P2_EBX_REG_27_ & n75378;
  assign n75388 = ~P2_P2_EBX_REG_28_ & n75387;
  assign n75389 = P2_P2_EBX_REG_28_ & ~n75387;
  assign n75390 = ~n75388 & ~n75389;
  assign n75391 = n75123 & ~n75390;
  assign n75392 = ~n75385 & ~n75386;
  assign n14221 = n75391 | ~n75392;
  assign n75394 = P2_P2_EBX_REG_29_ & ~n75122;
  assign n75395 = ~n75052 & n75125;
  assign n75396 = P2_P2_EBX_REG_27_ & P2_P2_EBX_REG_28_;
  assign n75397 = n75378 & n75396;
  assign n75398 = P2_P2_EBX_REG_29_ & ~n75397;
  assign n75399 = ~P2_P2_EBX_REG_29_ & n75397;
  assign n75400 = ~n75398 & ~n75399;
  assign n75401 = n75123 & ~n75400;
  assign n75402 = ~n75394 & ~n75395;
  assign n14226 = n75401 | ~n75402;
  assign n75404 = P2_P2_EBX_REG_30_ & ~n75122;
  assign n75405 = ~n75101 & n75125;
  assign n75406 = P2_P2_EBX_REG_29_ & n75397;
  assign n75407 = ~P2_P2_EBX_REG_30_ & n75406;
  assign n75408 = P2_P2_EBX_REG_30_ & ~n75406;
  assign n75409 = ~n75407 & ~n75408;
  assign n75410 = n75123 & ~n75409;
  assign n75411 = ~n75404 & ~n75405;
  assign n14231 = n75410 | ~n75411;
  assign n75413 = P2_P2_EBX_REG_31_ & ~n75122;
  assign n75414 = P2_P2_EBX_REG_30_ & n75406;
  assign n75415 = ~P2_P2_EBX_REG_31_ & n75414;
  assign n75416 = P2_P2_EBX_REG_31_ & ~n75414;
  assign n75417 = ~n75415 & ~n75416;
  assign n75418 = n75123 & ~n75417;
  assign n14236 = n75413 | n75418;
  assign n75420 = ~n68279 & ~n68318;
  assign n75421 = ~n69954 & n75420;
  assign n75422 = n68146 & n68154;
  assign n75423 = n68268 & ~n75422;
  assign n75424 = n75421 & ~n75423;
  assign n75425 = P2_P2_STATE2_REG_2_ & ~n75424;
  assign n75426 = n67996 & n75425;
  assign n75427 = ~n67629 & n75426;
  assign n75428 = ~P2_P2_EBX_REG_31_ & n75427;
  assign n75429 = n67914 & n75425;
  assign n75430 = ~n67632 & n75429;
  assign n75431 = n67632 & n75429;
  assign n75432 = ~n67629 & n75431;
  assign n75433 = ~n75428 & ~n75430;
  assign n75434 = ~n75432 & n75433;
  assign n75435 = P2_P2_EBX_REG_0_ & ~n75434;
  assign n75436 = n67629 & n75431;
  assign n75437 = P2_P2_REIP_REG_0_ & n75436;
  assign n75438 = P2_P2_EBX_REG_31_ & n75427;
  assign n75439 = P2_P2_EBX_REG_0_ & n75438;
  assign n75440 = n67991 & n75425;
  assign n75441 = ~P2_P2_INSTQUEUERD_ADDR_REG_0_ & n75440;
  assign n75442 = n67987 & n75425;
  assign n75443 = ~P2_P2_INSTQUEUERD_ADDR_REG_0_ & n75442;
  assign n75444 = ~n75441 & ~n75443;
  assign n75445 = ~n75437 & ~n75439;
  assign n75446 = n75444 & n75445;
  assign n75447 = n67629 & n75426;
  assign n75448 = P2_P2_REIP_REG_0_ & n75447;
  assign n75449 = P2_P2_STATE2_REG_1_ & ~n75424;
  assign n75450 = n73537 & n75449;
  assign n75451 = P2_P2_PHYADDRPOINTER_REG_0_ & n75450;
  assign n75452 = P2_P2_REIP_REG_0_ & n75424;
  assign n75453 = P2_P2_STATE2_REG_3_ & ~n75424;
  assign n75454 = P2_P2_PHYADDRPOINTER_REG_0_ & n75453;
  assign n75455 = ~n75452 & ~n75454;
  assign n75456 = ~n73537 & n75449;
  assign n75457 = P2_P2_PHYADDRPOINTER_REG_0_ & n75456;
  assign n75458 = n75455 & ~n75457;
  assign n75459 = ~n75435 & n75446;
  assign n75460 = ~n75448 & n75459;
  assign n75461 = ~n75451 & n75460;
  assign n14241 = ~n75458 | ~n75461;
  assign n75463 = P2_P2_EBX_REG_1_ & ~n75434;
  assign n75464 = ~P2_P2_REIP_REG_1_ & n75436;
  assign n75465 = ~n75132 & n75438;
  assign n75466 = ~n67638 & ~n67643;
  assign n75467 = n75440 & ~n75466;
  assign n75468 = n75442 & ~n75466;
  assign n75469 = ~n75467 & ~n75468;
  assign n75470 = ~n75464 & ~n75465;
  assign n75471 = n75469 & n75470;
  assign n75472 = ~P2_P2_REIP_REG_1_ & n75447;
  assign n75473 = ~P2_P2_PHYADDRPOINTER_REG_1_ & n75450;
  assign n75474 = P2_P2_REIP_REG_1_ & n75424;
  assign n75475 = P2_P2_PHYADDRPOINTER_REG_1_ & n75453;
  assign n75476 = ~n75474 & ~n75475;
  assign n75477 = P2_P2_PHYADDRPOINTER_REG_0_ & P2_P2_PHYADDRPOINTER_REG_1_;
  assign n75478 = ~P2_P2_PHYADDRPOINTER_REG_0_ & ~P2_P2_PHYADDRPOINTER_REG_1_;
  assign n75479 = ~n75477 & ~n75478;
  assign n75480 = n75456 & ~n75479;
  assign n75481 = n75476 & ~n75480;
  assign n75482 = ~n75463 & n75471;
  assign n75483 = ~n75472 & n75482;
  assign n75484 = ~n75473 & n75483;
  assign n14246 = ~n75481 | ~n75484;
  assign n75486 = P2_P2_EBX_REG_2_ & ~n75434;
  assign n75487 = P2_P2_REIP_REG_1_ & ~P2_P2_REIP_REG_2_;
  assign n75488 = ~P2_P2_REIP_REG_1_ & P2_P2_REIP_REG_2_;
  assign n75489 = ~n75487 & ~n75488;
  assign n75490 = n75436 & ~n75489;
  assign n75491 = ~P2_P2_EBX_REG_0_ & ~P2_P2_EBX_REG_1_;
  assign n75492 = P2_P2_EBX_REG_2_ & ~n75491;
  assign n75493 = ~P2_P2_EBX_REG_2_ & n75491;
  assign n75494 = ~n75492 & ~n75493;
  assign n75495 = n75438 & n75494;
  assign n75496 = ~n68116 & n75440;
  assign n75497 = ~n68116 & n75442;
  assign n75498 = ~n75496 & ~n75497;
  assign n75499 = ~n75490 & ~n75495;
  assign n75500 = n75498 & n75499;
  assign n75501 = n75447 & ~n75489;
  assign n75502 = ~n72871 & n75450;
  assign n75503 = P2_P2_REIP_REG_2_ & n75424;
  assign n75504 = P2_P2_PHYADDRPOINTER_REG_2_ & n75453;
  assign n75505 = ~n75503 & ~n75504;
  assign n75506 = ~P2_P2_PHYADDRPOINTER_REG_0_ & P2_P2_PHYADDRPOINTER_REG_1_;
  assign n75507 = ~n72871 & ~n75506;
  assign n75508 = n72871 & n75506;
  assign n75509 = ~n75507 & ~n75508;
  assign n75510 = n75456 & n75509;
  assign n75511 = n75505 & ~n75510;
  assign n75512 = ~n75486 & n75500;
  assign n75513 = ~n75501 & n75512;
  assign n75514 = ~n75502 & n75513;
  assign n14251 = ~n75511 | ~n75514;
  assign n75516 = P2_P2_EBX_REG_3_ & ~n75434;
  assign n75517 = P2_P2_REIP_REG_1_ & P2_P2_REIP_REG_2_;
  assign n75518 = ~P2_P2_REIP_REG_3_ & n75517;
  assign n75519 = P2_P2_REIP_REG_3_ & ~n75517;
  assign n75520 = ~n75518 & ~n75519;
  assign n75521 = n75436 & ~n75520;
  assign n75522 = ~P2_P2_EBX_REG_3_ & n75493;
  assign n75523 = P2_P2_EBX_REG_3_ & ~n75493;
  assign n75524 = ~n75522 & ~n75523;
  assign n75525 = n75438 & n75524;
  assign n75526 = ~P2_P2_INSTQUEUERD_ADDR_REG_3_ & n68164;
  assign n75527 = ~n68165 & ~n75526;
  assign n75528 = n75440 & ~n75527;
  assign n75529 = n75442 & ~n75527;
  assign n75530 = ~n75528 & ~n75529;
  assign n75531 = ~n75521 & ~n75525;
  assign n75532 = n75530 & n75531;
  assign n75533 = n75447 & ~n75520;
  assign n75534 = ~n72893 & n75450;
  assign n75535 = P2_P2_REIP_REG_3_ & n75424;
  assign n75536 = P2_P2_PHYADDRPOINTER_REG_3_ & n75453;
  assign n75537 = ~n75535 & ~n75536;
  assign n75538 = n72893 & n75508;
  assign n75539 = ~n72893 & ~n75508;
  assign n75540 = ~n75538 & ~n75539;
  assign n75541 = n75456 & n75540;
  assign n75542 = n75537 & ~n75541;
  assign n75543 = ~n75516 & n75532;
  assign n75544 = ~n75533 & n75543;
  assign n75545 = ~n75534 & n75544;
  assign n14256 = ~n75542 | ~n75545;
  assign n75547 = P2_P2_INSTQUEUERD_ADDR_REG_3_ & n68164;
  assign n75548 = ~P2_P2_INSTQUEUERD_ADDR_REG_4_ & n75547;
  assign n75549 = P2_P2_INSTQUEUERD_ADDR_REG_4_ & ~n75547;
  assign n75550 = ~n75548 & ~n75549;
  assign n75551 = n75442 & ~n75550;
  assign n75552 = n75440 & ~n75550;
  assign n75553 = ~n75551 & ~n75552;
  assign n75554 = P2_P2_EBX_REG_4_ & ~n75434;
  assign n75555 = P2_P2_EBX_REG_4_ & ~n75522;
  assign n75556 = ~P2_P2_EBX_REG_3_ & ~P2_P2_EBX_REG_4_;
  assign n75557 = n75493 & n75556;
  assign n75558 = ~n75555 & ~n75557;
  assign n75559 = n75438 & n75558;
  assign n75560 = n69953 & ~n75424;
  assign n75561 = P2_P2_REIP_REG_3_ & n75517;
  assign n75562 = ~P2_P2_REIP_REG_4_ & n75561;
  assign n75563 = P2_P2_REIP_REG_4_ & ~n75561;
  assign n75564 = ~n75562 & ~n75563;
  assign n75565 = n75436 & ~n75564;
  assign n75566 = ~n75559 & ~n75560;
  assign n75567 = ~n75565 & n75566;
  assign n75568 = n75447 & ~n75564;
  assign n75569 = ~n72914 & n75450;
  assign n75570 = n75553 & ~n75554;
  assign n75571 = n75567 & n75570;
  assign n75572 = ~n75568 & n75571;
  assign n75573 = ~n75569 & n75572;
  assign n75574 = P2_P2_REIP_REG_4_ & n75424;
  assign n75575 = P2_P2_PHYADDRPOINTER_REG_4_ & n75453;
  assign n75576 = ~n75574 & ~n75575;
  assign n75577 = ~n72914 & ~n75538;
  assign n75578 = n72893 & n72914;
  assign n75579 = n75508 & n75578;
  assign n75580 = ~n75577 & ~n75579;
  assign n75581 = n75456 & n75580;
  assign n75582 = n75576 & ~n75581;
  assign n14261 = ~n75573 | ~n75582;
  assign n75584 = P2_P2_INSTQUEUERD_ADDR_REG_4_ & n75547;
  assign n75585 = n75442 & n75584;
  assign n75586 = n75440 & n75584;
  assign n75587 = ~n75585 & ~n75586;
  assign n75588 = P2_P2_EBX_REG_5_ & ~n75434;
  assign n75589 = ~P2_P2_EBX_REG_5_ & n75557;
  assign n75590 = P2_P2_EBX_REG_5_ & ~n75557;
  assign n75591 = ~n75589 & ~n75590;
  assign n75592 = n75438 & n75591;
  assign n75593 = P2_P2_REIP_REG_4_ & n75561;
  assign n75594 = ~P2_P2_REIP_REG_5_ & n75593;
  assign n75595 = P2_P2_REIP_REG_5_ & ~n75593;
  assign n75596 = ~n75594 & ~n75595;
  assign n75597 = n75436 & ~n75596;
  assign n75598 = ~n75560 & ~n75592;
  assign n75599 = ~n75597 & n75598;
  assign n75600 = n75447 & ~n75596;
  assign n75601 = ~n72937 & n75450;
  assign n75602 = n75587 & ~n75588;
  assign n75603 = n75599 & n75602;
  assign n75604 = ~n75600 & n75603;
  assign n75605 = ~n75601 & n75604;
  assign n75606 = P2_P2_REIP_REG_5_ & n75424;
  assign n75607 = P2_P2_PHYADDRPOINTER_REG_5_ & n75453;
  assign n75608 = ~n75606 & ~n75607;
  assign n75609 = n72937 & n75579;
  assign n75610 = ~n72937 & ~n75579;
  assign n75611 = ~n75609 & ~n75610;
  assign n75612 = n75456 & n75611;
  assign n75613 = n75608 & ~n75612;
  assign n14266 = ~n75605 | ~n75613;
  assign n75615 = P2_P2_REIP_REG_5_ & n75593;
  assign n75616 = ~P2_P2_REIP_REG_6_ & n75615;
  assign n75617 = P2_P2_REIP_REG_6_ & ~n75615;
  assign n75618 = ~n75616 & ~n75617;
  assign n75619 = n75447 & ~n75618;
  assign n75620 = P2_P2_EBX_REG_6_ & ~n75434;
  assign n75621 = P2_P2_EBX_REG_6_ & ~n75589;
  assign n75622 = ~P2_P2_EBX_REG_5_ & ~P2_P2_EBX_REG_6_;
  assign n75623 = n75557 & n75622;
  assign n75624 = ~n75621 & ~n75623;
  assign n75625 = n75438 & n75624;
  assign n75626 = n75436 & ~n75618;
  assign n75627 = ~n75560 & ~n75625;
  assign n75628 = ~n75626 & n75627;
  assign n75629 = ~n72960 & ~n75609;
  assign n75630 = n72937 & n72960;
  assign n75631 = n75579 & n75630;
  assign n75632 = ~n75629 & ~n75631;
  assign n75633 = n75456 & n75632;
  assign n75634 = P2_P2_REIP_REG_6_ & n75424;
  assign n75635 = P2_P2_PHYADDRPOINTER_REG_6_ & n75453;
  assign n75636 = ~n75634 & ~n75635;
  assign n75637 = ~n72960 & n75450;
  assign n75638 = n75636 & ~n75637;
  assign n75639 = ~n75619 & ~n75620;
  assign n75640 = n75628 & n75639;
  assign n75641 = ~n75633 & n75640;
  assign n14271 = ~n75638 | ~n75641;
  assign n75643 = P2_P2_REIP_REG_6_ & n75615;
  assign n75644 = ~P2_P2_REIP_REG_7_ & n75643;
  assign n75645 = P2_P2_REIP_REG_7_ & ~n75643;
  assign n75646 = ~n75644 & ~n75645;
  assign n75647 = n75447 & ~n75646;
  assign n75648 = P2_P2_EBX_REG_7_ & ~n75434;
  assign n75649 = ~P2_P2_EBX_REG_7_ & n75623;
  assign n75650 = P2_P2_EBX_REG_7_ & ~n75623;
  assign n75651 = ~n75649 & ~n75650;
  assign n75652 = n75438 & n75651;
  assign n75653 = n75436 & ~n75646;
  assign n75654 = ~n75560 & ~n75652;
  assign n75655 = ~n75653 & n75654;
  assign n75656 = n72983 & n75631;
  assign n75657 = ~n72983 & ~n75631;
  assign n75658 = ~n75656 & ~n75657;
  assign n75659 = n75456 & n75658;
  assign n75660 = P2_P2_REIP_REG_7_ & n75424;
  assign n75661 = P2_P2_PHYADDRPOINTER_REG_7_ & n75453;
  assign n75662 = ~n75660 & ~n75661;
  assign n75663 = ~n72983 & n75450;
  assign n75664 = n75662 & ~n75663;
  assign n75665 = ~n75647 & ~n75648;
  assign n75666 = n75655 & n75665;
  assign n75667 = ~n75659 & n75666;
  assign n14276 = ~n75664 | ~n75667;
  assign n75669 = P2_P2_REIP_REG_7_ & n75643;
  assign n75670 = ~P2_P2_REIP_REG_8_ & n75669;
  assign n75671 = P2_P2_REIP_REG_8_ & ~n75669;
  assign n75672 = ~n75670 & ~n75671;
  assign n75673 = n75447 & ~n75672;
  assign n75674 = P2_P2_EBX_REG_8_ & ~n75434;
  assign n75675 = P2_P2_EBX_REG_8_ & ~n75649;
  assign n75676 = ~P2_P2_EBX_REG_7_ & ~P2_P2_EBX_REG_8_;
  assign n75677 = n75623 & n75676;
  assign n75678 = ~n75675 & ~n75677;
  assign n75679 = n75438 & n75678;
  assign n75680 = n75436 & ~n75672;
  assign n75681 = ~n75560 & ~n75679;
  assign n75682 = ~n75680 & n75681;
  assign n75683 = ~n73006 & ~n75656;
  assign n75684 = n72983 & n73006;
  assign n75685 = n75631 & n75684;
  assign n75686 = ~n75683 & ~n75685;
  assign n75687 = n75456 & n75686;
  assign n75688 = P2_P2_REIP_REG_8_ & n75424;
  assign n75689 = P2_P2_PHYADDRPOINTER_REG_8_ & n75453;
  assign n75690 = ~n75688 & ~n75689;
  assign n75691 = ~n73006 & n75450;
  assign n75692 = n75690 & ~n75691;
  assign n75693 = ~n75673 & ~n75674;
  assign n75694 = n75682 & n75693;
  assign n75695 = ~n75687 & n75694;
  assign n14281 = ~n75692 | ~n75695;
  assign n75697 = P2_P2_REIP_REG_8_ & n75669;
  assign n75698 = ~P2_P2_REIP_REG_9_ & n75697;
  assign n75699 = P2_P2_REIP_REG_9_ & ~n75697;
  assign n75700 = ~n75698 & ~n75699;
  assign n75701 = n75447 & ~n75700;
  assign n75702 = P2_P2_EBX_REG_9_ & ~n75434;
  assign n75703 = ~P2_P2_EBX_REG_9_ & n75677;
  assign n75704 = P2_P2_EBX_REG_9_ & ~n75677;
  assign n75705 = ~n75703 & ~n75704;
  assign n75706 = n75438 & n75705;
  assign n75707 = n75436 & ~n75700;
  assign n75708 = ~n75560 & ~n75706;
  assign n75709 = ~n75707 & n75708;
  assign n75710 = n73029 & n75685;
  assign n75711 = ~n73029 & ~n75685;
  assign n75712 = ~n75710 & ~n75711;
  assign n75713 = n75456 & n75712;
  assign n75714 = P2_P2_REIP_REG_9_ & n75424;
  assign n75715 = P2_P2_PHYADDRPOINTER_REG_9_ & n75453;
  assign n75716 = ~n75714 & ~n75715;
  assign n75717 = ~n73029 & n75450;
  assign n75718 = n75716 & ~n75717;
  assign n75719 = ~n75701 & ~n75702;
  assign n75720 = n75709 & n75719;
  assign n75721 = ~n75713 & n75720;
  assign n14286 = ~n75718 | ~n75721;
  assign n75723 = P2_P2_REIP_REG_9_ & n75697;
  assign n75724 = ~P2_P2_REIP_REG_10_ & n75723;
  assign n75725 = P2_P2_REIP_REG_10_ & ~n75723;
  assign n75726 = ~n75724 & ~n75725;
  assign n75727 = n75447 & ~n75726;
  assign n75728 = P2_P2_EBX_REG_10_ & ~n75434;
  assign n75729 = P2_P2_EBX_REG_10_ & ~n75703;
  assign n75730 = ~P2_P2_EBX_REG_9_ & ~P2_P2_EBX_REG_10_;
  assign n75731 = n75677 & n75730;
  assign n75732 = ~n75729 & ~n75731;
  assign n75733 = n75438 & n75732;
  assign n75734 = n75436 & ~n75726;
  assign n75735 = ~n75560 & ~n75733;
  assign n75736 = ~n75734 & n75735;
  assign n75737 = ~n73052 & ~n75710;
  assign n75738 = n73029 & n73052;
  assign n75739 = n75685 & n75738;
  assign n75740 = ~n75737 & ~n75739;
  assign n75741 = n75456 & n75740;
  assign n75742 = P2_P2_REIP_REG_10_ & n75424;
  assign n75743 = P2_P2_PHYADDRPOINTER_REG_10_ & n75453;
  assign n75744 = ~n75742 & ~n75743;
  assign n75745 = ~n73052 & n75450;
  assign n75746 = n75744 & ~n75745;
  assign n75747 = ~n75727 & ~n75728;
  assign n75748 = n75736 & n75747;
  assign n75749 = ~n75741 & n75748;
  assign n14291 = ~n75746 | ~n75749;
  assign n75751 = P2_P2_REIP_REG_10_ & n75723;
  assign n75752 = ~P2_P2_REIP_REG_11_ & n75751;
  assign n75753 = P2_P2_REIP_REG_11_ & ~n75751;
  assign n75754 = ~n75752 & ~n75753;
  assign n75755 = n75447 & ~n75754;
  assign n75756 = P2_P2_EBX_REG_11_ & ~n75434;
  assign n75757 = ~P2_P2_EBX_REG_11_ & n75731;
  assign n75758 = P2_P2_EBX_REG_11_ & ~n75731;
  assign n75759 = ~n75757 & ~n75758;
  assign n75760 = n75438 & n75759;
  assign n75761 = n75436 & ~n75754;
  assign n75762 = ~n75560 & ~n75760;
  assign n75763 = ~n75761 & n75762;
  assign n75764 = n73075 & n75739;
  assign n75765 = ~n73075 & ~n75739;
  assign n75766 = ~n75764 & ~n75765;
  assign n75767 = n75456 & n75766;
  assign n75768 = P2_P2_REIP_REG_11_ & n75424;
  assign n75769 = P2_P2_PHYADDRPOINTER_REG_11_ & n75453;
  assign n75770 = ~n75768 & ~n75769;
  assign n75771 = ~n73075 & n75450;
  assign n75772 = n75770 & ~n75771;
  assign n75773 = ~n75755 & ~n75756;
  assign n75774 = n75763 & n75773;
  assign n75775 = ~n75767 & n75774;
  assign n14296 = ~n75772 | ~n75775;
  assign n75777 = P2_P2_REIP_REG_11_ & n75751;
  assign n75778 = ~P2_P2_REIP_REG_12_ & n75777;
  assign n75779 = P2_P2_REIP_REG_12_ & ~n75777;
  assign n75780 = ~n75778 & ~n75779;
  assign n75781 = n75447 & ~n75780;
  assign n75782 = P2_P2_EBX_REG_12_ & ~n75434;
  assign n75783 = P2_P2_EBX_REG_12_ & ~n75757;
  assign n75784 = ~P2_P2_EBX_REG_11_ & ~P2_P2_EBX_REG_12_;
  assign n75785 = n75731 & n75784;
  assign n75786 = ~n75783 & ~n75785;
  assign n75787 = n75438 & n75786;
  assign n75788 = n75436 & ~n75780;
  assign n75789 = ~n75560 & ~n75787;
  assign n75790 = ~n75788 & n75789;
  assign n75791 = ~n73098 & ~n75764;
  assign n75792 = n73075 & n73098;
  assign n75793 = n75739 & n75792;
  assign n75794 = ~n75791 & ~n75793;
  assign n75795 = n75456 & n75794;
  assign n75796 = P2_P2_REIP_REG_12_ & n75424;
  assign n75797 = P2_P2_PHYADDRPOINTER_REG_12_ & n75453;
  assign n75798 = ~n75796 & ~n75797;
  assign n75799 = ~n73098 & n75450;
  assign n75800 = n75798 & ~n75799;
  assign n75801 = ~n75781 & ~n75782;
  assign n75802 = n75790 & n75801;
  assign n75803 = ~n75795 & n75802;
  assign n14301 = ~n75800 | ~n75803;
  assign n75805 = P2_P2_REIP_REG_12_ & n75777;
  assign n75806 = ~P2_P2_REIP_REG_13_ & n75805;
  assign n75807 = P2_P2_REIP_REG_13_ & ~n75805;
  assign n75808 = ~n75806 & ~n75807;
  assign n75809 = n75447 & ~n75808;
  assign n75810 = P2_P2_EBX_REG_13_ & ~n75434;
  assign n75811 = ~P2_P2_EBX_REG_13_ & n75785;
  assign n75812 = P2_P2_EBX_REG_13_ & ~n75785;
  assign n75813 = ~n75811 & ~n75812;
  assign n75814 = n75438 & n75813;
  assign n75815 = n75436 & ~n75808;
  assign n75816 = ~n75560 & ~n75814;
  assign n75817 = ~n75815 & n75816;
  assign n75818 = n73121 & n75793;
  assign n75819 = ~n73121 & ~n75793;
  assign n75820 = ~n75818 & ~n75819;
  assign n75821 = n75456 & n75820;
  assign n75822 = P2_P2_REIP_REG_13_ & n75424;
  assign n75823 = P2_P2_PHYADDRPOINTER_REG_13_ & n75453;
  assign n75824 = ~n75822 & ~n75823;
  assign n75825 = ~n73121 & n75450;
  assign n75826 = n75824 & ~n75825;
  assign n75827 = ~n75809 & ~n75810;
  assign n75828 = n75817 & n75827;
  assign n75829 = ~n75821 & n75828;
  assign n14306 = ~n75826 | ~n75829;
  assign n75831 = P2_P2_REIP_REG_13_ & n75805;
  assign n75832 = ~P2_P2_REIP_REG_14_ & n75831;
  assign n75833 = P2_P2_REIP_REG_14_ & ~n75831;
  assign n75834 = ~n75832 & ~n75833;
  assign n75835 = n75447 & ~n75834;
  assign n75836 = P2_P2_EBX_REG_14_ & ~n75434;
  assign n75837 = P2_P2_EBX_REG_14_ & ~n75811;
  assign n75838 = ~P2_P2_EBX_REG_13_ & ~P2_P2_EBX_REG_14_;
  assign n75839 = n75785 & n75838;
  assign n75840 = ~n75837 & ~n75839;
  assign n75841 = n75438 & n75840;
  assign n75842 = n75436 & ~n75834;
  assign n75843 = ~n75560 & ~n75841;
  assign n75844 = ~n75842 & n75843;
  assign n75845 = ~n73144 & ~n75818;
  assign n75846 = n73121 & n73144;
  assign n75847 = n75793 & n75846;
  assign n75848 = ~n75845 & ~n75847;
  assign n75849 = n75456 & n75848;
  assign n75850 = P2_P2_REIP_REG_14_ & n75424;
  assign n75851 = P2_P2_PHYADDRPOINTER_REG_14_ & n75453;
  assign n75852 = ~n75850 & ~n75851;
  assign n75853 = ~n73144 & n75450;
  assign n75854 = n75852 & ~n75853;
  assign n75855 = ~n75835 & ~n75836;
  assign n75856 = n75844 & n75855;
  assign n75857 = ~n75849 & n75856;
  assign n14311 = ~n75854 | ~n75857;
  assign n75859 = P2_P2_REIP_REG_14_ & n75831;
  assign n75860 = ~P2_P2_REIP_REG_15_ & n75859;
  assign n75861 = P2_P2_REIP_REG_15_ & ~n75859;
  assign n75862 = ~n75860 & ~n75861;
  assign n75863 = n75447 & ~n75862;
  assign n75864 = P2_P2_EBX_REG_15_ & ~n75434;
  assign n75865 = ~P2_P2_EBX_REG_15_ & n75839;
  assign n75866 = P2_P2_EBX_REG_15_ & ~n75839;
  assign n75867 = ~n75865 & ~n75866;
  assign n75868 = n75438 & n75867;
  assign n75869 = n75436 & ~n75862;
  assign n75870 = ~n75560 & ~n75868;
  assign n75871 = ~n75869 & n75870;
  assign n75872 = n73167 & n75847;
  assign n75873 = ~n73167 & ~n75847;
  assign n75874 = ~n75872 & ~n75873;
  assign n75875 = n75456 & n75874;
  assign n75876 = P2_P2_REIP_REG_15_ & n75424;
  assign n75877 = P2_P2_PHYADDRPOINTER_REG_15_ & n75453;
  assign n75878 = ~n75876 & ~n75877;
  assign n75879 = ~n73167 & n75450;
  assign n75880 = n75878 & ~n75879;
  assign n75881 = ~n75863 & ~n75864;
  assign n75882 = n75871 & n75881;
  assign n75883 = ~n75875 & n75882;
  assign n14316 = ~n75880 | ~n75883;
  assign n75885 = P2_P2_REIP_REG_15_ & n75859;
  assign n75886 = ~P2_P2_REIP_REG_16_ & n75885;
  assign n75887 = P2_P2_REIP_REG_16_ & ~n75885;
  assign n75888 = ~n75886 & ~n75887;
  assign n75889 = n75447 & ~n75888;
  assign n75890 = P2_P2_EBX_REG_16_ & ~n75434;
  assign n75891 = P2_P2_EBX_REG_16_ & ~n75865;
  assign n75892 = ~P2_P2_EBX_REG_15_ & ~P2_P2_EBX_REG_16_;
  assign n75893 = n75839 & n75892;
  assign n75894 = ~n75891 & ~n75893;
  assign n75895 = n75438 & n75894;
  assign n75896 = n75436 & ~n75888;
  assign n75897 = ~n75560 & ~n75895;
  assign n75898 = ~n75896 & n75897;
  assign n75899 = ~n73190 & ~n75872;
  assign n75900 = n73167 & n73190;
  assign n75901 = n75847 & n75900;
  assign n75902 = ~n75899 & ~n75901;
  assign n75903 = n75456 & n75902;
  assign n75904 = P2_P2_REIP_REG_16_ & n75424;
  assign n75905 = P2_P2_PHYADDRPOINTER_REG_16_ & n75453;
  assign n75906 = ~n75904 & ~n75905;
  assign n75907 = ~n73190 & n75450;
  assign n75908 = n75906 & ~n75907;
  assign n75909 = ~n75889 & ~n75890;
  assign n75910 = n75898 & n75909;
  assign n75911 = ~n75903 & n75910;
  assign n14321 = ~n75908 | ~n75911;
  assign n75913 = P2_P2_REIP_REG_16_ & n75885;
  assign n75914 = ~P2_P2_REIP_REG_17_ & n75913;
  assign n75915 = P2_P2_REIP_REG_17_ & ~n75913;
  assign n75916 = ~n75914 & ~n75915;
  assign n75917 = n75447 & ~n75916;
  assign n75918 = P2_P2_EBX_REG_17_ & ~n75434;
  assign n75919 = ~P2_P2_EBX_REG_17_ & n75893;
  assign n75920 = P2_P2_EBX_REG_17_ & ~n75893;
  assign n75921 = ~n75919 & ~n75920;
  assign n75922 = n75438 & n75921;
  assign n75923 = n75436 & ~n75916;
  assign n75924 = ~n75560 & ~n75922;
  assign n75925 = ~n75923 & n75924;
  assign n75926 = n73213 & n75901;
  assign n75927 = ~n73213 & ~n75901;
  assign n75928 = ~n75926 & ~n75927;
  assign n75929 = n75456 & n75928;
  assign n75930 = P2_P2_REIP_REG_17_ & n75424;
  assign n75931 = P2_P2_PHYADDRPOINTER_REG_17_ & n75453;
  assign n75932 = ~n75930 & ~n75931;
  assign n75933 = ~n73213 & n75450;
  assign n75934 = n75932 & ~n75933;
  assign n75935 = ~n75917 & ~n75918;
  assign n75936 = n75925 & n75935;
  assign n75937 = ~n75929 & n75936;
  assign n14326 = ~n75934 | ~n75937;
  assign n75939 = P2_P2_REIP_REG_17_ & n75913;
  assign n75940 = ~P2_P2_REIP_REG_18_ & n75939;
  assign n75941 = P2_P2_REIP_REG_18_ & ~n75939;
  assign n75942 = ~n75940 & ~n75941;
  assign n75943 = n75447 & ~n75942;
  assign n75944 = P2_P2_EBX_REG_18_ & ~n75434;
  assign n75945 = P2_P2_EBX_REG_18_ & ~n75919;
  assign n75946 = ~P2_P2_EBX_REG_17_ & ~P2_P2_EBX_REG_18_;
  assign n75947 = n75893 & n75946;
  assign n75948 = ~n75945 & ~n75947;
  assign n75949 = n75438 & n75948;
  assign n75950 = n75436 & ~n75942;
  assign n75951 = ~n75560 & ~n75949;
  assign n75952 = ~n75950 & n75951;
  assign n75953 = ~n73236 & ~n75926;
  assign n75954 = n73213 & n73236;
  assign n75955 = n75901 & n75954;
  assign n75956 = ~n75953 & ~n75955;
  assign n75957 = n75456 & n75956;
  assign n75958 = P2_P2_REIP_REG_18_ & n75424;
  assign n75959 = P2_P2_PHYADDRPOINTER_REG_18_ & n75453;
  assign n75960 = ~n75958 & ~n75959;
  assign n75961 = ~n73236 & n75450;
  assign n75962 = n75960 & ~n75961;
  assign n75963 = ~n75943 & ~n75944;
  assign n75964 = n75952 & n75963;
  assign n75965 = ~n75957 & n75964;
  assign n14331 = ~n75962 | ~n75965;
  assign n75967 = P2_P2_REIP_REG_18_ & n75939;
  assign n75968 = ~P2_P2_REIP_REG_19_ & n75967;
  assign n75969 = P2_P2_REIP_REG_19_ & ~n75967;
  assign n75970 = ~n75968 & ~n75969;
  assign n75971 = n75447 & ~n75970;
  assign n75972 = P2_P2_EBX_REG_19_ & ~n75434;
  assign n75973 = ~P2_P2_EBX_REG_19_ & n75947;
  assign n75974 = P2_P2_EBX_REG_19_ & ~n75947;
  assign n75975 = ~n75973 & ~n75974;
  assign n75976 = n75438 & n75975;
  assign n75977 = n75436 & ~n75970;
  assign n75978 = ~n75560 & ~n75976;
  assign n75979 = ~n75977 & n75978;
  assign n75980 = n73259 & n75955;
  assign n75981 = ~n73259 & ~n75955;
  assign n75982 = ~n75980 & ~n75981;
  assign n75983 = n75456 & n75982;
  assign n75984 = P2_P2_REIP_REG_19_ & n75424;
  assign n75985 = P2_P2_PHYADDRPOINTER_REG_19_ & n75453;
  assign n75986 = ~n75984 & ~n75985;
  assign n75987 = ~n73259 & n75450;
  assign n75988 = n75986 & ~n75987;
  assign n75989 = ~n75971 & ~n75972;
  assign n75990 = n75979 & n75989;
  assign n75991 = ~n75983 & n75990;
  assign n14336 = ~n75988 | ~n75991;
  assign n75993 = P2_P2_REIP_REG_19_ & n75967;
  assign n75994 = ~P2_P2_REIP_REG_20_ & n75993;
  assign n75995 = P2_P2_REIP_REG_20_ & ~n75993;
  assign n75996 = ~n75994 & ~n75995;
  assign n75997 = n75447 & ~n75996;
  assign n75998 = P2_P2_EBX_REG_20_ & ~n75434;
  assign n75999 = n75436 & ~n75996;
  assign n76000 = P2_P2_EBX_REG_20_ & ~n75973;
  assign n76001 = ~P2_P2_EBX_REG_19_ & ~P2_P2_EBX_REG_20_;
  assign n76002 = n75947 & n76001;
  assign n76003 = ~n76000 & ~n76002;
  assign n76004 = n75438 & n76003;
  assign n76005 = ~n75999 & ~n76004;
  assign n76006 = ~n73282 & ~n75980;
  assign n76007 = n73259 & n73282;
  assign n76008 = n75955 & n76007;
  assign n76009 = ~n76006 & ~n76008;
  assign n76010 = n75456 & n76009;
  assign n76011 = P2_P2_REIP_REG_20_ & n75424;
  assign n76012 = P2_P2_PHYADDRPOINTER_REG_20_ & n75453;
  assign n76013 = ~n76011 & ~n76012;
  assign n76014 = ~n73282 & n75450;
  assign n76015 = n76013 & ~n76014;
  assign n76016 = ~n75997 & ~n75998;
  assign n76017 = n76005 & n76016;
  assign n76018 = ~n76010 & n76017;
  assign n14341 = ~n76015 | ~n76018;
  assign n76020 = P2_P2_REIP_REG_20_ & n75993;
  assign n76021 = ~P2_P2_REIP_REG_21_ & n76020;
  assign n76022 = P2_P2_REIP_REG_21_ & ~n76020;
  assign n76023 = ~n76021 & ~n76022;
  assign n76024 = n75447 & ~n76023;
  assign n76025 = P2_P2_EBX_REG_21_ & ~n75434;
  assign n76026 = n75436 & ~n76023;
  assign n76027 = ~P2_P2_EBX_REG_21_ & n76002;
  assign n76028 = P2_P2_EBX_REG_21_ & ~n76002;
  assign n76029 = ~n76027 & ~n76028;
  assign n76030 = n75438 & n76029;
  assign n76031 = ~n76026 & ~n76030;
  assign n76032 = n73305 & n76008;
  assign n76033 = ~n73305 & ~n76008;
  assign n76034 = ~n76032 & ~n76033;
  assign n76035 = n75456 & n76034;
  assign n76036 = P2_P2_REIP_REG_21_ & n75424;
  assign n76037 = P2_P2_PHYADDRPOINTER_REG_21_ & n75453;
  assign n76038 = ~n76036 & ~n76037;
  assign n76039 = ~n73305 & n75450;
  assign n76040 = n76038 & ~n76039;
  assign n76041 = ~n76024 & ~n76025;
  assign n76042 = n76031 & n76041;
  assign n76043 = ~n76035 & n76042;
  assign n14346 = ~n76040 | ~n76043;
  assign n76045 = P2_P2_REIP_REG_21_ & n76020;
  assign n76046 = ~P2_P2_REIP_REG_22_ & n76045;
  assign n76047 = P2_P2_REIP_REG_22_ & ~n76045;
  assign n76048 = ~n76046 & ~n76047;
  assign n76049 = n75447 & ~n76048;
  assign n76050 = P2_P2_EBX_REG_22_ & ~n75434;
  assign n76051 = n75436 & ~n76048;
  assign n76052 = P2_P2_EBX_REG_22_ & ~n76027;
  assign n76053 = ~P2_P2_EBX_REG_21_ & ~P2_P2_EBX_REG_22_;
  assign n76054 = n76002 & n76053;
  assign n76055 = ~n76052 & ~n76054;
  assign n76056 = n75438 & n76055;
  assign n76057 = ~n76051 & ~n76056;
  assign n76058 = ~n73329 & ~n76032;
  assign n76059 = n73305 & n73329;
  assign n76060 = n76008 & n76059;
  assign n76061 = ~n76058 & ~n76060;
  assign n76062 = n75456 & n76061;
  assign n76063 = P2_P2_REIP_REG_22_ & n75424;
  assign n76064 = P2_P2_PHYADDRPOINTER_REG_22_ & n75453;
  assign n76065 = ~n76063 & ~n76064;
  assign n76066 = ~n73329 & n75450;
  assign n76067 = n76065 & ~n76066;
  assign n76068 = ~n76049 & ~n76050;
  assign n76069 = n76057 & n76068;
  assign n76070 = ~n76062 & n76069;
  assign n14351 = ~n76067 | ~n76070;
  assign n76072 = P2_P2_REIP_REG_22_ & n76045;
  assign n76073 = ~P2_P2_REIP_REG_23_ & n76072;
  assign n76074 = P2_P2_REIP_REG_23_ & ~n76072;
  assign n76075 = ~n76073 & ~n76074;
  assign n76076 = n75447 & ~n76075;
  assign n76077 = P2_P2_EBX_REG_23_ & ~n75434;
  assign n76078 = n75436 & ~n76075;
  assign n76079 = ~P2_P2_EBX_REG_23_ & n76054;
  assign n76080 = P2_P2_EBX_REG_23_ & ~n76054;
  assign n76081 = ~n76079 & ~n76080;
  assign n76082 = n75438 & n76081;
  assign n76083 = ~n76078 & ~n76082;
  assign n76084 = n73352 & n76060;
  assign n76085 = ~n73352 & ~n76060;
  assign n76086 = ~n76084 & ~n76085;
  assign n76087 = n75456 & n76086;
  assign n76088 = P2_P2_REIP_REG_23_ & n75424;
  assign n76089 = P2_P2_PHYADDRPOINTER_REG_23_ & n75453;
  assign n76090 = ~n76088 & ~n76089;
  assign n76091 = ~n73352 & n75450;
  assign n76092 = n76090 & ~n76091;
  assign n76093 = ~n76076 & ~n76077;
  assign n76094 = n76083 & n76093;
  assign n76095 = ~n76087 & n76094;
  assign n14356 = ~n76092 | ~n76095;
  assign n76097 = P2_P2_REIP_REG_23_ & n76072;
  assign n76098 = ~P2_P2_REIP_REG_24_ & n76097;
  assign n76099 = P2_P2_REIP_REG_24_ & ~n76097;
  assign n76100 = ~n76098 & ~n76099;
  assign n76101 = n75447 & ~n76100;
  assign n76102 = P2_P2_EBX_REG_24_ & ~n75434;
  assign n76103 = n75436 & ~n76100;
  assign n76104 = P2_P2_EBX_REG_24_ & ~n76079;
  assign n76105 = ~P2_P2_EBX_REG_23_ & ~P2_P2_EBX_REG_24_;
  assign n76106 = n76054 & n76105;
  assign n76107 = ~n76104 & ~n76106;
  assign n76108 = n75438 & n76107;
  assign n76109 = ~n76103 & ~n76108;
  assign n76110 = ~n73375 & ~n76084;
  assign n76111 = n73352 & n73375;
  assign n76112 = n76060 & n76111;
  assign n76113 = ~n76110 & ~n76112;
  assign n76114 = n75456 & n76113;
  assign n76115 = P2_P2_REIP_REG_24_ & n75424;
  assign n76116 = P2_P2_PHYADDRPOINTER_REG_24_ & n75453;
  assign n76117 = ~n76115 & ~n76116;
  assign n76118 = ~n73375 & n75450;
  assign n76119 = n76117 & ~n76118;
  assign n76120 = ~n76101 & ~n76102;
  assign n76121 = n76109 & n76120;
  assign n76122 = ~n76114 & n76121;
  assign n14361 = ~n76119 | ~n76122;
  assign n76124 = P2_P2_REIP_REG_24_ & n76097;
  assign n76125 = ~P2_P2_REIP_REG_25_ & n76124;
  assign n76126 = P2_P2_REIP_REG_25_ & ~n76124;
  assign n76127 = ~n76125 & ~n76126;
  assign n76128 = n75447 & ~n76127;
  assign n76129 = P2_P2_EBX_REG_25_ & ~n75434;
  assign n76130 = n75436 & ~n76127;
  assign n76131 = ~P2_P2_EBX_REG_25_ & n76106;
  assign n76132 = P2_P2_EBX_REG_25_ & ~n76106;
  assign n76133 = ~n76131 & ~n76132;
  assign n76134 = n75438 & n76133;
  assign n76135 = ~n76130 & ~n76134;
  assign n76136 = n73398 & n76112;
  assign n76137 = ~n73398 & ~n76112;
  assign n76138 = ~n76136 & ~n76137;
  assign n76139 = n75456 & n76138;
  assign n76140 = P2_P2_REIP_REG_25_ & n75424;
  assign n76141 = P2_P2_PHYADDRPOINTER_REG_25_ & n75453;
  assign n76142 = ~n76140 & ~n76141;
  assign n76143 = ~n73398 & n75450;
  assign n76144 = n76142 & ~n76143;
  assign n76145 = ~n76128 & ~n76129;
  assign n76146 = n76135 & n76145;
  assign n76147 = ~n76139 & n76146;
  assign n14366 = ~n76144 | ~n76147;
  assign n76149 = P2_P2_REIP_REG_25_ & n76124;
  assign n76150 = ~P2_P2_REIP_REG_26_ & n76149;
  assign n76151 = P2_P2_REIP_REG_26_ & ~n76149;
  assign n76152 = ~n76150 & ~n76151;
  assign n76153 = n75447 & ~n76152;
  assign n76154 = P2_P2_EBX_REG_26_ & ~n75434;
  assign n76155 = n75436 & ~n76152;
  assign n76156 = P2_P2_EBX_REG_26_ & ~n76131;
  assign n76157 = ~P2_P2_EBX_REG_25_ & ~P2_P2_EBX_REG_26_;
  assign n76158 = n76106 & n76157;
  assign n76159 = ~n76156 & ~n76158;
  assign n76160 = n75438 & n76159;
  assign n76161 = ~n76155 & ~n76160;
  assign n76162 = ~n73421 & ~n76136;
  assign n76163 = n73398 & n73421;
  assign n76164 = n76112 & n76163;
  assign n76165 = ~n76162 & ~n76164;
  assign n76166 = n75456 & n76165;
  assign n76167 = P2_P2_REIP_REG_26_ & n75424;
  assign n76168 = P2_P2_PHYADDRPOINTER_REG_26_ & n75453;
  assign n76169 = ~n76167 & ~n76168;
  assign n76170 = ~n73421 & n75450;
  assign n76171 = n76169 & ~n76170;
  assign n76172 = ~n76153 & ~n76154;
  assign n76173 = n76161 & n76172;
  assign n76174 = ~n76166 & n76173;
  assign n14371 = ~n76171 | ~n76174;
  assign n76176 = P2_P2_REIP_REG_26_ & n76149;
  assign n76177 = ~P2_P2_REIP_REG_27_ & n76176;
  assign n76178 = P2_P2_REIP_REG_27_ & ~n76176;
  assign n76179 = ~n76177 & ~n76178;
  assign n76180 = n75447 & ~n76179;
  assign n76181 = P2_P2_EBX_REG_27_ & ~n75434;
  assign n76182 = n75436 & ~n76179;
  assign n76183 = ~P2_P2_EBX_REG_27_ & n76158;
  assign n76184 = P2_P2_EBX_REG_27_ & ~n76158;
  assign n76185 = ~n76183 & ~n76184;
  assign n76186 = n75438 & n76185;
  assign n76187 = ~n76182 & ~n76186;
  assign n76188 = n73444 & n76164;
  assign n76189 = ~n73444 & ~n76164;
  assign n76190 = ~n76188 & ~n76189;
  assign n76191 = n75456 & n76190;
  assign n76192 = P2_P2_REIP_REG_27_ & n75424;
  assign n76193 = P2_P2_PHYADDRPOINTER_REG_27_ & n75453;
  assign n76194 = ~n76192 & ~n76193;
  assign n76195 = ~n73444 & n75450;
  assign n76196 = n76194 & ~n76195;
  assign n76197 = ~n76180 & ~n76181;
  assign n76198 = n76187 & n76197;
  assign n76199 = ~n76191 & n76198;
  assign n14376 = ~n76196 | ~n76199;
  assign n76201 = P2_P2_REIP_REG_27_ & n76176;
  assign n76202 = ~P2_P2_REIP_REG_28_ & n76201;
  assign n76203 = P2_P2_REIP_REG_28_ & ~n76201;
  assign n76204 = ~n76202 & ~n76203;
  assign n76205 = n75447 & ~n76204;
  assign n76206 = P2_P2_EBX_REG_28_ & ~n75434;
  assign n76207 = n75436 & ~n76204;
  assign n76208 = P2_P2_EBX_REG_28_ & ~n76183;
  assign n76209 = ~P2_P2_EBX_REG_27_ & ~P2_P2_EBX_REG_28_;
  assign n76210 = n76158 & n76209;
  assign n76211 = ~n76208 & ~n76210;
  assign n76212 = n75438 & n76211;
  assign n76213 = ~n76207 & ~n76212;
  assign n76214 = ~n73468 & ~n76188;
  assign n76215 = n73444 & n73468;
  assign n76216 = n76164 & n76215;
  assign n76217 = ~n76214 & ~n76216;
  assign n76218 = n75456 & n76217;
  assign n76219 = P2_P2_REIP_REG_28_ & n75424;
  assign n76220 = P2_P2_PHYADDRPOINTER_REG_28_ & n75453;
  assign n76221 = ~n76219 & ~n76220;
  assign n76222 = ~n73468 & n75450;
  assign n76223 = n76221 & ~n76222;
  assign n76224 = ~n76205 & ~n76206;
  assign n76225 = n76213 & n76224;
  assign n76226 = ~n76218 & n76225;
  assign n14381 = ~n76223 | ~n76226;
  assign n76228 = P2_P2_REIP_REG_28_ & n76201;
  assign n76229 = ~P2_P2_REIP_REG_29_ & n76228;
  assign n76230 = P2_P2_REIP_REG_29_ & ~n76228;
  assign n76231 = ~n76229 & ~n76230;
  assign n76232 = n75447 & ~n76231;
  assign n76233 = P2_P2_EBX_REG_29_ & ~n75434;
  assign n76234 = n75436 & ~n76231;
  assign n76235 = P2_P2_EBX_REG_29_ & ~n76210;
  assign n76236 = ~P2_P2_EBX_REG_29_ & n76210;
  assign n76237 = ~n76235 & ~n76236;
  assign n76238 = n75438 & n76237;
  assign n76239 = ~n76234 & ~n76238;
  assign n76240 = ~n73491 & ~n76216;
  assign n76241 = n73491 & n76216;
  assign n76242 = ~n76240 & ~n76241;
  assign n76243 = n75456 & n76242;
  assign n76244 = P2_P2_REIP_REG_29_ & n75424;
  assign n76245 = P2_P2_PHYADDRPOINTER_REG_29_ & n75453;
  assign n76246 = ~n76244 & ~n76245;
  assign n76247 = ~n73491 & n75450;
  assign n76248 = n76246 & ~n76247;
  assign n76249 = ~n76232 & ~n76233;
  assign n76250 = n76239 & n76249;
  assign n76251 = ~n76243 & n76250;
  assign n14386 = ~n76248 | ~n76251;
  assign n76253 = P2_P2_REIP_REG_29_ & n76228;
  assign n76254 = ~P2_P2_REIP_REG_30_ & n76253;
  assign n76255 = P2_P2_REIP_REG_30_ & ~n76253;
  assign n76256 = ~n76254 & ~n76255;
  assign n76257 = n75447 & ~n76256;
  assign n76258 = P2_P2_EBX_REG_30_ & ~n75434;
  assign n76259 = n75436 & ~n76256;
  assign n76260 = ~P2_P2_EBX_REG_30_ & n76236;
  assign n76261 = P2_P2_EBX_REG_30_ & ~n76236;
  assign n76262 = ~n76260 & ~n76261;
  assign n76263 = n75438 & n76262;
  assign n76264 = ~n76259 & ~n76263;
  assign n76265 = n73514 & n76241;
  assign n76266 = ~n73514 & ~n76241;
  assign n76267 = ~n76265 & ~n76266;
  assign n76268 = n75456 & n76267;
  assign n76269 = P2_P2_REIP_REG_30_ & n75424;
  assign n76270 = P2_P2_PHYADDRPOINTER_REG_30_ & n75453;
  assign n76271 = ~n76269 & ~n76270;
  assign n76272 = ~n73514 & n75450;
  assign n76273 = n76271 & ~n76272;
  assign n76274 = ~n76257 & ~n76258;
  assign n76275 = n76264 & n76274;
  assign n76276 = ~n76268 & n76275;
  assign n14391 = ~n76273 | ~n76276;
  assign n76278 = ~n73537 & n76265;
  assign n76279 = n73537 & ~n76265;
  assign n76280 = ~n76278 & ~n76279;
  assign n76281 = ~n73537 & n75450;
  assign n76282 = n76280 & ~n76281;
  assign n76283 = P2_P2_EBX_REG_31_ & ~n75434;
  assign n76284 = P2_P2_EBX_REG_31_ & n76260;
  assign n76285 = ~P2_P2_EBX_REG_31_ & ~n76260;
  assign n76286 = ~n76284 & ~n76285;
  assign n76287 = n75438 & ~n76286;
  assign n76288 = P2_P2_REIP_REG_30_ & n76253;
  assign n76289 = ~P2_P2_REIP_REG_31_ & n76288;
  assign n76290 = P2_P2_REIP_REG_31_ & ~n76288;
  assign n76291 = ~n76289 & ~n76290;
  assign n76292 = n75436 & ~n76291;
  assign n76293 = P2_P2_PHYADDRPOINTER_REG_31_ & n75453;
  assign n76294 = P2_P2_REIP_REG_31_ & n75424;
  assign n76295 = ~n76293 & ~n76294;
  assign n76296 = n75447 & ~n76291;
  assign n76297 = n76295 & ~n76296;
  assign n76298 = ~n76283 & ~n76287;
  assign n76299 = ~n76292 & n76298;
  assign n76300 = n76297 & n76299;
  assign n76301 = n76282 & n76300;
  assign n76302 = ~n75456 & ~n76281;
  assign n76303 = n76300 & n76302;
  assign n14396 = ~n76301 & ~n76303;
  assign n76305 = ~P2_P2_DATAWIDTH_REG_1_ & ~P2_P2_REIP_REG_1_;
  assign n76306 = ~P2_P2_DATAWIDTH_REG_30_ & ~P2_P2_DATAWIDTH_REG_31_;
  assign n76307 = P2_P2_DATAWIDTH_REG_0_ & P2_P2_DATAWIDTH_REG_1_;
  assign n76308 = ~P2_P2_DATAWIDTH_REG_28_ & ~P2_P2_DATAWIDTH_REG_29_;
  assign n76309 = ~P2_P2_DATAWIDTH_REG_26_ & ~P2_P2_DATAWIDTH_REG_27_;
  assign n76310 = n76306 & ~n76307;
  assign n76311 = n76308 & n76310;
  assign n76312 = n76309 & n76311;
  assign n76313 = ~P2_P2_DATAWIDTH_REG_22_ & ~P2_P2_DATAWIDTH_REG_23_;
  assign n76314 = ~P2_P2_DATAWIDTH_REG_24_ & n76313;
  assign n76315 = ~P2_P2_DATAWIDTH_REG_25_ & n76314;
  assign n76316 = ~P2_P2_DATAWIDTH_REG_18_ & ~P2_P2_DATAWIDTH_REG_19_;
  assign n76317 = ~P2_P2_DATAWIDTH_REG_20_ & n76316;
  assign n76318 = ~P2_P2_DATAWIDTH_REG_21_ & n76317;
  assign n76319 = n76315 & n76318;
  assign n76320 = ~P2_P2_DATAWIDTH_REG_14_ & ~P2_P2_DATAWIDTH_REG_15_;
  assign n76321 = ~P2_P2_DATAWIDTH_REG_16_ & n76320;
  assign n76322 = ~P2_P2_DATAWIDTH_REG_17_ & n76321;
  assign n76323 = ~P2_P2_DATAWIDTH_REG_10_ & ~P2_P2_DATAWIDTH_REG_11_;
  assign n76324 = ~P2_P2_DATAWIDTH_REG_12_ & n76323;
  assign n76325 = ~P2_P2_DATAWIDTH_REG_13_ & n76324;
  assign n76326 = n76322 & n76325;
  assign n76327 = ~P2_P2_DATAWIDTH_REG_6_ & ~P2_P2_DATAWIDTH_REG_7_;
  assign n76328 = ~P2_P2_DATAWIDTH_REG_8_ & n76327;
  assign n76329 = ~P2_P2_DATAWIDTH_REG_9_ & n76328;
  assign n76330 = ~P2_P2_DATAWIDTH_REG_2_ & ~P2_P2_DATAWIDTH_REG_3_;
  assign n76331 = ~P2_P2_DATAWIDTH_REG_4_ & n76330;
  assign n76332 = ~P2_P2_DATAWIDTH_REG_5_ & n76331;
  assign n76333 = n76329 & n76332;
  assign n76334 = n76312 & n76319;
  assign n76335 = n76326 & n76334;
  assign n76336 = n76333 & n76335;
  assign n76337 = n76305 & n76336;
  assign n76338 = P2_P2_BYTEENABLE_REG_3_ & ~n76336;
  assign n76339 = ~P2_P2_DATAWIDTH_REG_0_ & ~P2_P2_REIP_REG_0_;
  assign n76340 = ~P2_P2_DATAWIDTH_REG_1_ & n76339;
  assign n76341 = n76336 & n76340;
  assign n76342 = ~n76337 & ~n76338;
  assign n14401 = n76341 | ~n76342;
  assign n76344 = P2_P2_REIP_REG_0_ & P2_P2_REIP_REG_1_;
  assign n76345 = P2_P2_DATAWIDTH_REG_0_ & ~P2_P2_REIP_REG_0_;
  assign n76346 = ~P2_P2_DATAWIDTH_REG_0_ & ~P2_P2_DATAWIDTH_REG_1_;
  assign n76347 = ~n76345 & ~n76346;
  assign n76348 = ~P2_P2_REIP_REG_1_ & ~n76347;
  assign n76349 = ~n76344 & ~n76348;
  assign n76350 = n76336 & ~n76349;
  assign n76351 = P2_P2_BYTEENABLE_REG_2_ & ~n76336;
  assign n14406 = n76350 | n76351;
  assign n76353 = P2_P2_REIP_REG_1_ & n76336;
  assign n76354 = P2_P2_BYTEENABLE_REG_1_ & ~n76336;
  assign n76355 = ~n76353 & ~n76354;
  assign n14411 = n76341 | ~n76355;
  assign n76357 = ~P2_P2_REIP_REG_0_ & ~P2_P2_REIP_REG_1_;
  assign n76358 = n76336 & ~n76357;
  assign n76359 = P2_P2_BYTEENABLE_REG_0_ & ~n76336;
  assign n14416 = n76358 | n76359;
  assign n76361 = P2_P2_W_R_N_REG & ~n67372;
  assign n76362 = ~P2_P2_READREQUEST_REG & n67372;
  assign n14421 = n76361 | n76362;
  assign n76364 = n68036 & n68268;
  assign n76365 = ~n67984 & n68268;
  assign n76366 = P2_P2_FLUSH_REG & ~n76365;
  assign n14426 = n76364 | n76366;
  assign n76368 = P2_P2_MORE_REG & ~n76365;
  assign n76369 = ~n68030 & n76365;
  assign n14431 = n76368 | n76369;
  assign n76371 = BS & ~n67589;
  assign n76372 = P2_P2_STATEBS16_REG & n67589;
  assign n76373 = ~P2_P2_STATE_REG_0_ & n67544;
  assign n76374 = ~n76371 & ~n76372;
  assign n14436 = n76373 | ~n76374;
  assign n76376 = ~n67914 & ~n67987;
  assign n76377 = ~n67632 & ~n76376;
  assign n76378 = ~P2_P2_STATEBS16_REG & n67914;
  assign n76379 = ~n67541 & ~n76378;
  assign n76380 = P2_P2_STATE2_REG_2_ & ~n76377;
  assign n76381 = n76379 & n76380;
  assign n76382 = P2_P2_STATE2_REG_0_ & ~n76381;
  assign n76383 = ~n68284 & ~n76382;
  assign n76384 = ~n67541 & n67626;
  assign n76385 = ~n68274 & ~n76384;
  assign n76386 = ~P2_P2_STATE2_REG_0_ & ~n76385;
  assign n76387 = ~n68346 & ~n76386;
  assign n76388 = ~n75423 & n76387;
  assign n76389 = ~n76383 & ~n76388;
  assign n76390 = P2_P2_REQUESTPENDING_REG & n76388;
  assign n14441 = n76389 | n76390;
  assign n76392 = P2_P2_D_C_N_REG & ~n67372;
  assign n76393 = ~P2_P2_CODEFETCH_REG & n67372;
  assign n76394 = ~n76392 & ~n76393;
  assign n14446 = n76373 | ~n76394;
  assign n76396 = P2_P2_MEMORYFETCH_REG & n67372;
  assign n76397 = P2_P2_M_IO_N_REG & ~n67372;
  assign n14451 = n76396 | n76397;
  assign n76399 = P2_P2_STATE2_REG_0_ & n69953;
  assign n76400 = n67983 & n68268;
  assign n76401 = P2_P2_CODEFETCH_REG & ~n76400;
  assign n14456 = n76399 | n76401;
  assign n76403 = P2_P2_STATE_REG_0_ & P2_P2_ADS_N_REG;
  assign n14461 = ~n67589 | n76403;
  assign n76405 = P2_P2_STATE2_REG_2_ & ~n67996;
  assign n76406 = ~n67991 & n76405;
  assign n76407 = ~n69953 & ~n75423;
  assign n76408 = ~n76406 & ~n76407;
  assign n76409 = P2_P2_READREQUEST_REG & n76407;
  assign n14466 = n76408 | n76409;
  assign n76411 = P2_P2_STATE2_REG_2_ & n67913;
  assign n76412 = ~n76407 & ~n76411;
  assign n76413 = P2_P2_MEMORYFETCH_REG & n76407;
  assign n14471 = n76412 | n76413;
  assign n76415 = P2_P1_STATE_REG_1_ & ~P2_P1_STATE_REG_0_;
  assign n76416 = P2_P1_BYTEENABLE_REG_3_ & n76415;
  assign n76417 = P2_P1_BE_N_REG_3_ & ~n76415;
  assign n14476 = n76416 | n76417;
  assign n76419 = P2_P1_BYTEENABLE_REG_2_ & n76415;
  assign n76420 = P2_P1_BE_N_REG_2_ & ~n76415;
  assign n14481 = n76419 | n76420;
  assign n76422 = P2_P1_BYTEENABLE_REG_1_ & n76415;
  assign n76423 = P2_P1_BE_N_REG_1_ & ~n76415;
  assign n14486 = n76422 | n76423;
  assign n76425 = P2_P1_BYTEENABLE_REG_0_ & n76415;
  assign n76426 = P2_P1_BE_N_REG_0_ & ~n76415;
  assign n14491 = n76425 | n76426;
  assign n76428 = P2_P1_STATE_REG_2_ & n76415;
  assign n76429 = P2_P1_REIP_REG_30_ & n76428;
  assign n76430 = ~P2_P1_STATE_REG_2_ & n76415;
  assign n76431 = P2_P1_REIP_REG_31_ & n76430;
  assign n76432 = P2_P1_ADDRESS_REG_29_ & ~n76415;
  assign n76433 = ~n76429 & ~n76431;
  assign n14496 = n76432 | ~n76433;
  assign n76435 = P2_P1_REIP_REG_29_ & n76428;
  assign n76436 = P2_P1_REIP_REG_30_ & n76430;
  assign n76437 = P2_P1_ADDRESS_REG_28_ & ~n76415;
  assign n76438 = ~n76435 & ~n76436;
  assign n14501 = n76437 | ~n76438;
  assign n76440 = P2_P1_REIP_REG_28_ & n76428;
  assign n76441 = P2_P1_REIP_REG_29_ & n76430;
  assign n76442 = P2_P1_ADDRESS_REG_27_ & ~n76415;
  assign n76443 = ~n76440 & ~n76441;
  assign n14506 = n76442 | ~n76443;
  assign n76445 = P2_P1_REIP_REG_27_ & n76428;
  assign n76446 = P2_P1_REIP_REG_28_ & n76430;
  assign n76447 = P2_P1_ADDRESS_REG_26_ & ~n76415;
  assign n76448 = ~n76445 & ~n76446;
  assign n14511 = n76447 | ~n76448;
  assign n76450 = P2_P1_REIP_REG_26_ & n76428;
  assign n76451 = P2_P1_REIP_REG_27_ & n76430;
  assign n76452 = P2_P1_ADDRESS_REG_25_ & ~n76415;
  assign n76453 = ~n76450 & ~n76451;
  assign n14516 = n76452 | ~n76453;
  assign n76455 = P2_P1_REIP_REG_25_ & n76428;
  assign n76456 = P2_P1_REIP_REG_26_ & n76430;
  assign n76457 = P2_P1_ADDRESS_REG_24_ & ~n76415;
  assign n76458 = ~n76455 & ~n76456;
  assign n14521 = n76457 | ~n76458;
  assign n76460 = P2_P1_REIP_REG_24_ & n76428;
  assign n76461 = P2_P1_REIP_REG_25_ & n76430;
  assign n76462 = P2_P1_ADDRESS_REG_23_ & ~n76415;
  assign n76463 = ~n76460 & ~n76461;
  assign n14526 = n76462 | ~n76463;
  assign n76465 = P2_P1_REIP_REG_23_ & n76428;
  assign n76466 = P2_P1_REIP_REG_24_ & n76430;
  assign n76467 = P2_P1_ADDRESS_REG_22_ & ~n76415;
  assign n76468 = ~n76465 & ~n76466;
  assign n14531 = n76467 | ~n76468;
  assign n76470 = P2_P1_REIP_REG_22_ & n76428;
  assign n76471 = P2_P1_REIP_REG_23_ & n76430;
  assign n76472 = P2_P1_ADDRESS_REG_21_ & ~n76415;
  assign n76473 = ~n76470 & ~n76471;
  assign n14536 = n76472 | ~n76473;
  assign n76475 = P2_P1_REIP_REG_21_ & n76428;
  assign n76476 = P2_P1_REIP_REG_22_ & n76430;
  assign n76477 = P2_P1_ADDRESS_REG_20_ & ~n76415;
  assign n76478 = ~n76475 & ~n76476;
  assign n14541 = n76477 | ~n76478;
  assign n76480 = P2_P1_REIP_REG_20_ & n76428;
  assign n76481 = P2_P1_REIP_REG_21_ & n76430;
  assign n76482 = P2_P1_ADDRESS_REG_19_ & ~n76415;
  assign n76483 = ~n76480 & ~n76481;
  assign n14546 = n76482 | ~n76483;
  assign n76485 = P2_P1_REIP_REG_19_ & n76428;
  assign n76486 = P2_P1_REIP_REG_20_ & n76430;
  assign n76487 = P2_P1_ADDRESS_REG_18_ & ~n76415;
  assign n76488 = ~n76485 & ~n76486;
  assign n14551 = n76487 | ~n76488;
  assign n76490 = P2_P1_REIP_REG_18_ & n76428;
  assign n76491 = P2_P1_REIP_REG_19_ & n76430;
  assign n76492 = P2_P1_ADDRESS_REG_17_ & ~n76415;
  assign n76493 = ~n76490 & ~n76491;
  assign n14556 = n76492 | ~n76493;
  assign n76495 = P2_P1_REIP_REG_17_ & n76428;
  assign n76496 = P2_P1_REIP_REG_18_ & n76430;
  assign n76497 = P2_P1_ADDRESS_REG_16_ & ~n76415;
  assign n76498 = ~n76495 & ~n76496;
  assign n14561 = n76497 | ~n76498;
  assign n76500 = P2_P1_REIP_REG_16_ & n76428;
  assign n76501 = P2_P1_REIP_REG_17_ & n76430;
  assign n76502 = P2_P1_ADDRESS_REG_15_ & ~n76415;
  assign n76503 = ~n76500 & ~n76501;
  assign n14566 = n76502 | ~n76503;
  assign n76505 = P2_P1_REIP_REG_15_ & n76428;
  assign n76506 = P2_P1_REIP_REG_16_ & n76430;
  assign n76507 = P2_P1_ADDRESS_REG_14_ & ~n76415;
  assign n76508 = ~n76505 & ~n76506;
  assign n14571 = n76507 | ~n76508;
  assign n76510 = P2_P1_REIP_REG_14_ & n76428;
  assign n76511 = P2_P1_REIP_REG_15_ & n76430;
  assign n76512 = P2_P1_ADDRESS_REG_13_ & ~n76415;
  assign n76513 = ~n76510 & ~n76511;
  assign n14576 = n76512 | ~n76513;
  assign n76515 = P2_P1_REIP_REG_13_ & n76428;
  assign n76516 = P2_P1_REIP_REG_14_ & n76430;
  assign n76517 = P2_P1_ADDRESS_REG_12_ & ~n76415;
  assign n76518 = ~n76515 & ~n76516;
  assign n14581 = n76517 | ~n76518;
  assign n76520 = P2_P1_REIP_REG_12_ & n76428;
  assign n76521 = P2_P1_REIP_REG_13_ & n76430;
  assign n76522 = P2_P1_ADDRESS_REG_11_ & ~n76415;
  assign n76523 = ~n76520 & ~n76521;
  assign n14586 = n76522 | ~n76523;
  assign n76525 = P2_P1_REIP_REG_11_ & n76428;
  assign n76526 = P2_P1_REIP_REG_12_ & n76430;
  assign n76527 = P2_P1_ADDRESS_REG_10_ & ~n76415;
  assign n76528 = ~n76525 & ~n76526;
  assign n14591 = n76527 | ~n76528;
  assign n76530 = P2_P1_REIP_REG_10_ & n76428;
  assign n76531 = P2_P1_REIP_REG_11_ & n76430;
  assign n76532 = P2_P1_ADDRESS_REG_9_ & ~n76415;
  assign n76533 = ~n76530 & ~n76531;
  assign n14596 = n76532 | ~n76533;
  assign n76535 = P2_P1_REIP_REG_9_ & n76428;
  assign n76536 = P2_P1_REIP_REG_10_ & n76430;
  assign n76537 = P2_P1_ADDRESS_REG_8_ & ~n76415;
  assign n76538 = ~n76535 & ~n76536;
  assign n14601 = n76537 | ~n76538;
  assign n76540 = P2_P1_REIP_REG_8_ & n76428;
  assign n76541 = P2_P1_REIP_REG_9_ & n76430;
  assign n76542 = P2_P1_ADDRESS_REG_7_ & ~n76415;
  assign n76543 = ~n76540 & ~n76541;
  assign n14606 = n76542 | ~n76543;
  assign n76545 = P2_P1_REIP_REG_7_ & n76428;
  assign n76546 = P2_P1_REIP_REG_8_ & n76430;
  assign n76547 = P2_P1_ADDRESS_REG_6_ & ~n76415;
  assign n76548 = ~n76545 & ~n76546;
  assign n14611 = n76547 | ~n76548;
  assign n76550 = P2_P1_REIP_REG_6_ & n76428;
  assign n76551 = P2_P1_REIP_REG_7_ & n76430;
  assign n76552 = P2_P1_ADDRESS_REG_5_ & ~n76415;
  assign n76553 = ~n76550 & ~n76551;
  assign n14616 = n76552 | ~n76553;
  assign n76555 = P2_P1_REIP_REG_5_ & n76428;
  assign n76556 = P2_P1_REIP_REG_6_ & n76430;
  assign n76557 = P2_P1_ADDRESS_REG_4_ & ~n76415;
  assign n76558 = ~n76555 & ~n76556;
  assign n14621 = n76557 | ~n76558;
  assign n76560 = P2_P1_REIP_REG_4_ & n76428;
  assign n76561 = P2_P1_REIP_REG_5_ & n76430;
  assign n76562 = P2_P1_ADDRESS_REG_3_ & ~n76415;
  assign n76563 = ~n76560 & ~n76561;
  assign n14626 = n76562 | ~n76563;
  assign n76565 = P2_P1_REIP_REG_3_ & n76428;
  assign n76566 = P2_P1_REIP_REG_4_ & n76430;
  assign n76567 = P2_P1_ADDRESS_REG_2_ & ~n76415;
  assign n76568 = ~n76565 & ~n76566;
  assign n14631 = n76567 | ~n76568;
  assign n76570 = P2_P1_REIP_REG_2_ & n76428;
  assign n76571 = P2_P1_REIP_REG_3_ & n76430;
  assign n76572 = P2_P1_ADDRESS_REG_1_ & ~n76415;
  assign n76573 = ~n76570 & ~n76571;
  assign n14636 = n76572 | ~n76573;
  assign n76575 = P2_P1_REIP_REG_1_ & n76428;
  assign n76576 = P2_P1_REIP_REG_2_ & n76430;
  assign n76577 = P2_P1_ADDRESS_REG_0_ & ~n76415;
  assign n76578 = ~n76575 & ~n76576;
  assign n14641 = n76577 | ~n76578;
  assign n76580 = ~P2_P1_STATE_REG_2_ & P2_P1_STATE_REG_1_;
  assign n76581 = NA & n76580;
  assign n76582 = P2_P1_STATE_REG_0_ & ~n76581;
  assign n76583 = ~HOLD & ~P2_P1_REQUESTPENDING_REG;
  assign n76584 = P2_READY11_REG & P1_P1_ADS_N_REG;
  assign n76585 = ~n76583 & n76584;
  assign n76586 = n76580 & n76585;
  assign n76587 = ~P2_P1_STATE_REG_2_ & ~P2_P1_STATE_REG_1_;
  assign n76588 = HOLD & ~P2_P1_REQUESTPENDING_REG;
  assign n76589 = n76587 & n76588;
  assign n76590 = ~n76586 & ~n76589;
  assign n76591 = n76582 & ~n76590;
  assign n76592 = ~n76428 & ~n76591;
  assign n76593 = ~HOLD & P2_P1_REQUESTPENDING_REG;
  assign n76594 = P2_P1_STATE_REG_0_ & ~n76593;
  assign n76595 = ~n76583 & n76594;
  assign n76596 = ~NA & ~P2_P1_STATE_REG_0_;
  assign n76597 = n76583 & ~n76584;
  assign n76598 = ~n76584 & n76593;
  assign n76599 = P2_P1_STATE_REG_1_ & ~n76597;
  assign n76600 = ~n76598 & n76599;
  assign n76601 = ~n76595 & ~n76596;
  assign n76602 = ~n76600 & n76601;
  assign n76603 = P2_P1_STATE_REG_2_ & ~n76602;
  assign n14646 = ~n76592 | n76603;
  assign n76605 = P2_P1_STATE_REG_2_ & ~n76594;
  assign n76606 = P2_P1_STATE_REG_0_ & P2_P1_REQUESTPENDING_REG;
  assign n76607 = ~P2_P1_STATE_REG_2_ & n76606;
  assign n76608 = ~n76605 & ~n76607;
  assign n76609 = ~P2_P1_STATE_REG_1_ & ~n76608;
  assign n76610 = HOLD & ~n76584;
  assign n76611 = P2_P1_STATE_REG_0_ & ~n76610;
  assign n76612 = P2_P1_STATE_REG_2_ & ~n76611;
  assign n76613 = ~n76597 & ~n76612;
  assign n76614 = P2_P1_STATE_REG_1_ & n76613;
  assign n76615 = n76415 & n76584;
  assign n76616 = ~n76430 & ~n76615;
  assign n76617 = ~n76609 & ~n76614;
  assign n14651 = ~n76616 | ~n76617;
  assign n76619 = P2_P1_STATE_REG_1_ & ~n76598;
  assign n76620 = n76606 & ~n76619;
  assign n76621 = ~P2_P1_STATE_REG_2_ & ~n76620;
  assign n76622 = P2_P1_STATE_REG_2_ & n76594;
  assign n76623 = NA & ~P2_P1_STATE_REG_0_;
  assign n76624 = P2_P1_STATE_REG_2_ & ~n76593;
  assign n76625 = ~n76623 & ~n76624;
  assign n76626 = ~P2_P1_STATE_REG_1_ & ~n76625;
  assign n76627 = ~n76621 & ~n76622;
  assign n14656 = n76626 | ~n76627;
  assign n76629 = ~BS & ~n76587;
  assign n76630 = P2_P1_STATE_REG_0_ & n76580;
  assign n76631 = ~P2_P1_STATE_REG_1_ & ~P2_P1_STATE_REG_0_;
  assign n76632 = ~n76630 & ~n76631;
  assign n76633 = n76629 & ~n76632;
  assign n76634 = P2_P1_DATAWIDTH_REG_0_ & n76632;
  assign n14661 = n76633 | n76634;
  assign n76636 = P2_P1_DATAWIDTH_REG_1_ & n76632;
  assign n76637 = ~n76629 & ~n76632;
  assign n14666 = n76636 | n76637;
  assign n14671 = P2_P1_DATAWIDTH_REG_2_ & n76632;
  assign n14676 = P2_P1_DATAWIDTH_REG_3_ & n76632;
  assign n14681 = P2_P1_DATAWIDTH_REG_4_ & n76632;
  assign n14686 = P2_P1_DATAWIDTH_REG_5_ & n76632;
  assign n14691 = P2_P1_DATAWIDTH_REG_6_ & n76632;
  assign n14696 = P2_P1_DATAWIDTH_REG_7_ & n76632;
  assign n14701 = P2_P1_DATAWIDTH_REG_8_ & n76632;
  assign n14706 = P2_P1_DATAWIDTH_REG_9_ & n76632;
  assign n14711 = P2_P1_DATAWIDTH_REG_10_ & n76632;
  assign n14716 = P2_P1_DATAWIDTH_REG_11_ & n76632;
  assign n14721 = P2_P1_DATAWIDTH_REG_12_ & n76632;
  assign n14726 = P2_P1_DATAWIDTH_REG_13_ & n76632;
  assign n14731 = P2_P1_DATAWIDTH_REG_14_ & n76632;
  assign n14736 = P2_P1_DATAWIDTH_REG_15_ & n76632;
  assign n14741 = P2_P1_DATAWIDTH_REG_16_ & n76632;
  assign n14746 = P2_P1_DATAWIDTH_REG_17_ & n76632;
  assign n14751 = P2_P1_DATAWIDTH_REG_18_ & n76632;
  assign n14756 = P2_P1_DATAWIDTH_REG_19_ & n76632;
  assign n14761 = P2_P1_DATAWIDTH_REG_20_ & n76632;
  assign n14766 = P2_P1_DATAWIDTH_REG_21_ & n76632;
  assign n14771 = P2_P1_DATAWIDTH_REG_22_ & n76632;
  assign n14776 = P2_P1_DATAWIDTH_REG_23_ & n76632;
  assign n14781 = P2_P1_DATAWIDTH_REG_24_ & n76632;
  assign n14786 = P2_P1_DATAWIDTH_REG_25_ & n76632;
  assign n14791 = P2_P1_DATAWIDTH_REG_26_ & n76632;
  assign n14796 = P2_P1_DATAWIDTH_REG_27_ & n76632;
  assign n14801 = P2_P1_DATAWIDTH_REG_28_ & n76632;
  assign n14806 = P2_P1_DATAWIDTH_REG_29_ & n76632;
  assign n14811 = P2_P1_DATAWIDTH_REG_30_ & n76632;
  assign n14816 = P2_P1_DATAWIDTH_REG_31_ & n76632;
  assign n76669 = P2_P1_STATE2_REG_2_ & P2_P1_STATE2_REG_1_;
  assign n76670 = P2_P1_STATE2_REG_1_ & n76584;
  assign n76671 = ~P2_P1_STATE2_REG_0_ & ~n76670;
  assign n76672 = ~P2_P1_STATEBS16_REG & ~n76584;
  assign n76673 = P2_P1_STATE_REG_2_ & ~P2_P1_STATE_REG_1_;
  assign n76674 = ~n76580 & ~n76673;
  assign n76675 = ~P2_P1_STATE_REG_0_ & ~n76674;
  assign n76676 = n76672 & n76675;
  assign n76677 = P2_P1_INSTQUEUERD_ADDR_REG_1_ & P2_P1_INSTQUEUERD_ADDR_REG_0_;
  assign n76678 = ~P2_P1_INSTQUEUERD_ADDR_REG_2_ & n76677;
  assign n76679 = P2_P1_INSTQUEUERD_ADDR_REG_3_ & n76678;
  assign n76680 = P2_P1_INSTQUEUE_REG_11__5_ & n76679;
  assign n76681 = P2_P1_INSTQUEUERD_ADDR_REG_1_ & ~P2_P1_INSTQUEUERD_ADDR_REG_0_;
  assign n76682 = ~P2_P1_INSTQUEUERD_ADDR_REG_2_ & n76681;
  assign n76683 = P2_P1_INSTQUEUERD_ADDR_REG_3_ & n76682;
  assign n76684 = P2_P1_INSTQUEUE_REG_10__5_ & n76683;
  assign n76685 = ~n76680 & ~n76684;
  assign n76686 = ~P2_P1_INSTQUEUERD_ADDR_REG_1_ & P2_P1_INSTQUEUERD_ADDR_REG_0_;
  assign n76687 = ~P2_P1_INSTQUEUERD_ADDR_REG_2_ & n76686;
  assign n76688 = P2_P1_INSTQUEUERD_ADDR_REG_3_ & n76687;
  assign n76689 = P2_P1_INSTQUEUE_REG_9__5_ & n76688;
  assign n76690 = ~P2_P1_INSTQUEUERD_ADDR_REG_1_ & ~P2_P1_INSTQUEUERD_ADDR_REG_0_;
  assign n76691 = ~P2_P1_INSTQUEUERD_ADDR_REG_2_ & n76690;
  assign n76692 = P2_P1_INSTQUEUERD_ADDR_REG_3_ & n76691;
  assign n76693 = P2_P1_INSTQUEUE_REG_8__5_ & n76692;
  assign n76694 = ~n76689 & ~n76693;
  assign n76695 = P2_P1_INSTQUEUERD_ADDR_REG_3_ & P2_P1_INSTQUEUERD_ADDR_REG_2_;
  assign n76696 = n76677 & n76695;
  assign n76697 = P2_P1_INSTQUEUE_REG_15__5_ & n76696;
  assign n76698 = n76681 & n76695;
  assign n76699 = P2_P1_INSTQUEUE_REG_14__5_ & n76698;
  assign n76700 = n76686 & n76695;
  assign n76701 = P2_P1_INSTQUEUE_REG_13__5_ & n76700;
  assign n76702 = n76690 & n76695;
  assign n76703 = P2_P1_INSTQUEUE_REG_12__5_ & n76702;
  assign n76704 = ~n76697 & ~n76699;
  assign n76705 = ~n76701 & n76704;
  assign n76706 = ~n76703 & n76705;
  assign n76707 = ~P2_P1_INSTQUEUERD_ADDR_REG_3_ & P2_P1_INSTQUEUERD_ADDR_REG_2_;
  assign n76708 = n76677 & n76707;
  assign n76709 = P2_P1_INSTQUEUE_REG_7__5_ & n76708;
  assign n76710 = n76681 & n76707;
  assign n76711 = P2_P1_INSTQUEUE_REG_6__5_ & n76710;
  assign n76712 = n76686 & n76707;
  assign n76713 = P2_P1_INSTQUEUE_REG_5__5_ & n76712;
  assign n76714 = n76690 & n76707;
  assign n76715 = P2_P1_INSTQUEUE_REG_4__5_ & n76714;
  assign n76716 = ~n76709 & ~n76711;
  assign n76717 = ~n76713 & n76716;
  assign n76718 = ~n76715 & n76717;
  assign n76719 = ~P2_P1_INSTQUEUERD_ADDR_REG_3_ & n76678;
  assign n76720 = P2_P1_INSTQUEUE_REG_3__5_ & n76719;
  assign n76721 = ~P2_P1_INSTQUEUERD_ADDR_REG_3_ & ~P2_P1_INSTQUEUERD_ADDR_REG_2_;
  assign n76722 = n76681 & n76721;
  assign n76723 = P2_P1_INSTQUEUE_REG_2__5_ & n76722;
  assign n76724 = n76686 & n76721;
  assign n76725 = P2_P1_INSTQUEUE_REG_1__5_ & n76724;
  assign n76726 = ~P2_P1_INSTQUEUERD_ADDR_REG_3_ & n76691;
  assign n76727 = P2_P1_INSTQUEUE_REG_0__5_ & n76726;
  assign n76728 = ~n76720 & ~n76723;
  assign n76729 = ~n76725 & n76728;
  assign n76730 = ~n76727 & n76729;
  assign n76731 = n76685 & n76694;
  assign n76732 = n76706 & n76731;
  assign n76733 = n76718 & n76732;
  assign n76734 = n76730 & n76733;
  assign n76735 = P2_P1_INSTQUEUE_REG_11__6_ & n76679;
  assign n76736 = P2_P1_INSTQUEUE_REG_10__6_ & n76683;
  assign n76737 = ~n76735 & ~n76736;
  assign n76738 = P2_P1_INSTQUEUE_REG_9__6_ & n76688;
  assign n76739 = P2_P1_INSTQUEUE_REG_8__6_ & n76692;
  assign n76740 = ~n76738 & ~n76739;
  assign n76741 = P2_P1_INSTQUEUE_REG_15__6_ & n76696;
  assign n76742 = P2_P1_INSTQUEUE_REG_14__6_ & n76698;
  assign n76743 = P2_P1_INSTQUEUE_REG_13__6_ & n76700;
  assign n76744 = P2_P1_INSTQUEUE_REG_12__6_ & n76702;
  assign n76745 = ~n76741 & ~n76742;
  assign n76746 = ~n76743 & n76745;
  assign n76747 = ~n76744 & n76746;
  assign n76748 = P2_P1_INSTQUEUE_REG_7__6_ & n76708;
  assign n76749 = P2_P1_INSTQUEUE_REG_6__6_ & n76710;
  assign n76750 = P2_P1_INSTQUEUE_REG_5__6_ & n76712;
  assign n76751 = P2_P1_INSTQUEUE_REG_4__6_ & n76714;
  assign n76752 = ~n76748 & ~n76749;
  assign n76753 = ~n76750 & n76752;
  assign n76754 = ~n76751 & n76753;
  assign n76755 = P2_P1_INSTQUEUE_REG_3__6_ & n76719;
  assign n76756 = P2_P1_INSTQUEUE_REG_2__6_ & n76722;
  assign n76757 = P2_P1_INSTQUEUE_REG_1__6_ & n76724;
  assign n76758 = P2_P1_INSTQUEUE_REG_0__6_ & n76726;
  assign n76759 = ~n76755 & ~n76756;
  assign n76760 = ~n76757 & n76759;
  assign n76761 = ~n76758 & n76760;
  assign n76762 = n76737 & n76740;
  assign n76763 = n76747 & n76762;
  assign n76764 = n76754 & n76763;
  assign n76765 = n76761 & n76764;
  assign n76766 = n76734 & n76765;
  assign n76767 = P2_P1_INSTQUEUE_REG_11__4_ & n76679;
  assign n76768 = P2_P1_INSTQUEUE_REG_10__4_ & n76683;
  assign n76769 = ~n76767 & ~n76768;
  assign n76770 = P2_P1_INSTQUEUE_REG_9__4_ & n76688;
  assign n76771 = P2_P1_INSTQUEUE_REG_8__4_ & n76692;
  assign n76772 = ~n76770 & ~n76771;
  assign n76773 = P2_P1_INSTQUEUE_REG_15__4_ & n76696;
  assign n76774 = P2_P1_INSTQUEUE_REG_14__4_ & n76698;
  assign n76775 = P2_P1_INSTQUEUE_REG_13__4_ & n76700;
  assign n76776 = P2_P1_INSTQUEUE_REG_12__4_ & n76702;
  assign n76777 = ~n76773 & ~n76774;
  assign n76778 = ~n76775 & n76777;
  assign n76779 = ~n76776 & n76778;
  assign n76780 = P2_P1_INSTQUEUE_REG_7__4_ & n76708;
  assign n76781 = P2_P1_INSTQUEUE_REG_6__4_ & n76710;
  assign n76782 = P2_P1_INSTQUEUE_REG_5__4_ & n76712;
  assign n76783 = P2_P1_INSTQUEUE_REG_4__4_ & n76714;
  assign n76784 = ~n76780 & ~n76781;
  assign n76785 = ~n76782 & n76784;
  assign n76786 = ~n76783 & n76785;
  assign n76787 = P2_P1_INSTQUEUE_REG_3__4_ & n76719;
  assign n76788 = P2_P1_INSTQUEUE_REG_2__4_ & n76722;
  assign n76789 = P2_P1_INSTQUEUE_REG_1__4_ & n76724;
  assign n76790 = P2_P1_INSTQUEUE_REG_0__4_ & n76726;
  assign n76791 = ~n76787 & ~n76788;
  assign n76792 = ~n76789 & n76791;
  assign n76793 = ~n76790 & n76792;
  assign n76794 = n76769 & n76772;
  assign n76795 = n76779 & n76794;
  assign n76796 = n76786 & n76795;
  assign n76797 = n76793 & n76796;
  assign n76798 = P2_P1_INSTQUEUE_REG_11__7_ & n76679;
  assign n76799 = P2_P1_INSTQUEUE_REG_10__7_ & n76683;
  assign n76800 = ~n76798 & ~n76799;
  assign n76801 = P2_P1_INSTQUEUE_REG_9__7_ & n76688;
  assign n76802 = P2_P1_INSTQUEUE_REG_8__7_ & n76692;
  assign n76803 = ~n76801 & ~n76802;
  assign n76804 = P2_P1_INSTQUEUE_REG_15__7_ & n76696;
  assign n76805 = P2_P1_INSTQUEUE_REG_14__7_ & n76698;
  assign n76806 = P2_P1_INSTQUEUE_REG_13__7_ & n76700;
  assign n76807 = P2_P1_INSTQUEUE_REG_12__7_ & n76702;
  assign n76808 = ~n76804 & ~n76805;
  assign n76809 = ~n76806 & n76808;
  assign n76810 = ~n76807 & n76809;
  assign n76811 = P2_P1_INSTQUEUE_REG_7__7_ & n76708;
  assign n76812 = P2_P1_INSTQUEUE_REG_6__7_ & n76710;
  assign n76813 = P2_P1_INSTQUEUE_REG_5__7_ & n76712;
  assign n76814 = P2_P1_INSTQUEUE_REG_4__7_ & n76714;
  assign n76815 = ~n76811 & ~n76812;
  assign n76816 = ~n76813 & n76815;
  assign n76817 = ~n76814 & n76816;
  assign n76818 = P2_P1_INSTQUEUE_REG_3__7_ & n76719;
  assign n76819 = P2_P1_INSTQUEUE_REG_2__7_ & n76722;
  assign n76820 = P2_P1_INSTQUEUE_REG_1__7_ & n76724;
  assign n76821 = P2_P1_INSTQUEUE_REG_0__7_ & n76726;
  assign n76822 = ~n76818 & ~n76819;
  assign n76823 = ~n76820 & n76822;
  assign n76824 = ~n76821 & n76823;
  assign n76825 = n76800 & n76803;
  assign n76826 = n76810 & n76825;
  assign n76827 = n76817 & n76826;
  assign n76828 = n76824 & n76827;
  assign n76829 = P2_P1_INSTQUEUE_REG_11__3_ & n76679;
  assign n76830 = P2_P1_INSTQUEUE_REG_10__3_ & n76683;
  assign n76831 = ~n76829 & ~n76830;
  assign n76832 = P2_P1_INSTQUEUE_REG_9__3_ & n76688;
  assign n76833 = P2_P1_INSTQUEUE_REG_8__3_ & n76692;
  assign n76834 = ~n76832 & ~n76833;
  assign n76835 = P2_P1_INSTQUEUE_REG_15__3_ & n76696;
  assign n76836 = P2_P1_INSTQUEUE_REG_14__3_ & n76698;
  assign n76837 = P2_P1_INSTQUEUE_REG_13__3_ & n76700;
  assign n76838 = P2_P1_INSTQUEUE_REG_12__3_ & n76702;
  assign n76839 = ~n76835 & ~n76836;
  assign n76840 = ~n76837 & n76839;
  assign n76841 = ~n76838 & n76840;
  assign n76842 = P2_P1_INSTQUEUE_REG_7__3_ & n76708;
  assign n76843 = P2_P1_INSTQUEUE_REG_6__3_ & n76710;
  assign n76844 = P2_P1_INSTQUEUE_REG_5__3_ & n76712;
  assign n76845 = P2_P1_INSTQUEUE_REG_4__3_ & n76714;
  assign n76846 = ~n76842 & ~n76843;
  assign n76847 = ~n76844 & n76846;
  assign n76848 = ~n76845 & n76847;
  assign n76849 = P2_P1_INSTQUEUE_REG_3__3_ & n76719;
  assign n76850 = P2_P1_INSTQUEUE_REG_2__3_ & n76722;
  assign n76851 = P2_P1_INSTQUEUE_REG_1__3_ & n76724;
  assign n76852 = P2_P1_INSTQUEUE_REG_0__3_ & n76726;
  assign n76853 = ~n76849 & ~n76850;
  assign n76854 = ~n76851 & n76853;
  assign n76855 = ~n76852 & n76854;
  assign n76856 = n76831 & n76834;
  assign n76857 = n76841 & n76856;
  assign n76858 = n76848 & n76857;
  assign n76859 = n76855 & n76858;
  assign n76860 = P2_P1_INSTQUEUE_REG_11__2_ & n76679;
  assign n76861 = P2_P1_INSTQUEUE_REG_10__2_ & n76683;
  assign n76862 = ~n76860 & ~n76861;
  assign n76863 = P2_P1_INSTQUEUE_REG_9__2_ & n76688;
  assign n76864 = P2_P1_INSTQUEUE_REG_8__2_ & n76692;
  assign n76865 = ~n76863 & ~n76864;
  assign n76866 = P2_P1_INSTQUEUE_REG_15__2_ & n76696;
  assign n76867 = P2_P1_INSTQUEUE_REG_14__2_ & n76698;
  assign n76868 = P2_P1_INSTQUEUE_REG_13__2_ & n76700;
  assign n76869 = P2_P1_INSTQUEUE_REG_12__2_ & n76702;
  assign n76870 = ~n76866 & ~n76867;
  assign n76871 = ~n76868 & n76870;
  assign n76872 = ~n76869 & n76871;
  assign n76873 = P2_P1_INSTQUEUE_REG_7__2_ & n76708;
  assign n76874 = P2_P1_INSTQUEUE_REG_6__2_ & n76710;
  assign n76875 = P2_P1_INSTQUEUE_REG_5__2_ & n76712;
  assign n76876 = P2_P1_INSTQUEUE_REG_4__2_ & n76714;
  assign n76877 = ~n76873 & ~n76874;
  assign n76878 = ~n76875 & n76877;
  assign n76879 = ~n76876 & n76878;
  assign n76880 = P2_P1_INSTQUEUE_REG_3__2_ & n76719;
  assign n76881 = P2_P1_INSTQUEUE_REG_2__2_ & n76722;
  assign n76882 = P2_P1_INSTQUEUE_REG_1__2_ & n76724;
  assign n76883 = P2_P1_INSTQUEUE_REG_0__2_ & n76726;
  assign n76884 = ~n76880 & ~n76881;
  assign n76885 = ~n76882 & n76884;
  assign n76886 = ~n76883 & n76885;
  assign n76887 = n76862 & n76865;
  assign n76888 = n76872 & n76887;
  assign n76889 = n76879 & n76888;
  assign n76890 = n76886 & n76889;
  assign n76891 = ~n76828 & ~n76859;
  assign n76892 = n76890 & n76891;
  assign n76893 = n76766 & n76797;
  assign n76894 = n76892 & n76893;
  assign n76895 = P2_P1_INSTQUEUE_REG_11__1_ & n76679;
  assign n76896 = P2_P1_INSTQUEUE_REG_10__1_ & n76683;
  assign n76897 = ~n76895 & ~n76896;
  assign n76898 = P2_P1_INSTQUEUE_REG_9__1_ & n76688;
  assign n76899 = P2_P1_INSTQUEUE_REG_8__1_ & n76692;
  assign n76900 = ~n76898 & ~n76899;
  assign n76901 = P2_P1_INSTQUEUE_REG_15__1_ & n76696;
  assign n76902 = P2_P1_INSTQUEUE_REG_14__1_ & n76698;
  assign n76903 = P2_P1_INSTQUEUE_REG_13__1_ & n76700;
  assign n76904 = P2_P1_INSTQUEUE_REG_12__1_ & n76702;
  assign n76905 = ~n76901 & ~n76902;
  assign n76906 = ~n76903 & n76905;
  assign n76907 = ~n76904 & n76906;
  assign n76908 = P2_P1_INSTQUEUE_REG_7__1_ & n76708;
  assign n76909 = P2_P1_INSTQUEUE_REG_6__1_ & n76710;
  assign n76910 = P2_P1_INSTQUEUE_REG_5__1_ & n76712;
  assign n76911 = P2_P1_INSTQUEUE_REG_4__1_ & n76714;
  assign n76912 = ~n76908 & ~n76909;
  assign n76913 = ~n76910 & n76912;
  assign n76914 = ~n76911 & n76913;
  assign n76915 = P2_P1_INSTQUEUE_REG_3__1_ & n76719;
  assign n76916 = P2_P1_INSTQUEUE_REG_2__1_ & n76722;
  assign n76917 = P2_P1_INSTQUEUE_REG_1__1_ & n76724;
  assign n76918 = P2_P1_INSTQUEUE_REG_0__1_ & n76726;
  assign n76919 = ~n76915 & ~n76916;
  assign n76920 = ~n76917 & n76919;
  assign n76921 = ~n76918 & n76920;
  assign n76922 = n76897 & n76900;
  assign n76923 = n76907 & n76922;
  assign n76924 = n76914 & n76923;
  assign n76925 = n76921 & n76924;
  assign n76926 = P2_P1_INSTQUEUE_REG_11__0_ & n76679;
  assign n76927 = P2_P1_INSTQUEUE_REG_10__0_ & n76683;
  assign n76928 = ~n76926 & ~n76927;
  assign n76929 = P2_P1_INSTQUEUE_REG_9__0_ & n76688;
  assign n76930 = P2_P1_INSTQUEUE_REG_8__0_ & n76692;
  assign n76931 = ~n76929 & ~n76930;
  assign n76932 = P2_P1_INSTQUEUE_REG_15__0_ & n76696;
  assign n76933 = P2_P1_INSTQUEUE_REG_14__0_ & n76698;
  assign n76934 = P2_P1_INSTQUEUE_REG_13__0_ & n76700;
  assign n76935 = P2_P1_INSTQUEUE_REG_12__0_ & n76702;
  assign n76936 = ~n76932 & ~n76933;
  assign n76937 = ~n76934 & n76936;
  assign n76938 = ~n76935 & n76937;
  assign n76939 = P2_P1_INSTQUEUE_REG_7__0_ & n76708;
  assign n76940 = P2_P1_INSTQUEUE_REG_6__0_ & n76710;
  assign n76941 = P2_P1_INSTQUEUE_REG_5__0_ & n76712;
  assign n76942 = P2_P1_INSTQUEUE_REG_4__0_ & n76714;
  assign n76943 = ~n76939 & ~n76940;
  assign n76944 = ~n76941 & n76943;
  assign n76945 = ~n76942 & n76944;
  assign n76946 = P2_P1_INSTQUEUE_REG_3__0_ & n76719;
  assign n76947 = P2_P1_INSTQUEUE_REG_2__0_ & n76722;
  assign n76948 = P2_P1_INSTQUEUE_REG_1__0_ & n76724;
  assign n76949 = P2_P1_INSTQUEUE_REG_0__0_ & n76726;
  assign n76950 = ~n76946 & ~n76947;
  assign n76951 = ~n76948 & n76950;
  assign n76952 = ~n76949 & n76951;
  assign n76953 = n76928 & n76931;
  assign n76954 = n76938 & n76953;
  assign n76955 = n76945 & n76954;
  assign n76956 = n76952 & n76955;
  assign n76957 = n76925 & ~n76956;
  assign n76958 = n76894 & n76957;
  assign n76959 = n76676 & n76958;
  assign n76960 = ~P2_P1_STATE2_REG_1_ & ~n76959;
  assign n76961 = ~n76584 & n76675;
  assign n76962 = ~n76890 & ~n76925;
  assign n76963 = n76961 & n76962;
  assign n76964 = ~n76584 & ~n76890;
  assign n76965 = n76925 & n76964;
  assign n76966 = ~n76584 & n76890;
  assign n76967 = n76925 & ~n76961;
  assign n76968 = n76966 & ~n76967;
  assign n76969 = ~n76963 & ~n76965;
  assign n76970 = ~n76968 & n76969;
  assign n76971 = P2_P1_INSTQUEUERD_ADDR_REG_4_ & ~P2_P1_INSTQUEUEWR_ADDR_REG_4_;
  assign n76972 = ~P2_P1_INSTQUEUERD_ADDR_REG_3_ & P2_P1_INSTQUEUEWR_ADDR_REG_3_;
  assign n76973 = P2_P1_INSTQUEUERD_ADDR_REG_3_ & ~P2_P1_INSTQUEUEWR_ADDR_REG_3_;
  assign n76974 = ~P2_P1_INSTQUEUERD_ADDR_REG_2_ & P2_P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n76975 = P2_P1_INSTQUEUERD_ADDR_REG_2_ & ~P2_P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n76976 = P2_P1_INSTQUEUERD_ADDR_REG_0_ & ~P2_P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n76977 = P2_P1_INSTQUEUEWR_ADDR_REG_1_ & ~n76976;
  assign n76978 = ~P2_P1_INSTQUEUEWR_ADDR_REG_1_ & n76976;
  assign n76979 = ~P2_P1_INSTQUEUERD_ADDR_REG_1_ & ~n76978;
  assign n76980 = ~n76977 & ~n76979;
  assign n76981 = ~n76975 & ~n76980;
  assign n76982 = ~n76974 & ~n76981;
  assign n76983 = ~n76973 & ~n76982;
  assign n76984 = ~n76972 & ~n76983;
  assign n76985 = ~P2_P1_INSTQUEUERD_ADDR_REG_4_ & P2_P1_INSTQUEUEWR_ADDR_REG_4_;
  assign n76986 = n76984 & ~n76985;
  assign n76987 = ~n76971 & ~n76986;
  assign n76988 = ~n76971 & ~n76985;
  assign n76989 = ~n76984 & ~n76988;
  assign n76990 = n76984 & n76988;
  assign n76991 = ~n76989 & ~n76990;
  assign n76992 = ~n76972 & ~n76973;
  assign n76993 = ~n76982 & ~n76992;
  assign n76994 = n76982 & n76992;
  assign n76995 = ~n76993 & ~n76994;
  assign n76996 = ~P2_P1_INSTQUEUERD_ADDR_REG_1_ & P2_P1_INSTQUEUEWR_ADDR_REG_1_;
  assign n76997 = P2_P1_INSTQUEUERD_ADDR_REG_1_ & ~P2_P1_INSTQUEUEWR_ADDR_REG_1_;
  assign n76998 = ~n76996 & ~n76997;
  assign n76999 = ~n76976 & ~n76998;
  assign n77000 = n76976 & n76998;
  assign n77001 = ~n76999 & ~n77000;
  assign n77002 = ~n76974 & ~n76975;
  assign n77003 = ~n76980 & ~n77002;
  assign n77004 = n76980 & n77002;
  assign n77005 = ~n77003 & ~n77004;
  assign n77006 = n76991 & n76995;
  assign n77007 = n77001 & n77006;
  assign n77008 = n77005 & n77007;
  assign n77009 = n76987 & ~n77008;
  assign n77010 = ~n76925 & ~n77009;
  assign n77011 = n76925 & ~n77009;
  assign n77012 = ~n77010 & ~n77011;
  assign n77013 = ~n76828 & n76859;
  assign n77014 = ~n76734 & ~n76765;
  assign n77015 = n76797 & n77014;
  assign n77016 = n77013 & n77015;
  assign n77017 = n76956 & n77016;
  assign n77018 = n77012 & n77017;
  assign n77019 = ~n76890 & ~n77018;
  assign n77020 = ~n76859 & ~n76956;
  assign n77021 = ~n76828 & n77020;
  assign n77022 = n76893 & n77021;
  assign n77023 = ~n77010 & n77022;
  assign n77024 = ~n77011 & n77023;
  assign n77025 = n76890 & ~n77024;
  assign n77026 = ~n77019 & ~n77025;
  assign n77027 = n76970 & n77026;
  assign n77028 = ~P2_P1_FLUSH_REG & ~P2_P1_MORE_REG;
  assign n77029 = n77027 & ~n77028;
  assign n77030 = ~n76925 & n76956;
  assign n77031 = ~n76890 & n77030;
  assign n77032 = n77016 & n77031;
  assign n77033 = ~n77009 & n77032;
  assign n77034 = n76925 & n76956;
  assign n77035 = ~n76890 & n77034;
  assign n77036 = n77016 & n77035;
  assign n77037 = ~n77009 & n77036;
  assign n77038 = n76958 & ~n77009;
  assign n77039 = ~n76925 & ~n76956;
  assign n77040 = n76894 & n77039;
  assign n77041 = ~n77009 & n77040;
  assign n77042 = ~n77033 & ~n77037;
  assign n77043 = ~n77038 & n77042;
  assign n77044 = ~n77041 & n77043;
  assign n77045 = ~n76734 & n76765;
  assign n77046 = ~n76797 & n77045;
  assign n77047 = n76892 & n77046;
  assign n77048 = n77039 & n77047;
  assign n77049 = ~P2_P1_INSTQUEUERD_ADDR_REG_0_ & P2_P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n77050 = ~n76976 & ~n77049;
  assign n77051 = n77001 & n77050;
  assign n77052 = ~n77005 & ~n77051;
  assign n77053 = n77006 & ~n77052;
  assign n77054 = n76987 & ~n77053;
  assign n77055 = n77048 & ~n77054;
  assign n77056 = n77034 & n77047;
  assign n77057 = ~n77054 & n77056;
  assign n77058 = n76892 & n77015;
  assign n77059 = n76957 & n77058;
  assign n77060 = n76991 & ~n77052;
  assign n77061 = n76995 & n77060;
  assign n77062 = n76987 & ~n77061;
  assign n77063 = n77059 & ~n77062;
  assign n77064 = n77039 & n77058;
  assign n77065 = ~n77001 & ~n77050;
  assign n77066 = n77006 & ~n77065;
  assign n77067 = n77005 & n77066;
  assign n77068 = n76987 & ~n77067;
  assign n77069 = n77064 & ~n77068;
  assign n77070 = ~n77055 & ~n77057;
  assign n77071 = ~n77063 & n77070;
  assign n77072 = ~n77069 & n77071;
  assign n77073 = n77044 & n77072;
  assign n77074 = ~n77027 & ~n77073;
  assign n77075 = ~n76925 & ~n77068;
  assign n77076 = n76925 & ~n77062;
  assign n77077 = ~n77075 & ~n77076;
  assign n77078 = ~n76956 & n77058;
  assign n77079 = n77077 & n77078;
  assign n77080 = n76859 & n76890;
  assign n77081 = n76734 & ~n76765;
  assign n77082 = n77080 & n77081;
  assign n77083 = n77034 & n77082;
  assign n77084 = ~n76828 & n77083;
  assign n77085 = n76894 & ~n76956;
  assign n77086 = ~n77032 & ~n77084;
  assign n77087 = ~n77085 & n77086;
  assign n77088 = n76765 & n76859;
  assign n77089 = ~n76797 & n76890;
  assign n77090 = ~n76828 & n77034;
  assign n77091 = n77089 & n77090;
  assign n77092 = n76734 & ~n76890;
  assign n77093 = n76797 & n76828;
  assign n77094 = n77092 & n77093;
  assign n77095 = ~n77091 & ~n77094;
  assign n77096 = n77088 & ~n77095;
  assign n77097 = n77039 & n77093;
  assign n77098 = n77082 & n77097;
  assign n77099 = n76859 & ~n76890;
  assign n77100 = n76828 & n77030;
  assign n77101 = n77015 & n77099;
  assign n77102 = n77100 & n77101;
  assign n77103 = ~n76925 & n77058;
  assign n77104 = ~n77102 & ~n77103;
  assign n77105 = ~n77096 & ~n77098;
  assign n77106 = n77104 & n77105;
  assign n77107 = n76765 & ~n76828;
  assign n77108 = ~n77081 & ~n77107;
  assign n77109 = n76859 & n77108;
  assign n77110 = ~n76890 & ~n77109;
  assign n77111 = ~n76828 & ~n77081;
  assign n77112 = ~n77045 & n77111;
  assign n77113 = ~n76859 & n77112;
  assign n77114 = n76957 & ~n77113;
  assign n77115 = n77014 & n77034;
  assign n77116 = n76734 & n76828;
  assign n77117 = ~n76891 & ~n77116;
  assign n77118 = ~n76925 & n77117;
  assign n77119 = n76765 & n76797;
  assign n77120 = n76956 & n77119;
  assign n77121 = ~n77115 & ~n77118;
  assign n77122 = ~n77120 & n77121;
  assign n77123 = ~n77114 & n77122;
  assign n77124 = n76890 & ~n77123;
  assign n77125 = ~n76859 & ~n77119;
  assign n77126 = n76734 & n77125;
  assign n77127 = n76828 & n76925;
  assign n77128 = n76956 & ~n77127;
  assign n77129 = n76859 & ~n77128;
  assign n77130 = ~n76734 & n77129;
  assign n77131 = ~n76828 & ~n77014;
  assign n77132 = ~n76957 & n77131;
  assign n77133 = ~n76797 & ~n77132;
  assign n77134 = n76765 & ~n76925;
  assign n77135 = n76828 & n77134;
  assign n77136 = n76797 & ~n76925;
  assign n77137 = n77045 & n77136;
  assign n77138 = ~n77014 & n77030;
  assign n77139 = ~n77135 & ~n77137;
  assign n77140 = ~n77138 & n77139;
  assign n77141 = ~n77126 & ~n77130;
  assign n77142 = ~n77133 & n77141;
  assign n77143 = n77140 & n77142;
  assign n77144 = ~n77110 & ~n77124;
  assign n77145 = n77143 & n77144;
  assign n77146 = n77106 & n77145;
  assign n77147 = ~n77083 & n77146;
  assign n77148 = P2_P1_INSTQUEUERD_ADDR_REG_0_ & ~n77147;
  assign n77149 = n77087 & ~n77148;
  assign n77150 = ~P2_P1_INSTQUEUERD_ADDR_REG_2_ & ~n77149;
  assign n77151 = P2_P1_INSTQUEUERD_ADDR_REG_1_ & n77150;
  assign n77152 = P2_P1_INSTQUEUERD_ADDR_REG_2_ & ~n77087;
  assign n77153 = ~P2_P1_INSTQUEUERD_ADDR_REG_1_ & n77152;
  assign n77154 = ~P2_P1_INSTQUEUERD_ADDR_REG_2_ & P2_P1_INSTQUEUERD_ADDR_REG_1_;
  assign n77155 = P2_P1_INSTQUEUERD_ADDR_REG_2_ & ~P2_P1_INSTQUEUERD_ADDR_REG_1_;
  assign n77156 = ~n77154 & ~n77155;
  assign n77157 = n77036 & ~n77156;
  assign n77158 = P2_P1_INSTQUEUERD_ADDR_REG_2_ & ~n76677;
  assign n77159 = ~n76678 & ~n77158;
  assign n77160 = ~n77034 & ~n77039;
  assign n77161 = n77159 & ~n77160;
  assign n77162 = n77047 & n77161;
  assign n77163 = ~n77157 & ~n77162;
  assign n77164 = n76925 & n77088;
  assign n77165 = ~n77089 & ~n77094;
  assign n77166 = n77164 & ~n77165;
  assign n77167 = n77093 & ~n77160;
  assign n77168 = n77082 & n77167;
  assign n77169 = ~n77166 & ~n77168;
  assign n77170 = n77104 & n77169;
  assign n77171 = n77145 & n77170;
  assign n77172 = n77158 & ~n77171;
  assign n77173 = n77163 & ~n77172;
  assign n77174 = ~n77151 & ~n77153;
  assign n77175 = n77173 & n77174;
  assign n77176 = n76797 & n76956;
  assign n77177 = ~n76859 & ~n77030;
  assign n77178 = n77111 & ~n77176;
  assign n77179 = n77177 & n77178;
  assign n77180 = ~n77137 & n77179;
  assign n77181 = n76890 & ~n77180;
  assign n77182 = ~n76890 & ~n77017;
  assign n77183 = n76957 & ~n77112;
  assign n77184 = ~n77181 & ~n77182;
  assign n77185 = ~n77183 & n77184;
  assign n77186 = n77054 & n77056;
  assign n77187 = n77009 & n77036;
  assign n77188 = n77009 & n77040;
  assign n77189 = ~n77187 & ~n77188;
  assign n77190 = ~n76584 & ~n77189;
  assign n77191 = ~n77186 & ~n77190;
  assign n77192 = n77048 & n77054;
  assign n77193 = ~n77045 & n77089;
  assign n77194 = ~n77192 & ~n77193;
  assign n77195 = n77009 & n77032;
  assign n77196 = n76958 & n77009;
  assign n77197 = ~n77195 & ~n77196;
  assign n77198 = n76961 & ~n77197;
  assign n77199 = n77194 & ~n77198;
  assign n77200 = n77185 & n77191;
  assign n77201 = n77199 & n77200;
  assign n77202 = ~n77175 & ~n77201;
  assign n77203 = P2_P1_INSTQUEUERD_ADDR_REG_2_ & n77201;
  assign n77204 = ~n77202 & ~n77203;
  assign n77205 = P2_P1_INSTQUEUERD_ADDR_REG_1_ & n76707;
  assign n77206 = ~n77149 & n77205;
  assign n77207 = P2_P1_INSTQUEUERD_ADDR_REG_2_ & n76677;
  assign n77208 = P2_P1_INSTQUEUERD_ADDR_REG_3_ & ~n77207;
  assign n77209 = ~n77170 & n77208;
  assign n77210 = P2_P1_INSTQUEUERD_ADDR_REG_2_ & P2_P1_INSTQUEUERD_ADDR_REG_1_;
  assign n77211 = ~P2_P1_INSTQUEUERD_ADDR_REG_3_ & n77210;
  assign n77212 = P2_P1_INSTQUEUERD_ADDR_REG_3_ & ~n77210;
  assign n77213 = ~n77211 & ~n77212;
  assign n77214 = n77036 & ~n77213;
  assign n77215 = ~n77209 & ~n77214;
  assign n77216 = ~n76797 & n77084;
  assign n77217 = n76797 & n77084;
  assign n77218 = ~n76958 & ~n77040;
  assign n77219 = ~n77032 & n77218;
  assign n77220 = ~n77216 & ~n77217;
  assign n77221 = n77219 & n77220;
  assign n77222 = n77145 & n77221;
  assign n77223 = n77212 & ~n77222;
  assign n77224 = P2_P1_INSTQUEUERD_ADDR_REG_3_ & ~P2_P1_INSTQUEUERD_ADDR_REG_0_;
  assign n77225 = ~n77145 & n77224;
  assign n77226 = ~n76677 & n76721;
  assign n77227 = ~P2_P1_INSTQUEUERD_ADDR_REG_2_ & ~n76677;
  assign n77228 = P2_P1_INSTQUEUERD_ADDR_REG_3_ & ~n77227;
  assign n77229 = ~n77226 & ~n77228;
  assign n77230 = ~n77160 & n77229;
  assign n77231 = n77047 & n77230;
  assign n77232 = ~n77225 & ~n77231;
  assign n77233 = n77215 & ~n77223;
  assign n77234 = n77232 & n77233;
  assign n77235 = ~n77206 & n77234;
  assign n77236 = ~n77201 & ~n77235;
  assign n77237 = P2_P1_INSTQUEUERD_ADDR_REG_3_ & n77201;
  assign n77238 = ~n77236 & ~n77237;
  assign n77239 = ~n77204 & ~n77238;
  assign n77240 = P2_P1_INSTQUEUERD_ADDR_REG_4_ & n77201;
  assign n77241 = P2_P1_INSTQUEUERD_ADDR_REG_3_ & n77210;
  assign n77242 = ~P2_P1_INSTQUEUERD_ADDR_REG_4_ & n77241;
  assign n77243 = P2_P1_INSTQUEUERD_ADDR_REG_4_ & ~n77241;
  assign n77244 = ~n77242 & ~n77243;
  assign n77245 = n77036 & ~n77244;
  assign n77246 = ~n77201 & n77245;
  assign n77247 = ~n77240 & ~n77246;
  assign n77248 = ~n77239 & n77247;
  assign n77249 = ~P2_P1_INSTQUEUEWR_ADDR_REG_3_ & ~n77238;
  assign n77250 = ~P2_P1_INSTQUEUEWR_ADDR_REG_4_ & ~n77247;
  assign n77251 = P2_P1_INSTQUEUEWR_ADDR_REG_2_ & n77204;
  assign n77252 = P2_P1_INSTQUEUEWR_ADDR_REG_3_ & n77238;
  assign n77253 = n77045 & n77091;
  assign n77254 = ~n77048 & ~n77253;
  assign n77255 = n77083 & n77093;
  assign n77256 = n77146 & ~n77255;
  assign n77257 = n77254 & n77256;
  assign n77258 = ~P2_P1_INSTQUEUERD_ADDR_REG_0_ & ~n77257;
  assign n77259 = P2_P1_INSTQUEUERD_ADDR_REG_0_ & ~n77087;
  assign n77260 = P2_P1_INSTQUEUERD_ADDR_REG_0_ & n77036;
  assign n77261 = ~n77258 & ~n77259;
  assign n77262 = ~n77260 & n77261;
  assign n77263 = ~n77201 & ~n77262;
  assign n77264 = P2_P1_INSTQUEUERD_ADDR_REG_0_ & n77201;
  assign n77265 = ~n77263 & ~n77264;
  assign n77266 = P2_P1_INSTQUEUEWR_ADDR_REG_0_ & n77265;
  assign n77267 = ~P2_P1_INSTQUEUEWR_ADDR_REG_1_ & ~n77266;
  assign n77268 = ~P2_P1_INSTQUEUEWR_ADDR_REG_2_ & ~n77204;
  assign n77269 = ~P2_P1_INSTQUEUERD_ADDR_REG_1_ & ~n77149;
  assign n77270 = ~P2_P1_INSTQUEUERD_ADDR_REG_1_ & n77036;
  assign n77271 = ~n76677 & ~n76690;
  assign n77272 = ~n77254 & n77271;
  assign n77273 = ~n77270 & ~n77272;
  assign n77274 = n76681 & ~n77256;
  assign n77275 = n77273 & ~n77274;
  assign n77276 = ~n77269 & n77275;
  assign n77277 = ~n77201 & ~n77276;
  assign n77278 = P2_P1_INSTQUEUERD_ADDR_REG_1_ & n77201;
  assign n77279 = ~n77277 & ~n77278;
  assign n77280 = P2_P1_INSTQUEUEWR_ADDR_REG_1_ & n77266;
  assign n77281 = ~n77279 & ~n77280;
  assign n77282 = ~n77267 & ~n77268;
  assign n77283 = ~n77281 & n77282;
  assign n77284 = ~n77251 & ~n77252;
  assign n77285 = ~n77283 & n77284;
  assign n77286 = ~n77249 & ~n77250;
  assign n77287 = ~n77285 & n77286;
  assign n77288 = P2_P1_INSTQUEUEWR_ADDR_REG_4_ & n77247;
  assign n77289 = ~n77287 & ~n77288;
  assign n77290 = ~n77029 & ~n77074;
  assign n77291 = ~n77079 & n77290;
  assign n77292 = n77248 & n77291;
  assign n77293 = ~n77289 & n77292;
  assign n77294 = n76960 & n77293;
  assign n77295 = P2_P1_STATE2_REG_0_ & ~n77294;
  assign n77296 = ~n76671 & ~n77295;
  assign n77297 = P2_P1_STATE2_REG_2_ & n77296;
  assign n77298 = P2_P1_STATE2_REG_0_ & ~n77297;
  assign n77299 = n76669 & n77298;
  assign n77300 = P2_P1_STATE2_REG_3_ & ~n77298;
  assign n14821 = n77299 | n77300;
  assign n77302 = ~P2_P1_STATE2_REG_2_ & ~n76584;
  assign n77303 = P2_P1_STATE2_REG_0_ & ~n77302;
  assign n77304 = ~P2_P1_STATE2_REG_0_ & ~P2_P1_STATEBS16_REG;
  assign n77305 = ~n77303 & ~n77304;
  assign n77306 = P2_P1_STATE2_REG_1_ & n77305;
  assign n77307 = P2_P1_STATE2_REG_2_ & ~P2_P1_STATE2_REG_1_;
  assign n77308 = ~n77306 & ~n77307;
  assign n77309 = P2_P1_STATE2_REG_2_ & ~n77298;
  assign n14826 = ~n77308 | n77309;
  assign n77311 = P2_P1_STATE2_REG_0_ & n77307;
  assign n77312 = ~n77297 & n77311;
  assign n77313 = ~P2_P1_STATE2_REG_2_ & P2_P1_STATE2_REG_0_;
  assign n77314 = n76584 & n77313;
  assign n77315 = ~n77297 & ~n77314;
  assign n77316 = P2_P1_STATE2_REG_1_ & ~n77315;
  assign n77317 = ~P2_P1_STATE2_REG_3_ & ~P2_P1_STATE2_REG_1_;
  assign n77318 = ~n76584 & n77317;
  assign n77319 = n77298 & n77318;
  assign n77320 = P2_P1_STATE2_REG_1_ & ~P2_P1_STATE2_REG_0_;
  assign n77321 = ~P2_P1_STATE2_REG_2_ & n77320;
  assign n77322 = ~P2_P1_STATEBS16_REG & n77321;
  assign n77323 = ~n77312 & ~n77316;
  assign n77324 = ~n77319 & n77323;
  assign n14831 = n77322 | ~n77324;
  assign n77326 = P2_P1_STATE2_REG_3_ & ~P2_P1_INSTQUEUERD_ADDR_REG_4_;
  assign n77327 = ~P2_P1_STATE2_REG_2_ & ~P2_P1_STATE2_REG_1_;
  assign n77328 = n77326 & n77327;
  assign n77329 = ~n77297 & ~n77328;
  assign n77330 = ~P2_P1_STATE2_REG_0_ & n77329;
  assign n77331 = P2_P1_INSTADDRPOINTER_REG_0_ & P2_P1_INSTADDRPOINTER_REG_31_;
  assign n77332 = P2_P1_INSTADDRPOINTER_REG_0_ & ~P2_P1_INSTADDRPOINTER_REG_31_;
  assign n77333 = ~n77331 & ~n77332;
  assign n77334 = P2_P1_FLUSH_REG & n77333;
  assign n77335 = P2_P1_INSTQUEUERD_ADDR_REG_0_ & ~P2_P1_FLUSH_REG;
  assign n77336 = ~n77334 & ~n77335;
  assign n77337 = P2_P1_INSTADDRPOINTER_REG_0_ & ~P2_P1_INSTADDRPOINTER_REG_1_;
  assign n77338 = ~P2_P1_INSTADDRPOINTER_REG_0_ & P2_P1_INSTADDRPOINTER_REG_1_;
  assign n77339 = ~n77337 & ~n77338;
  assign n77340 = P2_P1_INSTADDRPOINTER_REG_31_ & ~n77339;
  assign n77341 = P2_P1_INSTADDRPOINTER_REG_1_ & ~P2_P1_INSTADDRPOINTER_REG_31_;
  assign n77342 = ~n77340 & ~n77341;
  assign n77343 = ~n77333 & n77342;
  assign n77344 = P2_P1_FLUSH_REG & n77343;
  assign n77345 = P2_P1_INSTQUEUERD_ADDR_REG_1_ & ~P2_P1_FLUSH_REG;
  assign n77346 = ~n77344 & ~n77345;
  assign n77347 = n77336 & n77346;
  assign n77348 = P2_P1_INSTQUEUERD_ADDR_REG_3_ & ~P2_P1_FLUSH_REG;
  assign n77349 = ~n77333 & ~n77342;
  assign n77350 = P2_P1_FLUSH_REG & n77349;
  assign n77351 = P2_P1_INSTQUEUERD_ADDR_REG_2_ & ~P2_P1_FLUSH_REG;
  assign n77352 = ~n77350 & ~n77351;
  assign n77353 = ~n77347 & n77348;
  assign n77354 = ~n77352 & n77353;
  assign n77355 = P2_P1_INSTQUEUERD_ADDR_REG_4_ & ~P2_P1_FLUSH_REG;
  assign n77356 = ~n77354 & ~n77355;
  assign n77357 = n76669 & n77356;
  assign n77358 = ~n77297 & ~n77357;
  assign n77359 = P2_P1_STATE2_REG_0_ & ~n77358;
  assign n77360 = P2_P1_STATE2_REG_3_ & P2_P1_STATE2_REG_0_;
  assign n77361 = n77327 & n77360;
  assign n77362 = ~n77314 & ~n77361;
  assign n77363 = ~n77293 & n77311;
  assign n77364 = n77362 & ~n77363;
  assign n77365 = ~n77330 & ~n77359;
  assign n14836 = ~n77364 | ~n77365;
  assign n77367 = P2_P1_INSTQUEUEWR_ADDR_REG_1_ & P2_P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n77368 = P2_P1_INSTQUEUEWR_ADDR_REG_2_ & n77367;
  assign n77369 = P2_P1_INSTQUEUEWR_ADDR_REG_3_ & n77368;
  assign n77370 = P2_P1_STATE2_REG_3_ & ~n77369;
  assign n77371 = ~P2_P1_STATE2_REG_2_ & P2_P1_STATE2_REG_1_;
  assign n77372 = ~n77307 & ~n77371;
  assign n77373 = ~n77326 & n77372;
  assign n77374 = ~P2_P1_STATE2_REG_0_ & ~n77373;
  assign n77375 = ~n77370 & n77374;
  assign n77376 = ~P2_P1_INSTQUEUEWR_ADDR_REG_2_ & n77367;
  assign n77377 = P2_P1_INSTQUEUEWR_ADDR_REG_2_ & ~n77367;
  assign n77378 = ~n77376 & ~n77377;
  assign n77379 = ~P2_P1_INSTQUEUEWR_ADDR_REG_3_ & n77368;
  assign n77380 = P2_P1_INSTQUEUEWR_ADDR_REG_3_ & ~n77368;
  assign n77381 = ~n77379 & ~n77380;
  assign n77382 = ~n77378 & ~n77381;
  assign n77383 = ~P2_P1_INSTQUEUEWR_ADDR_REG_1_ & P2_P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n77384 = P2_P1_INSTQUEUEWR_ADDR_REG_1_ & ~P2_P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n77385 = ~n77383 & ~n77384;
  assign n77386 = ~P2_P1_INSTQUEUEWR_ADDR_REG_0_ & ~n77385;
  assign n77387 = n77382 & n77386;
  assign n77388 = ~n77369 & ~n77387;
  assign n77389 = ~P2_P1_STATE2_REG_3_ & ~P2_P1_STATE2_REG_2_;
  assign n77390 = ~P2_P1_STATEBS16_REG & n77389;
  assign n77391 = ~P2_P1_STATE2_REG_2_ & ~n77390;
  assign n77392 = P2_P1_INSTQUEUEWR_ADDR_REG_0_ & ~n77385;
  assign n77393 = ~P2_P1_INSTQUEUEWR_ADDR_REG_0_ & n77385;
  assign n77394 = ~n77392 & ~n77393;
  assign n77395 = ~P2_P1_INSTQUEUEWR_ADDR_REG_0_ & ~n77394;
  assign n77396 = P2_P1_INSTQUEUEWR_ADDR_REG_0_ & n77394;
  assign n77397 = ~n77395 & ~n77396;
  assign n77398 = ~P2_P1_INSTQUEUEWR_ADDR_REG_0_ & ~n77397;
  assign n77399 = ~n77378 & ~n77386;
  assign n77400 = n77378 & n77386;
  assign n77401 = ~n77399 & ~n77400;
  assign n77402 = P2_P1_INSTQUEUEWR_ADDR_REG_0_ & ~n77394;
  assign n77403 = ~n77401 & ~n77402;
  assign n77404 = n77401 & n77402;
  assign n77405 = ~n77403 & ~n77404;
  assign n77406 = ~n77378 & n77381;
  assign n77407 = n77386 & n77406;
  assign n77408 = ~n77378 & n77386;
  assign n77409 = ~n77381 & ~n77408;
  assign n77410 = ~n77407 & ~n77409;
  assign n77411 = n77401 & ~n77410;
  assign n77412 = ~n77402 & ~n77410;
  assign n77413 = ~n77411 & ~n77412;
  assign n77414 = ~n77401 & n77410;
  assign n77415 = n77402 & n77414;
  assign n77416 = n77413 & ~n77415;
  assign n77417 = ~n77405 & ~n77416;
  assign n77418 = n77398 & n77417;
  assign n77419 = ~n77401 & ~n77410;
  assign n77420 = n77402 & n77419;
  assign n77421 = ~n77418 & ~n77420;
  assign n77422 = n77391 & ~n77421;
  assign n77423 = n77388 & ~n77422;
  assign n77424 = n77375 & ~n77423;
  assign n77425 = P2_P1_INSTQUEUE_REG_15__7_ & ~n77424;
  assign n77426 = P2_P1_STATE2_REG_3_ & n77374;
  assign n77427 = ~n76828 & n77426;
  assign n77428 = n77369 & n77427;
  assign n77429 = P2_P1_STATEBS16_REG & n77389;
  assign n77430 = n77421 & n77429;
  assign n77431 = n77391 & ~n77430;
  assign n77432 = ~n77388 & ~n77431;
  assign n77433 = P2_BUF1_REG_7_ & n12802;
  assign n77434 = ~SEL & DIN_6_;
  assign n77435 = P3_DATAO_REG_0_ & n77434;
  assign n77436 = ~SEL & DIN_5_;
  assign n77437 = P3_DATAO_REG_0_ & n77436;
  assign n77438 = ~SEL & DIN_3_;
  assign n77439 = P3_DATAO_REG_1_ & n77438;
  assign n77440 = ~SEL & DIN_2_;
  assign n77441 = P3_DATAO_REG_1_ & n77440;
  assign n77442 = ~SEL & DIN_1_;
  assign n77443 = P3_DATAO_REG_2_ & n77442;
  assign n77444 = ~SEL & DIN_0_;
  assign n77445 = P3_DATAO_REG_3_ & n77444;
  assign n77446 = n77443 & ~n77445;
  assign n77447 = ~n77443 & n77445;
  assign n77448 = ~n77446 & ~n77447;
  assign n77449 = n77441 & ~n77448;
  assign n77450 = P3_DATAO_REG_1_ & P3_DATAO_REG_2_;
  assign n77451 = n77442 & n77444;
  assign n77452 = n77450 & n77451;
  assign n77453 = ~n77441 & n77448;
  assign n77454 = n77452 & ~n77453;
  assign n77455 = ~n77449 & ~n77454;
  assign n77456 = n77439 & ~n77455;
  assign n77457 = P3_DATAO_REG_2_ & n77440;
  assign n77458 = P3_DATAO_REG_4_ & n77444;
  assign n77459 = P3_DATAO_REG_3_ & n77442;
  assign n77460 = n77458 & ~n77459;
  assign n77461 = ~n77458 & n77459;
  assign n77462 = ~n77460 & ~n77461;
  assign n77463 = n77457 & ~n77462;
  assign n77464 = ~n77457 & n77462;
  assign n77465 = P3_DATAO_REG_2_ & P3_DATAO_REG_3_;
  assign n77466 = n77451 & n77465;
  assign n77467 = ~n77463 & ~n77464;
  assign n77468 = ~n77466 & n77467;
  assign n77469 = n77466 & ~n77467;
  assign n77470 = ~n77468 & ~n77469;
  assign n77471 = n77439 & ~n77470;
  assign n77472 = ~n77455 & ~n77470;
  assign n77473 = ~n77456 & ~n77471;
  assign n77474 = ~n77472 & n77473;
  assign n77475 = ~SEL & DIN_4_;
  assign n77476 = P3_DATAO_REG_1_ & n77475;
  assign n77477 = ~n77464 & n77466;
  assign n77478 = ~n77463 & ~n77477;
  assign n77479 = P3_DATAO_REG_2_ & n77438;
  assign n77480 = P3_DATAO_REG_3_ & n77440;
  assign n77481 = P3_DATAO_REG_5_ & n77444;
  assign n77482 = P3_DATAO_REG_4_ & n77442;
  assign n77483 = n77481 & ~n77482;
  assign n77484 = ~n77481 & n77482;
  assign n77485 = ~n77483 & ~n77484;
  assign n77486 = n77480 & ~n77485;
  assign n77487 = ~n77480 & n77485;
  assign n77488 = P3_DATAO_REG_3_ & P3_DATAO_REG_4_;
  assign n77489 = n77451 & n77488;
  assign n77490 = ~n77486 & ~n77487;
  assign n77491 = ~n77489 & n77490;
  assign n77492 = n77487 & n77489;
  assign n77493 = n77480 & n77489;
  assign n77494 = ~n77485 & n77493;
  assign n77495 = ~n77491 & ~n77492;
  assign n77496 = ~n77494 & n77495;
  assign n77497 = n77479 & ~n77496;
  assign n77498 = ~n77479 & n77496;
  assign n77499 = ~n77497 & ~n77498;
  assign n77500 = n77478 & ~n77499;
  assign n77501 = ~n77479 & ~n77496;
  assign n77502 = ~n77478 & n77501;
  assign n77503 = ~n77478 & n77479;
  assign n77504 = n77496 & n77503;
  assign n77505 = ~n77500 & ~n77502;
  assign n77506 = ~n77504 & n77505;
  assign n77507 = n77476 & ~n77506;
  assign n77508 = ~n77476 & n77506;
  assign n77509 = ~n77507 & ~n77508;
  assign n77510 = n77474 & ~n77509;
  assign n77511 = n77476 & n77506;
  assign n77512 = ~n77476 & ~n77506;
  assign n77513 = ~n77511 & ~n77512;
  assign n77514 = ~n77474 & ~n77513;
  assign n77515 = ~n77510 & ~n77514;
  assign n77516 = n77437 & ~n77515;
  assign n77517 = ~n77437 & n77515;
  assign n77518 = P3_DATAO_REG_0_ & n77475;
  assign n77519 = P3_DATAO_REG_0_ & n77438;
  assign n77520 = ~n77449 & ~n77453;
  assign n77521 = ~n77452 & n77520;
  assign n77522 = n77452 & ~n77520;
  assign n77523 = ~n77521 & ~n77522;
  assign n77524 = n77519 & ~n77523;
  assign n77525 = ~n77519 & n77523;
  assign n77526 = P3_DATAO_REG_1_ & n77442;
  assign n77527 = P3_DATAO_REG_0_ & n77444;
  assign n77528 = n77526 & n77527;
  assign n77529 = P3_DATAO_REG_0_ & n77440;
  assign n77530 = n77528 & n77529;
  assign n77531 = ~n77528 & ~n77529;
  assign n77532 = P3_DATAO_REG_2_ & n77444;
  assign n77533 = n77526 & ~n77532;
  assign n77534 = ~n77526 & n77532;
  assign n77535 = ~n77533 & ~n77534;
  assign n77536 = ~n77531 & ~n77535;
  assign n77537 = ~n77530 & ~n77536;
  assign n77538 = ~n77525 & ~n77537;
  assign n77539 = ~n77524 & ~n77538;
  assign n77540 = n77518 & ~n77539;
  assign n77541 = ~n77439 & n77470;
  assign n77542 = ~n77471 & ~n77541;
  assign n77543 = n77455 & ~n77542;
  assign n77544 = ~n77439 & ~n77470;
  assign n77545 = ~n77455 & n77544;
  assign n77546 = n77456 & n77470;
  assign n77547 = ~n77543 & ~n77545;
  assign n77548 = ~n77546 & n77547;
  assign n77549 = ~n77518 & n77539;
  assign n77550 = n77548 & ~n77549;
  assign n77551 = ~n77540 & ~n77550;
  assign n77552 = ~n77517 & ~n77551;
  assign n77553 = ~n77516 & ~n77552;
  assign n77554 = n77435 & ~n77553;
  assign n77555 = ~n77474 & ~n77512;
  assign n77556 = ~n77511 & ~n77555;
  assign n77557 = P3_DATAO_REG_1_ & n77436;
  assign n77558 = P3_DATAO_REG_2_ & n77475;
  assign n77559 = ~n77480 & ~n77489;
  assign n77560 = ~n77485 & ~n77559;
  assign n77561 = ~n77493 & ~n77560;
  assign n77562 = P3_DATAO_REG_3_ & n77438;
  assign n77563 = P3_DATAO_REG_4_ & n77440;
  assign n77564 = P3_DATAO_REG_6_ & n77444;
  assign n77565 = P3_DATAO_REG_5_ & n77442;
  assign n77566 = n77564 & ~n77565;
  assign n77567 = ~n77564 & n77565;
  assign n77568 = ~n77566 & ~n77567;
  assign n77569 = n77563 & ~n77568;
  assign n77570 = ~n77563 & n77568;
  assign n77571 = P3_DATAO_REG_4_ & P3_DATAO_REG_5_;
  assign n77572 = n77451 & n77571;
  assign n77573 = ~n77569 & ~n77570;
  assign n77574 = ~n77572 & n77573;
  assign n77575 = n77570 & n77572;
  assign n77576 = n77563 & n77572;
  assign n77577 = ~n77568 & n77576;
  assign n77578 = ~n77574 & ~n77575;
  assign n77579 = ~n77577 & n77578;
  assign n77580 = n77562 & ~n77579;
  assign n77581 = ~n77562 & n77579;
  assign n77582 = ~n77580 & ~n77581;
  assign n77583 = n77561 & ~n77582;
  assign n77584 = ~n77562 & ~n77579;
  assign n77585 = ~n77561 & n77584;
  assign n77586 = ~n77561 & n77562;
  assign n77587 = n77579 & n77586;
  assign n77588 = ~n77583 & ~n77585;
  assign n77589 = ~n77587 & n77588;
  assign n77590 = n77558 & ~n77589;
  assign n77591 = ~n77558 & n77589;
  assign n77592 = ~n77590 & ~n77591;
  assign n77593 = ~n77478 & ~n77496;
  assign n77594 = ~n77497 & ~n77503;
  assign n77595 = ~n77593 & n77594;
  assign n77596 = ~n77592 & n77595;
  assign n77597 = ~n77558 & ~n77589;
  assign n77598 = ~n77595 & n77597;
  assign n77599 = n77558 & ~n77595;
  assign n77600 = n77589 & n77599;
  assign n77601 = ~n77596 & ~n77598;
  assign n77602 = ~n77600 & n77601;
  assign n77603 = n77557 & ~n77602;
  assign n77604 = ~n77557 & n77602;
  assign n77605 = ~n77603 & ~n77604;
  assign n77606 = n77556 & ~n77605;
  assign n77607 = ~n77557 & ~n77602;
  assign n77608 = ~n77556 & n77607;
  assign n77609 = ~n77556 & n77557;
  assign n77610 = n77602 & n77609;
  assign n77611 = ~n77606 & ~n77608;
  assign n77612 = ~n77610 & n77611;
  assign n77613 = ~n77435 & n77553;
  assign n77614 = n77612 & ~n77613;
  assign n77615 = ~n77554 & ~n77614;
  assign n77616 = ~n77556 & ~n77602;
  assign n77617 = ~n77603 & ~n77609;
  assign n77618 = ~n77616 & n77617;
  assign n77619 = P3_DATAO_REG_1_ & n77434;
  assign n77620 = ~n77558 & n77595;
  assign n77621 = n77589 & ~n77620;
  assign n77622 = ~n77599 & ~n77621;
  assign n77623 = P3_DATAO_REG_2_ & n77436;
  assign n77624 = P3_DATAO_REG_3_ & n77475;
  assign n77625 = ~n77563 & ~n77572;
  assign n77626 = ~n77568 & ~n77625;
  assign n77627 = ~n77576 & ~n77626;
  assign n77628 = P3_DATAO_REG_4_ & n77438;
  assign n77629 = P3_DATAO_REG_5_ & n77440;
  assign n77630 = P3_DATAO_REG_7_ & n77444;
  assign n77631 = P3_DATAO_REG_6_ & n77442;
  assign n77632 = n77630 & ~n77631;
  assign n77633 = ~n77630 & n77631;
  assign n77634 = ~n77632 & ~n77633;
  assign n77635 = n77629 & ~n77634;
  assign n77636 = ~n77629 & n77634;
  assign n77637 = P3_DATAO_REG_5_ & P3_DATAO_REG_6_;
  assign n77638 = n77451 & n77637;
  assign n77639 = ~n77635 & ~n77636;
  assign n77640 = ~n77638 & n77639;
  assign n77641 = n77636 & n77638;
  assign n77642 = n77629 & n77638;
  assign n77643 = ~n77634 & n77642;
  assign n77644 = ~n77640 & ~n77641;
  assign n77645 = ~n77643 & n77644;
  assign n77646 = n77628 & ~n77645;
  assign n77647 = ~n77628 & n77645;
  assign n77648 = ~n77646 & ~n77647;
  assign n77649 = n77627 & ~n77648;
  assign n77650 = ~n77628 & ~n77645;
  assign n77651 = ~n77627 & n77650;
  assign n77652 = ~n77627 & n77628;
  assign n77653 = n77645 & n77652;
  assign n77654 = ~n77649 & ~n77651;
  assign n77655 = ~n77653 & n77654;
  assign n77656 = n77624 & ~n77655;
  assign n77657 = ~n77624 & n77655;
  assign n77658 = ~n77656 & ~n77657;
  assign n77659 = ~n77561 & ~n77579;
  assign n77660 = ~n77580 & ~n77586;
  assign n77661 = ~n77659 & n77660;
  assign n77662 = ~n77658 & n77661;
  assign n77663 = ~n77624 & ~n77655;
  assign n77664 = ~n77661 & n77663;
  assign n77665 = n77624 & ~n77661;
  assign n77666 = n77655 & n77665;
  assign n77667 = ~n77662 & ~n77664;
  assign n77668 = ~n77666 & n77667;
  assign n77669 = n77623 & ~n77668;
  assign n77670 = ~n77623 & n77668;
  assign n77671 = ~n77669 & ~n77670;
  assign n77672 = n77622 & ~n77671;
  assign n77673 = ~n77623 & ~n77668;
  assign n77674 = ~n77622 & n77673;
  assign n77675 = ~n77622 & n77623;
  assign n77676 = n77668 & n77675;
  assign n77677 = ~n77672 & ~n77674;
  assign n77678 = ~n77676 & n77677;
  assign n77679 = n77619 & ~n77678;
  assign n77680 = ~n77619 & n77678;
  assign n77681 = ~n77679 & ~n77680;
  assign n77682 = n77618 & ~n77681;
  assign n77683 = n77619 & n77678;
  assign n77684 = ~n77619 & ~n77678;
  assign n77685 = ~n77683 & ~n77684;
  assign n77686 = ~n77618 & ~n77685;
  assign n77687 = ~n77682 & ~n77686;
  assign n77688 = ~SEL & DIN_7_;
  assign n77689 = P3_DATAO_REG_0_ & n77688;
  assign n77690 = ~n77687 & ~n77689;
  assign n77691 = n77687 & n77689;
  assign n77692 = ~n77690 & ~n77691;
  assign n77693 = n77615 & ~n77692;
  assign n77694 = n77687 & ~n77689;
  assign n77695 = ~n77687 & n77689;
  assign n77696 = ~n77694 & ~n77695;
  assign n77697 = ~n77615 & ~n77696;
  assign n77698 = ~n77693 & ~n77697;
  assign n77699 = ~n12802 & ~n77698;
  assign n77700 = ~n77433 & ~n77699;
  assign n77701 = n77374 & ~n77700;
  assign n77702 = n77432 & n77701;
  assign n77703 = P2_BUF1_REG_23_ & n12802;
  assign n77704 = ~SEL & DIN_23_;
  assign n77705 = P3_DATAO_REG_0_ & n77704;
  assign n77706 = ~SEL & DIN_21_;
  assign n77707 = P3_DATAO_REG_1_ & n77706;
  assign n77708 = ~SEL & DIN_20_;
  assign n77709 = P3_DATAO_REG_1_ & n77708;
  assign n77710 = ~SEL & DIN_19_;
  assign n77711 = P3_DATAO_REG_1_ & n77710;
  assign n77712 = ~SEL & DIN_18_;
  assign n77713 = P3_DATAO_REG_2_ & n77712;
  assign n77714 = ~SEL & DIN_17_;
  assign n77715 = P3_DATAO_REG_2_ & n77714;
  assign n77716 = ~SEL & DIN_15_;
  assign n77717 = P3_DATAO_REG_4_ & n77716;
  assign n77718 = ~SEL & DIN_14_;
  assign n77719 = P3_DATAO_REG_4_ & n77718;
  assign n77720 = ~SEL & DIN_13_;
  assign n77721 = P3_DATAO_REG_5_ & n77720;
  assign n77722 = ~SEL & DIN_12_;
  assign n77723 = P3_DATAO_REG_5_ & n77722;
  assign n77724 = ~SEL & DIN_11_;
  assign n77725 = P3_DATAO_REG_6_ & n77724;
  assign n77726 = ~SEL & DIN_10_;
  assign n77727 = P3_DATAO_REG_6_ & n77726;
  assign n77728 = P3_DATAO_REG_13_ & n77438;
  assign n77729 = P3_DATAO_REG_13_ & n77440;
  assign n77730 = P3_DATAO_REG_14_ & n77442;
  assign n77731 = P3_DATAO_REG_15_ & n77444;
  assign n77732 = n77730 & ~n77731;
  assign n77733 = ~n77730 & n77731;
  assign n77734 = ~n77732 & ~n77733;
  assign n77735 = n77729 & ~n77734;
  assign n77736 = P3_DATAO_REG_13_ & P3_DATAO_REG_14_;
  assign n77737 = n77451 & n77736;
  assign n77738 = ~n77729 & n77734;
  assign n77739 = n77737 & ~n77738;
  assign n77740 = ~n77735 & ~n77739;
  assign n77741 = n77728 & ~n77740;
  assign n77742 = ~n77728 & n77740;
  assign n77743 = ~n77741 & ~n77742;
  assign n77744 = P3_DATAO_REG_14_ & n77440;
  assign n77745 = P3_DATAO_REG_15_ & n77442;
  assign n77746 = P3_DATAO_REG_16_ & n77444;
  assign n77747 = n77745 & ~n77746;
  assign n77748 = ~n77745 & n77746;
  assign n77749 = ~n77747 & ~n77748;
  assign n77750 = n77744 & ~n77749;
  assign n77751 = ~n77744 & n77749;
  assign n77752 = P3_DATAO_REG_14_ & P3_DATAO_REG_15_;
  assign n77753 = n77451 & n77752;
  assign n77754 = ~n77750 & ~n77751;
  assign n77755 = ~n77753 & n77754;
  assign n77756 = n77753 & ~n77754;
  assign n77757 = ~n77755 & ~n77756;
  assign n77758 = ~n77743 & n77757;
  assign n77759 = n77743 & ~n77757;
  assign n77760 = ~n77758 & ~n77759;
  assign n77761 = P3_DATAO_REG_12_ & n77475;
  assign n77762 = ~n77760 & ~n77761;
  assign n77763 = n77760 & n77761;
  assign n77764 = P3_DATAO_REG_12_ & n77438;
  assign n77765 = P3_DATAO_REG_12_ & n77440;
  assign n77766 = P3_DATAO_REG_13_ & n77442;
  assign n77767 = P3_DATAO_REG_14_ & n77444;
  assign n77768 = n77766 & ~n77767;
  assign n77769 = ~n77766 & n77767;
  assign n77770 = ~n77768 & ~n77769;
  assign n77771 = n77765 & ~n77770;
  assign n77772 = P3_DATAO_REG_12_ & P3_DATAO_REG_13_;
  assign n77773 = n77451 & n77772;
  assign n77774 = ~n77765 & n77770;
  assign n77775 = n77773 & ~n77774;
  assign n77776 = ~n77771 & ~n77775;
  assign n77777 = n77764 & ~n77776;
  assign n77778 = ~n77735 & ~n77738;
  assign n77779 = ~n77737 & n77778;
  assign n77780 = n77737 & ~n77778;
  assign n77781 = ~n77779 & ~n77780;
  assign n77782 = n77764 & ~n77781;
  assign n77783 = ~n77776 & ~n77781;
  assign n77784 = ~n77777 & ~n77782;
  assign n77785 = ~n77783 & n77784;
  assign n77786 = ~n77762 & ~n77763;
  assign n77787 = n77785 & n77786;
  assign n77788 = ~n77785 & ~n77786;
  assign n77789 = ~n77787 & ~n77788;
  assign n77790 = P3_DATAO_REG_11_ & n77436;
  assign n77791 = n77789 & n77790;
  assign n77792 = ~n77789 & ~n77790;
  assign n77793 = ~n77791 & ~n77792;
  assign n77794 = P3_DATAO_REG_11_ & n77475;
  assign n77795 = ~n77764 & n77781;
  assign n77796 = ~n77782 & ~n77795;
  assign n77797 = n77776 & ~n77796;
  assign n77798 = ~n77764 & ~n77781;
  assign n77799 = ~n77776 & n77798;
  assign n77800 = n77777 & n77781;
  assign n77801 = ~n77797 & ~n77799;
  assign n77802 = ~n77800 & n77801;
  assign n77803 = n77794 & n77802;
  assign n77804 = ~n77794 & ~n77802;
  assign n77805 = P3_DATAO_REG_11_ & n77438;
  assign n77806 = P3_DATAO_REG_11_ & n77440;
  assign n77807 = P3_DATAO_REG_12_ & n77442;
  assign n77808 = P3_DATAO_REG_13_ & n77444;
  assign n77809 = n77807 & ~n77808;
  assign n77810 = ~n77807 & n77808;
  assign n77811 = ~n77809 & ~n77810;
  assign n77812 = n77806 & ~n77811;
  assign n77813 = P3_DATAO_REG_11_ & P3_DATAO_REG_12_;
  assign n77814 = n77451 & n77813;
  assign n77815 = ~n77806 & n77811;
  assign n77816 = n77814 & ~n77815;
  assign n77817 = ~n77812 & ~n77816;
  assign n77818 = n77805 & ~n77817;
  assign n77819 = ~n77771 & ~n77774;
  assign n77820 = ~n77773 & n77819;
  assign n77821 = n77773 & ~n77819;
  assign n77822 = ~n77820 & ~n77821;
  assign n77823 = n77805 & ~n77822;
  assign n77824 = ~n77817 & ~n77822;
  assign n77825 = ~n77818 & ~n77823;
  assign n77826 = ~n77824 & n77825;
  assign n77827 = ~n77804 & ~n77826;
  assign n77828 = ~n77803 & ~n77827;
  assign n77829 = ~n77793 & ~n77828;
  assign n77830 = n77793 & n77828;
  assign n77831 = ~n77829 & ~n77830;
  assign n77832 = P3_DATAO_REG_10_ & n77434;
  assign n77833 = ~n77831 & ~n77832;
  assign n77834 = n77831 & n77832;
  assign n77835 = P3_DATAO_REG_10_ & n77436;
  assign n77836 = P3_DATAO_REG_10_ & n77475;
  assign n77837 = ~n77805 & n77822;
  assign n77838 = ~n77823 & ~n77837;
  assign n77839 = n77817 & ~n77838;
  assign n77840 = ~n77805 & ~n77822;
  assign n77841 = ~n77817 & n77840;
  assign n77842 = n77818 & n77822;
  assign n77843 = ~n77839 & ~n77841;
  assign n77844 = ~n77842 & n77843;
  assign n77845 = n77836 & n77844;
  assign n77846 = ~n77836 & ~n77844;
  assign n77847 = P3_DATAO_REG_10_ & n77438;
  assign n77848 = P3_DATAO_REG_10_ & n77440;
  assign n77849 = P3_DATAO_REG_11_ & n77442;
  assign n77850 = P3_DATAO_REG_12_ & n77444;
  assign n77851 = n77849 & ~n77850;
  assign n77852 = ~n77849 & n77850;
  assign n77853 = ~n77851 & ~n77852;
  assign n77854 = n77848 & ~n77853;
  assign n77855 = P3_DATAO_REG_10_ & P3_DATAO_REG_11_;
  assign n77856 = n77451 & n77855;
  assign n77857 = ~n77848 & n77853;
  assign n77858 = n77856 & ~n77857;
  assign n77859 = ~n77854 & ~n77858;
  assign n77860 = n77847 & ~n77859;
  assign n77861 = ~n77812 & ~n77815;
  assign n77862 = ~n77814 & n77861;
  assign n77863 = n77814 & ~n77861;
  assign n77864 = ~n77862 & ~n77863;
  assign n77865 = n77847 & ~n77864;
  assign n77866 = ~n77859 & ~n77864;
  assign n77867 = ~n77860 & ~n77865;
  assign n77868 = ~n77866 & n77867;
  assign n77869 = ~n77846 & ~n77868;
  assign n77870 = ~n77845 & ~n77869;
  assign n77871 = n77835 & ~n77870;
  assign n77872 = n77794 & ~n77802;
  assign n77873 = ~n77794 & n77802;
  assign n77874 = ~n77872 & ~n77873;
  assign n77875 = n77826 & ~n77874;
  assign n77876 = ~n77803 & ~n77804;
  assign n77877 = ~n77826 & ~n77876;
  assign n77878 = ~n77875 & ~n77877;
  assign n77879 = n77835 & ~n77878;
  assign n77880 = ~n77870 & ~n77878;
  assign n77881 = ~n77871 & ~n77879;
  assign n77882 = ~n77880 & n77881;
  assign n77883 = ~n77833 & ~n77834;
  assign n77884 = n77882 & n77883;
  assign n77885 = ~n77882 & ~n77883;
  assign n77886 = ~n77884 & ~n77885;
  assign n77887 = P3_DATAO_REG_9_ & n77688;
  assign n77888 = n77886 & n77887;
  assign n77889 = ~n77886 & ~n77887;
  assign n77890 = ~n77888 & ~n77889;
  assign n77891 = ~n77835 & n77878;
  assign n77892 = ~n77879 & ~n77891;
  assign n77893 = n77870 & ~n77892;
  assign n77894 = ~n77835 & ~n77878;
  assign n77895 = ~n77870 & n77894;
  assign n77896 = n77871 & n77878;
  assign n77897 = ~n77893 & ~n77895;
  assign n77898 = ~n77896 & n77897;
  assign n77899 = P3_DATAO_REG_9_ & n77434;
  assign n77900 = n77898 & n77899;
  assign n77901 = ~n77898 & ~n77899;
  assign n77902 = P3_DATAO_REG_9_ & n77436;
  assign n77903 = ~n77847 & n77864;
  assign n77904 = ~n77865 & ~n77903;
  assign n77905 = n77859 & ~n77904;
  assign n77906 = ~n77847 & ~n77864;
  assign n77907 = ~n77859 & n77906;
  assign n77908 = n77860 & n77864;
  assign n77909 = ~n77905 & ~n77907;
  assign n77910 = ~n77908 & n77909;
  assign n77911 = P3_DATAO_REG_9_ & n77475;
  assign n77912 = n77910 & n77911;
  assign n77913 = ~n77910 & ~n77911;
  assign n77914 = P3_DATAO_REG_9_ & n77438;
  assign n77915 = P3_DATAO_REG_9_ & n77440;
  assign n77916 = P3_DATAO_REG_10_ & n77442;
  assign n77917 = P3_DATAO_REG_11_ & n77444;
  assign n77918 = n77916 & ~n77917;
  assign n77919 = ~n77916 & n77917;
  assign n77920 = ~n77918 & ~n77919;
  assign n77921 = n77915 & ~n77920;
  assign n77922 = P3_DATAO_REG_9_ & P3_DATAO_REG_10_;
  assign n77923 = n77451 & n77922;
  assign n77924 = ~n77915 & n77920;
  assign n77925 = n77923 & ~n77924;
  assign n77926 = ~n77921 & ~n77925;
  assign n77927 = n77914 & ~n77926;
  assign n77928 = ~n77854 & ~n77857;
  assign n77929 = ~n77856 & n77928;
  assign n77930 = n77856 & ~n77928;
  assign n77931 = ~n77929 & ~n77930;
  assign n77932 = n77914 & ~n77931;
  assign n77933 = ~n77926 & ~n77931;
  assign n77934 = ~n77927 & ~n77932;
  assign n77935 = ~n77933 & n77934;
  assign n77936 = ~n77913 & ~n77935;
  assign n77937 = ~n77912 & ~n77936;
  assign n77938 = n77902 & ~n77937;
  assign n77939 = n77836 & ~n77844;
  assign n77940 = ~n77836 & n77844;
  assign n77941 = ~n77939 & ~n77940;
  assign n77942 = n77868 & ~n77941;
  assign n77943 = ~n77845 & ~n77846;
  assign n77944 = ~n77868 & ~n77943;
  assign n77945 = ~n77942 & ~n77944;
  assign n77946 = n77902 & ~n77945;
  assign n77947 = ~n77937 & ~n77945;
  assign n77948 = ~n77938 & ~n77946;
  assign n77949 = ~n77947 & n77948;
  assign n77950 = ~n77901 & ~n77949;
  assign n77951 = ~n77900 & ~n77950;
  assign n77952 = ~n77890 & ~n77951;
  assign n77953 = n77890 & n77951;
  assign n77954 = ~n77952 & ~n77953;
  assign n77955 = ~SEL & DIN_8_;
  assign n77956 = P3_DATAO_REG_8_ & n77955;
  assign n77957 = ~n77954 & ~n77956;
  assign n77958 = n77954 & n77956;
  assign n77959 = P3_DATAO_REG_8_ & n77688;
  assign n77960 = ~n77898 & n77899;
  assign n77961 = n77898 & ~n77899;
  assign n77962 = ~n77960 & ~n77961;
  assign n77963 = n77949 & ~n77962;
  assign n77964 = ~n77900 & ~n77901;
  assign n77965 = ~n77949 & ~n77964;
  assign n77966 = ~n77963 & ~n77965;
  assign n77967 = n77959 & ~n77966;
  assign n77968 = ~n77959 & n77966;
  assign n77969 = P3_DATAO_REG_8_ & n77434;
  assign n77970 = P3_DATAO_REG_8_ & n77436;
  assign n77971 = ~n77910 & n77911;
  assign n77972 = n77910 & ~n77911;
  assign n77973 = ~n77971 & ~n77972;
  assign n77974 = n77935 & ~n77973;
  assign n77975 = ~n77912 & ~n77913;
  assign n77976 = ~n77935 & ~n77975;
  assign n77977 = ~n77974 & ~n77976;
  assign n77978 = n77970 & ~n77977;
  assign n77979 = ~n77914 & n77931;
  assign n77980 = ~n77932 & ~n77979;
  assign n77981 = n77926 & ~n77980;
  assign n77982 = ~n77914 & ~n77931;
  assign n77983 = ~n77926 & n77982;
  assign n77984 = n77927 & n77931;
  assign n77985 = ~n77981 & ~n77983;
  assign n77986 = ~n77984 & n77985;
  assign n77987 = P3_DATAO_REG_8_ & n77475;
  assign n77988 = n77986 & n77987;
  assign n77989 = ~n77986 & ~n77987;
  assign n77990 = P3_DATAO_REG_8_ & n77438;
  assign n77991 = P3_DATAO_REG_8_ & n77440;
  assign n77992 = P3_DATAO_REG_9_ & n77442;
  assign n77993 = P3_DATAO_REG_10_ & n77444;
  assign n77994 = n77992 & ~n77993;
  assign n77995 = ~n77992 & n77993;
  assign n77996 = ~n77994 & ~n77995;
  assign n77997 = n77991 & ~n77996;
  assign n77998 = P3_DATAO_REG_8_ & P3_DATAO_REG_9_;
  assign n77999 = n77451 & n77998;
  assign n78000 = ~n77991 & n77996;
  assign n78001 = n77999 & ~n78000;
  assign n78002 = ~n77997 & ~n78001;
  assign n78003 = n77990 & ~n78002;
  assign n78004 = ~n77921 & ~n77924;
  assign n78005 = ~n77923 & n78004;
  assign n78006 = n77923 & ~n78004;
  assign n78007 = ~n78005 & ~n78006;
  assign n78008 = n77990 & ~n78007;
  assign n78009 = ~n78002 & ~n78007;
  assign n78010 = ~n78003 & ~n78008;
  assign n78011 = ~n78009 & n78010;
  assign n78012 = ~n77989 & ~n78011;
  assign n78013 = ~n77988 & ~n78012;
  assign n78014 = n77970 & ~n78013;
  assign n78015 = ~n77977 & ~n78013;
  assign n78016 = ~n77978 & ~n78014;
  assign n78017 = ~n78015 & n78016;
  assign n78018 = n77969 & ~n78017;
  assign n78019 = ~n77902 & n77945;
  assign n78020 = ~n77946 & ~n78019;
  assign n78021 = n77937 & ~n78020;
  assign n78022 = ~n77902 & ~n77945;
  assign n78023 = ~n77937 & n78022;
  assign n78024 = n77938 & n77945;
  assign n78025 = ~n78021 & ~n78023;
  assign n78026 = ~n78024 & n78025;
  assign n78027 = ~n77969 & n78017;
  assign n78028 = n78026 & ~n78027;
  assign n78029 = ~n78018 & ~n78028;
  assign n78030 = ~n77968 & ~n78029;
  assign n78031 = ~n77967 & ~n78030;
  assign n78032 = ~n77957 & ~n77958;
  assign n78033 = n78031 & n78032;
  assign n78034 = ~n78031 & ~n78032;
  assign n78035 = ~n78033 & ~n78034;
  assign n78036 = ~SEL & DIN_9_;
  assign n78037 = P3_DATAO_REG_7_ & n78036;
  assign n78038 = n78035 & n78037;
  assign n78039 = ~n78035 & ~n78037;
  assign n78040 = ~n78038 & ~n78039;
  assign n78041 = P3_DATAO_REG_7_ & n77955;
  assign n78042 = n77959 & ~n78029;
  assign n78043 = ~n77959 & n78029;
  assign n78044 = ~n78042 & ~n78043;
  assign n78045 = n77966 & ~n78044;
  assign n78046 = ~n77966 & n78044;
  assign n78047 = ~n78045 & ~n78046;
  assign n78048 = n78041 & n78047;
  assign n78049 = ~n78041 & ~n78047;
  assign n78050 = P3_DATAO_REG_7_ & n77688;
  assign n78051 = ~n77970 & n78013;
  assign n78052 = ~n78014 & ~n78051;
  assign n78053 = n77977 & ~n78052;
  assign n78054 = ~n77970 & ~n78013;
  assign n78055 = ~n77977 & n78054;
  assign n78056 = n77978 & n78013;
  assign n78057 = ~n78053 & ~n78055;
  assign n78058 = ~n78056 & n78057;
  assign n78059 = P3_DATAO_REG_7_ & n77434;
  assign n78060 = n78058 & n78059;
  assign n78061 = ~n78058 & ~n78059;
  assign n78062 = P3_DATAO_REG_7_ & n77436;
  assign n78063 = ~n77990 & n78007;
  assign n78064 = ~n78008 & ~n78063;
  assign n78065 = n78002 & ~n78064;
  assign n78066 = ~n77990 & ~n78007;
  assign n78067 = ~n78002 & n78066;
  assign n78068 = n78003 & n78007;
  assign n78069 = ~n78065 & ~n78067;
  assign n78070 = ~n78068 & n78069;
  assign n78071 = P3_DATAO_REG_7_ & n77475;
  assign n78072 = n78070 & n78071;
  assign n78073 = ~n78070 & ~n78071;
  assign n78074 = P3_DATAO_REG_7_ & n77438;
  assign n78075 = P3_DATAO_REG_7_ & P3_DATAO_REG_8_;
  assign n78076 = n77451 & n78075;
  assign n78077 = P3_DATAO_REG_7_ & n77440;
  assign n78078 = n78076 & n78077;
  assign n78079 = ~n78076 & ~n78077;
  assign n78080 = P3_DATAO_REG_9_ & n77444;
  assign n78081 = P3_DATAO_REG_8_ & n77442;
  assign n78082 = n78080 & ~n78081;
  assign n78083 = ~n78080 & n78081;
  assign n78084 = ~n78082 & ~n78083;
  assign n78085 = ~n78079 & ~n78084;
  assign n78086 = ~n78078 & ~n78085;
  assign n78087 = n78074 & ~n78086;
  assign n78088 = ~n77997 & ~n78000;
  assign n78089 = ~n77999 & n78088;
  assign n78090 = n77999 & ~n78088;
  assign n78091 = ~n78089 & ~n78090;
  assign n78092 = n78074 & ~n78091;
  assign n78093 = ~n78086 & ~n78091;
  assign n78094 = ~n78087 & ~n78092;
  assign n78095 = ~n78093 & n78094;
  assign n78096 = ~n78073 & ~n78095;
  assign n78097 = ~n78072 & ~n78096;
  assign n78098 = n78062 & ~n78097;
  assign n78099 = ~n77986 & n77987;
  assign n78100 = n77986 & ~n77987;
  assign n78101 = ~n78099 & ~n78100;
  assign n78102 = n78011 & ~n78101;
  assign n78103 = ~n77988 & ~n77989;
  assign n78104 = ~n78011 & ~n78103;
  assign n78105 = ~n78102 & ~n78104;
  assign n78106 = n78062 & ~n78105;
  assign n78107 = ~n78097 & ~n78105;
  assign n78108 = ~n78098 & ~n78106;
  assign n78109 = ~n78107 & n78108;
  assign n78110 = ~n78061 & ~n78109;
  assign n78111 = ~n78060 & ~n78110;
  assign n78112 = n78050 & ~n78111;
  assign n78113 = ~n78018 & ~n78027;
  assign n78114 = ~n78026 & n78113;
  assign n78115 = n78026 & ~n78113;
  assign n78116 = ~n78114 & ~n78115;
  assign n78117 = n78050 & ~n78116;
  assign n78118 = ~n78111 & ~n78116;
  assign n78119 = ~n78112 & ~n78117;
  assign n78120 = ~n78118 & n78119;
  assign n78121 = ~n78049 & ~n78120;
  assign n78122 = ~n78048 & ~n78121;
  assign n78123 = ~n78040 & ~n78122;
  assign n78124 = n78040 & n78122;
  assign n78125 = ~n78123 & ~n78124;
  assign n78126 = n77727 & n78125;
  assign n78127 = ~n77727 & ~n78125;
  assign n78128 = P3_DATAO_REG_6_ & n78036;
  assign n78129 = ~n78050 & n78116;
  assign n78130 = ~n78117 & ~n78129;
  assign n78131 = n78111 & ~n78130;
  assign n78132 = ~n78050 & ~n78116;
  assign n78133 = ~n78111 & n78132;
  assign n78134 = n78112 & n78116;
  assign n78135 = ~n78131 & ~n78133;
  assign n78136 = ~n78134 & n78135;
  assign n78137 = P3_DATAO_REG_6_ & n77955;
  assign n78138 = n78136 & n78137;
  assign n78139 = ~n78136 & ~n78137;
  assign n78140 = P3_DATAO_REG_6_ & n77688;
  assign n78141 = ~n78058 & n78059;
  assign n78142 = n78058 & ~n78059;
  assign n78143 = ~n78141 & ~n78142;
  assign n78144 = n78109 & ~n78143;
  assign n78145 = ~n78060 & ~n78061;
  assign n78146 = ~n78109 & ~n78145;
  assign n78147 = ~n78144 & ~n78146;
  assign n78148 = n78140 & ~n78147;
  assign n78149 = ~n78062 & n78105;
  assign n78150 = ~n78106 & ~n78149;
  assign n78151 = n78097 & ~n78150;
  assign n78152 = ~n78062 & ~n78105;
  assign n78153 = ~n78097 & n78152;
  assign n78154 = n78098 & n78105;
  assign n78155 = ~n78151 & ~n78153;
  assign n78156 = ~n78154 & n78155;
  assign n78157 = P3_DATAO_REG_6_ & n77434;
  assign n78158 = n78156 & n78157;
  assign n78159 = ~n78156 & ~n78157;
  assign n78160 = P3_DATAO_REG_6_ & n77436;
  assign n78161 = ~n78070 & n78071;
  assign n78162 = n78070 & ~n78071;
  assign n78163 = ~n78161 & ~n78162;
  assign n78164 = n78095 & ~n78163;
  assign n78165 = ~n78072 & ~n78073;
  assign n78166 = ~n78095 & ~n78165;
  assign n78167 = ~n78164 & ~n78166;
  assign n78168 = n78160 & ~n78167;
  assign n78169 = ~n78074 & n78091;
  assign n78170 = ~n78092 & ~n78169;
  assign n78171 = n78086 & ~n78170;
  assign n78172 = ~n78074 & ~n78091;
  assign n78173 = ~n78086 & n78172;
  assign n78174 = n78087 & n78091;
  assign n78175 = ~n78171 & ~n78173;
  assign n78176 = ~n78174 & n78175;
  assign n78177 = P3_DATAO_REG_6_ & n77475;
  assign n78178 = n78176 & n78177;
  assign n78179 = ~n78176 & ~n78177;
  assign n78180 = P3_DATAO_REG_6_ & n77438;
  assign n78181 = n78077 & ~n78084;
  assign n78182 = ~n78077 & n78084;
  assign n78183 = ~n78181 & ~n78182;
  assign n78184 = ~n78076 & n78183;
  assign n78185 = n78076 & n78182;
  assign n78186 = n78078 & ~n78084;
  assign n78187 = ~n78184 & ~n78185;
  assign n78188 = ~n78186 & n78187;
  assign n78189 = n78180 & ~n78188;
  assign n78190 = P3_DATAO_REG_6_ & P3_DATAO_REG_7_;
  assign n78191 = n77451 & n78190;
  assign n78192 = P3_DATAO_REG_6_ & n77440;
  assign n78193 = n78191 & n78192;
  assign n78194 = ~n78191 & ~n78192;
  assign n78195 = P3_DATAO_REG_8_ & n77444;
  assign n78196 = P3_DATAO_REG_7_ & n77442;
  assign n78197 = n78195 & ~n78196;
  assign n78198 = ~n78195 & n78196;
  assign n78199 = ~n78197 & ~n78198;
  assign n78200 = ~n78194 & ~n78199;
  assign n78201 = ~n78193 & ~n78200;
  assign n78202 = n78180 & ~n78201;
  assign n78203 = ~n78188 & ~n78201;
  assign n78204 = ~n78189 & ~n78202;
  assign n78205 = ~n78203 & n78204;
  assign n78206 = ~n78179 & ~n78205;
  assign n78207 = ~n78178 & ~n78206;
  assign n78208 = n78160 & ~n78207;
  assign n78209 = ~n78167 & ~n78207;
  assign n78210 = ~n78168 & ~n78208;
  assign n78211 = ~n78209 & n78210;
  assign n78212 = ~n78159 & ~n78211;
  assign n78213 = ~n78158 & ~n78212;
  assign n78214 = n78140 & ~n78213;
  assign n78215 = ~n78147 & ~n78213;
  assign n78216 = ~n78148 & ~n78214;
  assign n78217 = ~n78215 & n78216;
  assign n78218 = ~n78139 & ~n78217;
  assign n78219 = ~n78138 & ~n78218;
  assign n78220 = n78128 & ~n78219;
  assign n78221 = ~n78048 & ~n78049;
  assign n78222 = n78120 & n78221;
  assign n78223 = ~n78120 & ~n78221;
  assign n78224 = ~n78222 & ~n78223;
  assign n78225 = n78128 & ~n78224;
  assign n78226 = ~n78219 & ~n78224;
  assign n78227 = ~n78220 & ~n78225;
  assign n78228 = ~n78226 & n78227;
  assign n78229 = ~n78127 & ~n78228;
  assign n78230 = ~n78126 & ~n78229;
  assign n78231 = n77725 & ~n78230;
  assign n78232 = ~n77725 & n78230;
  assign n78233 = ~n78231 & ~n78232;
  assign n78234 = ~n78035 & n78037;
  assign n78235 = n78035 & ~n78037;
  assign n78236 = ~n78122 & ~n78235;
  assign n78237 = ~n78234 & ~n78236;
  assign n78238 = P3_DATAO_REG_7_ & n77726;
  assign n78239 = ~n77957 & ~n78031;
  assign n78240 = ~n77958 & ~n78239;
  assign n78241 = P3_DATAO_REG_8_ & n78036;
  assign n78242 = P3_DATAO_REG_9_ & n77955;
  assign n78243 = ~n77886 & n77887;
  assign n78244 = n77886 & ~n77887;
  assign n78245 = ~n77951 & ~n78244;
  assign n78246 = ~n78243 & ~n78245;
  assign n78247 = n78242 & ~n78246;
  assign n78248 = ~n78242 & n78246;
  assign n78249 = ~n78247 & ~n78248;
  assign n78250 = ~n77833 & ~n77882;
  assign n78251 = ~n77834 & ~n78250;
  assign n78252 = P3_DATAO_REG_10_ & n77688;
  assign n78253 = ~n77789 & n77790;
  assign n78254 = n77789 & ~n77790;
  assign n78255 = ~n77828 & ~n78254;
  assign n78256 = ~n78253 & ~n78255;
  assign n78257 = P3_DATAO_REG_11_ & n77434;
  assign n78258 = ~n77762 & ~n77785;
  assign n78259 = ~n77763 & ~n78258;
  assign n78260 = P3_DATAO_REG_12_ & n77436;
  assign n78261 = n77728 & ~n77757;
  assign n78262 = ~n77728 & n77757;
  assign n78263 = ~n77740 & ~n78262;
  assign n78264 = ~n78261 & ~n78263;
  assign n78265 = P3_DATAO_REG_13_ & n77475;
  assign n78266 = ~n77751 & n77753;
  assign n78267 = ~n77750 & ~n78266;
  assign n78268 = P3_DATAO_REG_14_ & n77438;
  assign n78269 = P3_DATAO_REG_16_ & n77442;
  assign n78270 = P3_DATAO_REG_17_ & n77444;
  assign n78271 = n78269 & ~n78270;
  assign n78272 = ~n78269 & n78270;
  assign n78273 = ~n78271 & ~n78272;
  assign n78274 = P3_DATAO_REG_15_ & n77440;
  assign n78275 = P3_DATAO_REG_15_ & P3_DATAO_REG_16_;
  assign n78276 = n77451 & n78275;
  assign n78277 = n78274 & ~n78276;
  assign n78278 = ~n78274 & n78276;
  assign n78279 = ~n78277 & ~n78278;
  assign n78280 = n78273 & ~n78279;
  assign n78281 = ~n78274 & ~n78276;
  assign n78282 = n78274 & n78276;
  assign n78283 = ~n78281 & ~n78282;
  assign n78284 = ~n78273 & ~n78283;
  assign n78285 = ~n78280 & ~n78284;
  assign n78286 = n78268 & ~n78285;
  assign n78287 = ~n78268 & n78285;
  assign n78288 = ~n78286 & ~n78287;
  assign n78289 = n78267 & ~n78288;
  assign n78290 = ~n78268 & ~n78285;
  assign n78291 = ~n78267 & n78290;
  assign n78292 = ~n78267 & n78268;
  assign n78293 = n78285 & n78292;
  assign n78294 = ~n78289 & ~n78291;
  assign n78295 = ~n78293 & n78294;
  assign n78296 = n78265 & ~n78295;
  assign n78297 = ~n78265 & n78295;
  assign n78298 = ~n78296 & ~n78297;
  assign n78299 = n78264 & ~n78298;
  assign n78300 = n78265 & n78295;
  assign n78301 = ~n78265 & ~n78295;
  assign n78302 = ~n78300 & ~n78301;
  assign n78303 = ~n78264 & ~n78302;
  assign n78304 = ~n78299 & ~n78303;
  assign n78305 = n78260 & ~n78304;
  assign n78306 = ~n78260 & n78304;
  assign n78307 = ~n78305 & ~n78306;
  assign n78308 = n78259 & ~n78307;
  assign n78309 = ~n78260 & ~n78304;
  assign n78310 = ~n78259 & n78309;
  assign n78311 = ~n78259 & n78260;
  assign n78312 = n78304 & n78311;
  assign n78313 = ~n78308 & ~n78310;
  assign n78314 = ~n78312 & n78313;
  assign n78315 = n78257 & ~n78314;
  assign n78316 = ~n78257 & n78314;
  assign n78317 = ~n78315 & ~n78316;
  assign n78318 = n78256 & ~n78317;
  assign n78319 = n78257 & n78314;
  assign n78320 = ~n78257 & ~n78314;
  assign n78321 = ~n78319 & ~n78320;
  assign n78322 = ~n78256 & ~n78321;
  assign n78323 = ~n78318 & ~n78322;
  assign n78324 = n78252 & ~n78323;
  assign n78325 = ~n78252 & n78323;
  assign n78326 = ~n78324 & ~n78325;
  assign n78327 = n78251 & ~n78326;
  assign n78328 = ~n78252 & ~n78323;
  assign n78329 = ~n78251 & n78328;
  assign n78330 = ~n78251 & n78252;
  assign n78331 = n78323 & n78330;
  assign n78332 = ~n78327 & ~n78329;
  assign n78333 = ~n78331 & n78332;
  assign n78334 = ~n78249 & ~n78333;
  assign n78335 = n78249 & n78333;
  assign n78336 = ~n78334 & ~n78335;
  assign n78337 = n78241 & n78336;
  assign n78338 = ~n78241 & ~n78336;
  assign n78339 = ~n78337 & ~n78338;
  assign n78340 = n78240 & ~n78339;
  assign n78341 = ~n78241 & n78336;
  assign n78342 = ~n78240 & n78341;
  assign n78343 = ~n78240 & n78241;
  assign n78344 = ~n78336 & n78343;
  assign n78345 = ~n78340 & ~n78342;
  assign n78346 = ~n78344 & n78345;
  assign n78347 = n78238 & ~n78346;
  assign n78348 = ~n78238 & n78346;
  assign n78349 = ~n78347 & ~n78348;
  assign n78350 = n78237 & ~n78349;
  assign n78351 = n78238 & n78346;
  assign n78352 = ~n78238 & ~n78346;
  assign n78353 = ~n78351 & ~n78352;
  assign n78354 = ~n78237 & ~n78353;
  assign n78355 = ~n78350 & ~n78354;
  assign n78356 = ~n78233 & n78355;
  assign n78357 = n78233 & ~n78355;
  assign n78358 = ~n78356 & ~n78357;
  assign n78359 = n77723 & n78358;
  assign n78360 = ~n77723 & ~n78358;
  assign n78361 = P3_DATAO_REG_5_ & n77724;
  assign n78362 = ~n78128 & n78224;
  assign n78363 = ~n78225 & ~n78362;
  assign n78364 = n78219 & ~n78363;
  assign n78365 = ~n78128 & ~n78224;
  assign n78366 = ~n78219 & n78365;
  assign n78367 = n78220 & n78224;
  assign n78368 = ~n78364 & ~n78366;
  assign n78369 = ~n78367 & n78368;
  assign n78370 = P3_DATAO_REG_5_ & n77726;
  assign n78371 = n78369 & n78370;
  assign n78372 = ~n78369 & ~n78370;
  assign n78373 = P3_DATAO_REG_5_ & n78036;
  assign n78374 = ~n78140 & n78213;
  assign n78375 = ~n78214 & ~n78374;
  assign n78376 = n78147 & ~n78375;
  assign n78377 = ~n78140 & ~n78213;
  assign n78378 = ~n78147 & n78377;
  assign n78379 = n78148 & n78213;
  assign n78380 = ~n78376 & ~n78378;
  assign n78381 = ~n78379 & n78380;
  assign n78382 = P3_DATAO_REG_5_ & n77955;
  assign n78383 = n78381 & n78382;
  assign n78384 = ~n78381 & ~n78382;
  assign n78385 = P3_DATAO_REG_5_ & n77688;
  assign n78386 = ~n78160 & n78207;
  assign n78387 = ~n78208 & ~n78386;
  assign n78388 = n78167 & ~n78387;
  assign n78389 = ~n78160 & ~n78207;
  assign n78390 = ~n78167 & n78389;
  assign n78391 = n78168 & n78207;
  assign n78392 = ~n78388 & ~n78390;
  assign n78393 = ~n78391 & n78392;
  assign n78394 = P3_DATAO_REG_5_ & n77434;
  assign n78395 = n78393 & n78394;
  assign n78396 = ~n78393 & ~n78394;
  assign n78397 = P3_DATAO_REG_5_ & n77436;
  assign n78398 = P3_DATAO_REG_5_ & n77475;
  assign n78399 = P3_DATAO_REG_5_ & n77438;
  assign n78400 = n78192 & ~n78199;
  assign n78401 = ~n78192 & n78199;
  assign n78402 = ~n78400 & ~n78401;
  assign n78403 = ~n78191 & n78402;
  assign n78404 = n78191 & n78401;
  assign n78405 = n78193 & ~n78199;
  assign n78406 = ~n78403 & ~n78404;
  assign n78407 = ~n78405 & n78406;
  assign n78408 = n78399 & ~n78407;
  assign n78409 = ~n77629 & ~n77638;
  assign n78410 = ~n77634 & ~n78409;
  assign n78411 = ~n77642 & ~n78410;
  assign n78412 = n78399 & ~n78411;
  assign n78413 = ~n78407 & ~n78411;
  assign n78414 = ~n78408 & ~n78412;
  assign n78415 = ~n78413 & n78414;
  assign n78416 = n78398 & ~n78415;
  assign n78417 = ~n78180 & n78188;
  assign n78418 = ~n78189 & ~n78417;
  assign n78419 = n78201 & ~n78418;
  assign n78420 = ~n78180 & ~n78188;
  assign n78421 = ~n78201 & n78420;
  assign n78422 = n78188 & n78202;
  assign n78423 = ~n78419 & ~n78421;
  assign n78424 = ~n78422 & n78423;
  assign n78425 = ~n78398 & n78415;
  assign n78426 = n78424 & ~n78425;
  assign n78427 = ~n78416 & ~n78426;
  assign n78428 = n78397 & ~n78427;
  assign n78429 = ~n78176 & n78177;
  assign n78430 = n78176 & ~n78177;
  assign n78431 = ~n78429 & ~n78430;
  assign n78432 = n78205 & ~n78431;
  assign n78433 = ~n78178 & ~n78179;
  assign n78434 = ~n78205 & ~n78433;
  assign n78435 = ~n78432 & ~n78434;
  assign n78436 = n78397 & ~n78435;
  assign n78437 = ~n78427 & ~n78435;
  assign n78438 = ~n78428 & ~n78436;
  assign n78439 = ~n78437 & n78438;
  assign n78440 = ~n78396 & ~n78439;
  assign n78441 = ~n78395 & ~n78440;
  assign n78442 = n78385 & ~n78441;
  assign n78443 = ~n78156 & n78157;
  assign n78444 = n78156 & ~n78157;
  assign n78445 = ~n78443 & ~n78444;
  assign n78446 = n78211 & ~n78445;
  assign n78447 = ~n78158 & ~n78159;
  assign n78448 = ~n78211 & ~n78447;
  assign n78449 = ~n78446 & ~n78448;
  assign n78450 = n78385 & ~n78449;
  assign n78451 = ~n78441 & ~n78449;
  assign n78452 = ~n78442 & ~n78450;
  assign n78453 = ~n78451 & n78452;
  assign n78454 = ~n78384 & ~n78453;
  assign n78455 = ~n78383 & ~n78454;
  assign n78456 = n78373 & ~n78455;
  assign n78457 = ~n78136 & n78137;
  assign n78458 = n78136 & ~n78137;
  assign n78459 = ~n78457 & ~n78458;
  assign n78460 = n78217 & ~n78459;
  assign n78461 = ~n78138 & ~n78139;
  assign n78462 = ~n78217 & ~n78461;
  assign n78463 = ~n78460 & ~n78462;
  assign n78464 = n78373 & ~n78463;
  assign n78465 = ~n78455 & ~n78463;
  assign n78466 = ~n78456 & ~n78464;
  assign n78467 = ~n78465 & n78466;
  assign n78468 = ~n78372 & ~n78467;
  assign n78469 = ~n78371 & ~n78468;
  assign n78470 = n78361 & ~n78469;
  assign n78471 = ~n78126 & ~n78127;
  assign n78472 = n78228 & n78471;
  assign n78473 = ~n78228 & ~n78471;
  assign n78474 = ~n78472 & ~n78473;
  assign n78475 = n78361 & ~n78474;
  assign n78476 = ~n78469 & ~n78474;
  assign n78477 = ~n78470 & ~n78475;
  assign n78478 = ~n78476 & n78477;
  assign n78479 = ~n78360 & ~n78478;
  assign n78480 = ~n78359 & ~n78479;
  assign n78481 = n77721 & ~n78480;
  assign n78482 = ~n77721 & n78480;
  assign n78483 = ~n78481 & ~n78482;
  assign n78484 = P3_DATAO_REG_6_ & n77722;
  assign n78485 = n77725 & ~n78355;
  assign n78486 = ~n77725 & n78355;
  assign n78487 = ~n78230 & ~n78486;
  assign n78488 = ~n78485 & ~n78487;
  assign n78489 = n78484 & ~n78488;
  assign n78490 = ~n78484 & n78488;
  assign n78491 = ~n78237 & n78238;
  assign n78492 = ~n78237 & n78346;
  assign n78493 = ~n78351 & ~n78491;
  assign n78494 = ~n78492 & n78493;
  assign n78495 = P3_DATAO_REG_7_ & n77724;
  assign n78496 = ~n78240 & n78336;
  assign n78497 = ~n78337 & ~n78343;
  assign n78498 = ~n78496 & n78497;
  assign n78499 = n77726 & ~n78498;
  assign n78500 = ~n77726 & n78498;
  assign n78501 = P3_DATAO_REG_8_ & ~n78499;
  assign n78502 = ~n78500 & n78501;
  assign n78503 = ~n78242 & ~n78333;
  assign n78504 = ~n78251 & ~n78323;
  assign n78505 = ~n78324 & ~n78330;
  assign n78506 = ~n78504 & n78505;
  assign n78507 = P3_DATAO_REG_10_ & n77955;
  assign n78508 = ~n78259 & ~n78304;
  assign n78509 = ~n78305 & ~n78311;
  assign n78510 = ~n78508 & n78509;
  assign n78511 = P3_DATAO_REG_12_ & n77434;
  assign n78512 = ~n78264 & ~n78301;
  assign n78513 = ~n78300 & ~n78512;
  assign n78514 = P3_DATAO_REG_13_ & n77436;
  assign n78515 = P3_DATAO_REG_15_ & n77438;
  assign n78516 = ~n78273 & ~n78281;
  assign n78517 = ~n78282 & ~n78516;
  assign n78518 = n78515 & ~n78517;
  assign n78519 = ~n78515 & n78517;
  assign n78520 = ~n78518 & ~n78519;
  assign n78521 = P3_DATAO_REG_16_ & n77440;
  assign n78522 = P3_DATAO_REG_17_ & n77442;
  assign n78523 = P3_DATAO_REG_18_ & n77444;
  assign n78524 = n78522 & ~n78523;
  assign n78525 = ~n78522 & n78523;
  assign n78526 = ~n78524 & ~n78525;
  assign n78527 = n78521 & ~n78526;
  assign n78528 = ~n78521 & n78526;
  assign n78529 = P3_DATAO_REG_16_ & P3_DATAO_REG_17_;
  assign n78530 = n77451 & n78529;
  assign n78531 = ~n78527 & ~n78528;
  assign n78532 = ~n78530 & n78531;
  assign n78533 = ~n78521 & ~n78524;
  assign n78534 = ~n78527 & ~n78533;
  assign n78535 = n78530 & ~n78534;
  assign n78536 = ~n78532 & ~n78535;
  assign n78537 = ~n78520 & n78536;
  assign n78538 = n78520 & ~n78536;
  assign n78539 = ~n78537 & ~n78538;
  assign n78540 = P3_DATAO_REG_14_ & n77475;
  assign n78541 = ~n78539 & ~n78540;
  assign n78542 = n78539 & n78540;
  assign n78543 = ~n78267 & ~n78285;
  assign n78544 = ~n78286 & ~n78292;
  assign n78545 = ~n78543 & n78544;
  assign n78546 = ~n78541 & ~n78542;
  assign n78547 = n78545 & n78546;
  assign n78548 = ~n78545 & ~n78546;
  assign n78549 = ~n78547 & ~n78548;
  assign n78550 = n78514 & ~n78549;
  assign n78551 = ~n78514 & n78549;
  assign n78552 = ~n78550 & ~n78551;
  assign n78553 = n78513 & ~n78552;
  assign n78554 = ~n78514 & ~n78549;
  assign n78555 = ~n78513 & n78554;
  assign n78556 = ~n78513 & n78514;
  assign n78557 = n78549 & n78556;
  assign n78558 = ~n78553 & ~n78555;
  assign n78559 = ~n78557 & n78558;
  assign n78560 = n78511 & ~n78559;
  assign n78561 = ~n78511 & n78559;
  assign n78562 = ~n78560 & ~n78561;
  assign n78563 = n78510 & ~n78562;
  assign n78564 = n78511 & n78559;
  assign n78565 = ~n78511 & ~n78559;
  assign n78566 = ~n78564 & ~n78565;
  assign n78567 = ~n78510 & ~n78566;
  assign n78568 = ~n78563 & ~n78567;
  assign n78569 = P3_DATAO_REG_11_ & n77688;
  assign n78570 = ~n78256 & ~n78320;
  assign n78571 = ~n78319 & ~n78570;
  assign n78572 = ~n78568 & ~n78569;
  assign n78573 = ~n78571 & n78572;
  assign n78574 = ~n78568 & n78569;
  assign n78575 = n78568 & ~n78569;
  assign n78576 = ~n78574 & ~n78575;
  assign n78577 = n78571 & ~n78576;
  assign n78578 = ~n78573 & ~n78577;
  assign n78579 = n78569 & ~n78571;
  assign n78580 = n78568 & n78579;
  assign n78581 = n78578 & ~n78580;
  assign n78582 = n78507 & ~n78581;
  assign n78583 = ~n78507 & n78581;
  assign n78584 = ~n78582 & ~n78583;
  assign n78585 = n78506 & ~n78584;
  assign n78586 = n78507 & n78581;
  assign n78587 = ~n78507 & ~n78581;
  assign n78588 = ~n78586 & ~n78587;
  assign n78589 = ~n78506 & ~n78588;
  assign n78590 = ~n78585 & ~n78589;
  assign n78591 = P3_DATAO_REG_9_ & n78036;
  assign n78592 = n78590 & ~n78591;
  assign n78593 = n78246 & ~n78333;
  assign n78594 = ~n78248 & ~n78593;
  assign n78595 = ~n78503 & ~n78592;
  assign n78596 = n78594 & n78595;
  assign n78597 = ~n78590 & n78591;
  assign n78598 = n78596 & ~n78597;
  assign n78599 = ~n78590 & ~n78591;
  assign n78600 = n78590 & n78591;
  assign n78601 = n78242 & n78333;
  assign n78602 = ~n78246 & ~n78503;
  assign n78603 = ~n78601 & ~n78602;
  assign n78604 = ~n78599 & ~n78600;
  assign n78605 = n78603 & n78604;
  assign n78606 = ~n78598 & ~n78605;
  assign n78607 = n78502 & ~n78606;
  assign n78608 = ~n78502 & n78606;
  assign n78609 = ~n78607 & ~n78608;
  assign n78610 = n78495 & ~n78609;
  assign n78611 = ~n78495 & n78609;
  assign n78612 = ~n78610 & ~n78611;
  assign n78613 = n78494 & ~n78612;
  assign n78614 = ~n78495 & ~n78609;
  assign n78615 = ~n78494 & n78614;
  assign n78616 = ~n78494 & n78495;
  assign n78617 = n78609 & n78616;
  assign n78618 = ~n78613 & ~n78615;
  assign n78619 = ~n78617 & n78618;
  assign n78620 = ~n78489 & ~n78490;
  assign n78621 = ~n78619 & n78620;
  assign n78622 = n78619 & ~n78620;
  assign n78623 = ~n78621 & ~n78622;
  assign n78624 = ~n78483 & n78623;
  assign n78625 = n78483 & ~n78623;
  assign n78626 = ~n78624 & ~n78625;
  assign n78627 = n77719 & n78626;
  assign n78628 = ~n77719 & ~n78626;
  assign n78629 = P3_DATAO_REG_4_ & n77720;
  assign n78630 = P3_DATAO_REG_4_ & n77722;
  assign n78631 = P3_DATAO_REG_4_ & n77724;
  assign n78632 = ~n78369 & n78370;
  assign n78633 = n78369 & ~n78370;
  assign n78634 = ~n78632 & ~n78633;
  assign n78635 = n78467 & ~n78634;
  assign n78636 = ~n78371 & ~n78372;
  assign n78637 = ~n78467 & ~n78636;
  assign n78638 = ~n78635 & ~n78637;
  assign n78639 = n78631 & ~n78638;
  assign n78640 = ~n78373 & n78463;
  assign n78641 = ~n78464 & ~n78640;
  assign n78642 = n78455 & ~n78641;
  assign n78643 = ~n78373 & ~n78463;
  assign n78644 = ~n78455 & n78643;
  assign n78645 = n78456 & n78463;
  assign n78646 = ~n78642 & ~n78644;
  assign n78647 = ~n78645 & n78646;
  assign n78648 = P3_DATAO_REG_4_ & n77726;
  assign n78649 = n78647 & n78648;
  assign n78650 = ~n78647 & ~n78648;
  assign n78651 = P3_DATAO_REG_4_ & n78036;
  assign n78652 = ~n78385 & n78449;
  assign n78653 = ~n78450 & ~n78652;
  assign n78654 = n78441 & ~n78653;
  assign n78655 = ~n78385 & ~n78449;
  assign n78656 = ~n78441 & n78655;
  assign n78657 = n78442 & n78449;
  assign n78658 = ~n78654 & ~n78656;
  assign n78659 = ~n78657 & n78658;
  assign n78660 = P3_DATAO_REG_4_ & n77955;
  assign n78661 = n78659 & n78660;
  assign n78662 = ~n78659 & ~n78660;
  assign n78663 = P3_DATAO_REG_4_ & n77688;
  assign n78664 = ~n78397 & n78435;
  assign n78665 = ~n78436 & ~n78664;
  assign n78666 = n78427 & ~n78665;
  assign n78667 = ~n78397 & ~n78435;
  assign n78668 = ~n78427 & n78667;
  assign n78669 = n78428 & n78435;
  assign n78670 = ~n78666 & ~n78668;
  assign n78671 = ~n78669 & n78670;
  assign n78672 = P3_DATAO_REG_4_ & n77434;
  assign n78673 = n78671 & n78672;
  assign n78674 = ~n78671 & ~n78672;
  assign n78675 = P3_DATAO_REG_4_ & n77436;
  assign n78676 = n78398 & ~n78424;
  assign n78677 = ~n78398 & n78424;
  assign n78678 = ~n78676 & ~n78677;
  assign n78679 = n78415 & ~n78678;
  assign n78680 = ~n78398 & ~n78424;
  assign n78681 = ~n78415 & n78680;
  assign n78682 = n78416 & n78424;
  assign n78683 = ~n78679 & ~n78681;
  assign n78684 = ~n78682 & n78683;
  assign n78685 = n78675 & ~n78684;
  assign n78686 = P3_DATAO_REG_4_ & n77475;
  assign n78687 = ~n77627 & ~n77645;
  assign n78688 = ~n77646 & ~n77652;
  assign n78689 = ~n78687 & n78688;
  assign n78690 = n78686 & ~n78689;
  assign n78691 = ~n78399 & n78407;
  assign n78692 = ~n78408 & ~n78691;
  assign n78693 = n78411 & ~n78692;
  assign n78694 = ~n78399 & ~n78407;
  assign n78695 = ~n78411 & n78694;
  assign n78696 = n78407 & n78412;
  assign n78697 = ~n78693 & ~n78695;
  assign n78698 = ~n78696 & n78697;
  assign n78699 = ~n78686 & n78689;
  assign n78700 = n78698 & ~n78699;
  assign n78701 = ~n78690 & ~n78700;
  assign n78702 = n78675 & ~n78701;
  assign n78703 = ~n78684 & ~n78701;
  assign n78704 = ~n78685 & ~n78702;
  assign n78705 = ~n78703 & n78704;
  assign n78706 = ~n78674 & ~n78705;
  assign n78707 = ~n78673 & ~n78706;
  assign n78708 = n78663 & ~n78707;
  assign n78709 = ~n78393 & n78394;
  assign n78710 = n78393 & ~n78394;
  assign n78711 = ~n78709 & ~n78710;
  assign n78712 = n78439 & ~n78711;
  assign n78713 = ~n78395 & ~n78396;
  assign n78714 = ~n78439 & ~n78713;
  assign n78715 = ~n78712 & ~n78714;
  assign n78716 = n78663 & ~n78715;
  assign n78717 = ~n78707 & ~n78715;
  assign n78718 = ~n78708 & ~n78716;
  assign n78719 = ~n78717 & n78718;
  assign n78720 = ~n78662 & ~n78719;
  assign n78721 = ~n78661 & ~n78720;
  assign n78722 = n78651 & ~n78721;
  assign n78723 = ~n78381 & n78382;
  assign n78724 = n78381 & ~n78382;
  assign n78725 = ~n78723 & ~n78724;
  assign n78726 = n78453 & ~n78725;
  assign n78727 = ~n78383 & ~n78384;
  assign n78728 = ~n78453 & ~n78727;
  assign n78729 = ~n78726 & ~n78728;
  assign n78730 = n78651 & ~n78729;
  assign n78731 = ~n78721 & ~n78729;
  assign n78732 = ~n78722 & ~n78730;
  assign n78733 = ~n78731 & n78732;
  assign n78734 = ~n78650 & ~n78733;
  assign n78735 = ~n78649 & ~n78734;
  assign n78736 = n78631 & ~n78735;
  assign n78737 = ~n78638 & ~n78735;
  assign n78738 = ~n78639 & ~n78736;
  assign n78739 = ~n78737 & n78738;
  assign n78740 = n78630 & ~n78739;
  assign n78741 = ~n78361 & n78474;
  assign n78742 = ~n78475 & ~n78741;
  assign n78743 = n78469 & ~n78742;
  assign n78744 = ~n78361 & ~n78474;
  assign n78745 = ~n78469 & n78744;
  assign n78746 = n78470 & n78474;
  assign n78747 = ~n78743 & ~n78745;
  assign n78748 = ~n78746 & n78747;
  assign n78749 = ~n78630 & n78739;
  assign n78750 = n78748 & ~n78749;
  assign n78751 = ~n78740 & ~n78750;
  assign n78752 = n78629 & ~n78751;
  assign n78753 = ~n78359 & ~n78360;
  assign n78754 = n78478 & n78753;
  assign n78755 = ~n78478 & ~n78753;
  assign n78756 = ~n78754 & ~n78755;
  assign n78757 = n78629 & ~n78756;
  assign n78758 = ~n78751 & ~n78756;
  assign n78759 = ~n78752 & ~n78757;
  assign n78760 = ~n78758 & n78759;
  assign n78761 = ~n78628 & ~n78760;
  assign n78762 = ~n78627 & ~n78761;
  assign n78763 = n77717 & ~n78762;
  assign n78764 = ~n77717 & n78762;
  assign n78765 = ~n78763 & ~n78764;
  assign n78766 = n77721 & ~n78623;
  assign n78767 = ~n77721 & n78623;
  assign n78768 = ~n78480 & ~n78767;
  assign n78769 = ~n78766 & ~n78768;
  assign n78770 = P3_DATAO_REG_5_ & n77718;
  assign n78771 = ~n78490 & n78619;
  assign n78772 = ~n78489 & ~n78771;
  assign n78773 = P3_DATAO_REG_6_ & n77720;
  assign n78774 = ~n78494 & ~n78609;
  assign n78775 = ~n78610 & ~n78616;
  assign n78776 = ~n78774 & n78775;
  assign n78777 = P3_DATAO_REG_7_ & n77722;
  assign n78778 = P3_DATAO_REG_8_ & ~n78500;
  assign n78779 = n78606 & n78778;
  assign n78780 = ~n78499 & ~n78779;
  assign n78781 = P3_DATAO_REG_8_ & n77724;
  assign n78782 = P3_DATAO_REG_10_ & n78036;
  assign n78783 = ~n78506 & ~n78587;
  assign n78784 = ~n78586 & ~n78783;
  assign n78785 = n78782 & ~n78784;
  assign n78786 = ~n78782 & n78784;
  assign n78787 = ~n78785 & ~n78786;
  assign n78788 = P3_DATAO_REG_11_ & n77955;
  assign n78789 = ~n78568 & ~n78571;
  assign n78790 = ~n78574 & ~n78579;
  assign n78791 = ~n78789 & n78790;
  assign n78792 = n78788 & ~n78791;
  assign n78793 = ~n78788 & n78791;
  assign n78794 = ~n78792 & ~n78793;
  assign n78795 = ~n78510 & ~n78565;
  assign n78796 = ~n78564 & ~n78795;
  assign n78797 = P3_DATAO_REG_12_ & n77688;
  assign n78798 = ~n78513 & ~n78549;
  assign n78799 = ~n78550 & ~n78556;
  assign n78800 = ~n78798 & n78799;
  assign n78801 = P3_DATAO_REG_13_ & n77434;
  assign n78802 = n78515 & ~n78536;
  assign n78803 = ~n78515 & n78536;
  assign n78804 = ~n78517 & ~n78803;
  assign n78805 = ~n78802 & ~n78804;
  assign n78806 = P3_DATAO_REG_15_ & n77475;
  assign n78807 = P3_DATAO_REG_17_ & n77440;
  assign n78808 = P3_DATAO_REG_18_ & n77442;
  assign n78809 = P3_DATAO_REG_19_ & n77444;
  assign n78810 = n78808 & ~n78809;
  assign n78811 = ~n78808 & n78809;
  assign n78812 = ~n78810 & ~n78811;
  assign n78813 = n78807 & ~n78812;
  assign n78814 = ~n78807 & n78812;
  assign n78815 = P3_DATAO_REG_17_ & P3_DATAO_REG_18_;
  assign n78816 = n77451 & n78815;
  assign n78817 = ~n78813 & ~n78814;
  assign n78818 = ~n78816 & n78817;
  assign n78819 = n78807 & ~n78810;
  assign n78820 = ~n78807 & n78810;
  assign n78821 = ~n78819 & ~n78820;
  assign n78822 = n78816 & n78821;
  assign n78823 = ~n78818 & ~n78822;
  assign n78824 = P3_DATAO_REG_16_ & n77438;
  assign n78825 = ~n78528 & n78530;
  assign n78826 = ~n78527 & ~n78825;
  assign n78827 = ~n78823 & ~n78824;
  assign n78828 = ~n78826 & n78827;
  assign n78829 = n78823 & n78824;
  assign n78830 = ~n78827 & ~n78829;
  assign n78831 = n78826 & n78830;
  assign n78832 = ~n78828 & ~n78831;
  assign n78833 = n78824 & ~n78826;
  assign n78834 = n78823 & n78833;
  assign n78835 = n78832 & ~n78834;
  assign n78836 = n78806 & ~n78835;
  assign n78837 = ~n78806 & n78835;
  assign n78838 = ~n78836 & ~n78837;
  assign n78839 = n78805 & ~n78838;
  assign n78840 = n78806 & n78832;
  assign n78841 = ~n78834 & n78840;
  assign n78842 = ~n78806 & ~n78835;
  assign n78843 = ~n78841 & ~n78842;
  assign n78844 = ~n78805 & ~n78843;
  assign n78845 = ~n78839 & ~n78844;
  assign n78846 = P3_DATAO_REG_14_ & n77436;
  assign n78847 = ~n78541 & ~n78545;
  assign n78848 = ~n78542 & ~n78847;
  assign n78849 = ~n78845 & ~n78846;
  assign n78850 = ~n78848 & n78849;
  assign n78851 = ~n78845 & n78846;
  assign n78852 = n78845 & ~n78846;
  assign n78853 = ~n78851 & ~n78852;
  assign n78854 = n78848 & ~n78853;
  assign n78855 = ~n78850 & ~n78854;
  assign n78856 = n78846 & ~n78848;
  assign n78857 = n78845 & n78856;
  assign n78858 = n78855 & ~n78857;
  assign n78859 = n78801 & ~n78858;
  assign n78860 = ~n78801 & n78858;
  assign n78861 = ~n78859 & ~n78860;
  assign n78862 = n78800 & ~n78861;
  assign n78863 = n78801 & ~n78857;
  assign n78864 = n78855 & n78863;
  assign n78865 = ~n78801 & ~n78858;
  assign n78866 = ~n78864 & ~n78865;
  assign n78867 = ~n78800 & ~n78866;
  assign n78868 = ~n78862 & ~n78867;
  assign n78869 = n78797 & ~n78868;
  assign n78870 = ~n78797 & n78868;
  assign n78871 = ~n78869 & ~n78870;
  assign n78872 = n78796 & ~n78871;
  assign n78873 = ~n78797 & ~n78868;
  assign n78874 = ~n78796 & n78873;
  assign n78875 = ~n78796 & n78797;
  assign n78876 = n78868 & n78875;
  assign n78877 = ~n78872 & ~n78874;
  assign n78878 = ~n78876 & n78877;
  assign n78879 = n78794 & ~n78878;
  assign n78880 = ~n78794 & n78878;
  assign n78881 = ~n78879 & ~n78880;
  assign n78882 = ~n78787 & n78881;
  assign n78883 = n78787 & ~n78881;
  assign n78884 = ~n78882 & ~n78883;
  assign n78885 = P3_DATAO_REG_9_ & n77726;
  assign n78886 = n78884 & n78885;
  assign n78887 = ~n78884 & ~n78885;
  assign n78888 = ~n78886 & ~n78887;
  assign n78889 = ~n78596 & ~n78597;
  assign n78890 = ~n78888 & ~n78889;
  assign n78891 = n78888 & n78889;
  assign n78892 = ~n78890 & ~n78891;
  assign n78893 = n78781 & ~n78892;
  assign n78894 = ~n78781 & n78892;
  assign n78895 = ~n78893 & ~n78894;
  assign n78896 = n78780 & ~n78895;
  assign n78897 = ~n78781 & ~n78892;
  assign n78898 = ~n78780 & n78897;
  assign n78899 = ~n78780 & n78781;
  assign n78900 = n78892 & n78899;
  assign n78901 = ~n78896 & ~n78898;
  assign n78902 = ~n78900 & n78901;
  assign n78903 = n78777 & ~n78902;
  assign n78904 = ~n78777 & n78902;
  assign n78905 = ~n78903 & ~n78904;
  assign n78906 = n78776 & ~n78905;
  assign n78907 = n78777 & n78902;
  assign n78908 = ~n78777 & ~n78902;
  assign n78909 = ~n78907 & ~n78908;
  assign n78910 = ~n78776 & ~n78909;
  assign n78911 = ~n78906 & ~n78910;
  assign n78912 = n78773 & ~n78911;
  assign n78913 = ~n78773 & n78911;
  assign n78914 = ~n78912 & ~n78913;
  assign n78915 = n78772 & ~n78914;
  assign n78916 = ~n78773 & ~n78911;
  assign n78917 = ~n78772 & n78916;
  assign n78918 = ~n78772 & n78773;
  assign n78919 = n78911 & n78918;
  assign n78920 = ~n78915 & ~n78917;
  assign n78921 = ~n78919 & n78920;
  assign n78922 = n78770 & ~n78921;
  assign n78923 = ~n78770 & n78921;
  assign n78924 = ~n78922 & ~n78923;
  assign n78925 = n78769 & ~n78924;
  assign n78926 = n78770 & n78921;
  assign n78927 = ~n78770 & ~n78921;
  assign n78928 = ~n78926 & ~n78927;
  assign n78929 = ~n78769 & ~n78928;
  assign n78930 = ~n78925 & ~n78929;
  assign n78931 = ~n78765 & n78930;
  assign n78932 = n78765 & ~n78930;
  assign n78933 = ~n78931 & ~n78932;
  assign n78934 = ~SEL & DIN_16_;
  assign n78935 = P3_DATAO_REG_3_ & n78934;
  assign n78936 = ~n78933 & ~n78935;
  assign n78937 = n78933 & n78935;
  assign n78938 = P3_DATAO_REG_3_ & n77716;
  assign n78939 = ~n78627 & ~n78628;
  assign n78940 = ~n78760 & ~n78939;
  assign n78941 = n78760 & n78939;
  assign n78942 = ~n78940 & ~n78941;
  assign n78943 = n78938 & ~n78942;
  assign n78944 = ~n78938 & n78942;
  assign n78945 = ~n78629 & n78756;
  assign n78946 = ~n78757 & ~n78945;
  assign n78947 = n78751 & ~n78946;
  assign n78948 = ~n78629 & ~n78756;
  assign n78949 = ~n78751 & n78948;
  assign n78950 = n78752 & n78756;
  assign n78951 = ~n78947 & ~n78949;
  assign n78952 = ~n78950 & n78951;
  assign n78953 = P3_DATAO_REG_3_ & n77718;
  assign n78954 = n78952 & n78953;
  assign n78955 = ~n78952 & ~n78953;
  assign n78956 = P3_DATAO_REG_3_ & n77720;
  assign n78957 = ~n78631 & n78735;
  assign n78958 = ~n78736 & ~n78957;
  assign n78959 = n78638 & ~n78958;
  assign n78960 = ~n78631 & ~n78735;
  assign n78961 = ~n78638 & n78960;
  assign n78962 = n78639 & n78735;
  assign n78963 = ~n78959 & ~n78961;
  assign n78964 = ~n78962 & n78963;
  assign n78965 = P3_DATAO_REG_3_ & n77722;
  assign n78966 = n78964 & n78965;
  assign n78967 = ~n78964 & ~n78965;
  assign n78968 = P3_DATAO_REG_3_ & n77724;
  assign n78969 = ~n78651 & n78729;
  assign n78970 = ~n78730 & ~n78969;
  assign n78971 = n78721 & ~n78970;
  assign n78972 = ~n78651 & ~n78729;
  assign n78973 = ~n78721 & n78972;
  assign n78974 = n78722 & n78729;
  assign n78975 = ~n78971 & ~n78973;
  assign n78976 = ~n78974 & n78975;
  assign n78977 = P3_DATAO_REG_3_ & n77726;
  assign n78978 = n78976 & n78977;
  assign n78979 = ~n78976 & ~n78977;
  assign n78980 = P3_DATAO_REG_3_ & n78036;
  assign n78981 = ~n78663 & n78715;
  assign n78982 = ~n78716 & ~n78981;
  assign n78983 = n78707 & ~n78982;
  assign n78984 = ~n78663 & ~n78715;
  assign n78985 = ~n78707 & n78984;
  assign n78986 = n78708 & n78715;
  assign n78987 = ~n78983 & ~n78985;
  assign n78988 = ~n78986 & n78987;
  assign n78989 = P3_DATAO_REG_3_ & n77955;
  assign n78990 = n78988 & n78989;
  assign n78991 = ~n78988 & ~n78989;
  assign n78992 = P3_DATAO_REG_3_ & n77688;
  assign n78993 = P3_DATAO_REG_3_ & n77434;
  assign n78994 = P3_DATAO_REG_3_ & n77436;
  assign n78995 = n78686 & ~n78698;
  assign n78996 = ~n78686 & n78698;
  assign n78997 = ~n78995 & ~n78996;
  assign n78998 = n78689 & ~n78997;
  assign n78999 = ~n78686 & ~n78698;
  assign n79000 = ~n78689 & n78999;
  assign n79001 = n78690 & n78698;
  assign n79002 = ~n78998 & ~n79000;
  assign n79003 = ~n79001 & n79002;
  assign n79004 = n78994 & ~n79003;
  assign n79005 = ~n77624 & n77661;
  assign n79006 = n77655 & ~n79005;
  assign n79007 = ~n77665 & ~n79006;
  assign n79008 = n78994 & ~n79007;
  assign n79009 = ~n79003 & ~n79007;
  assign n79010 = ~n79004 & ~n79008;
  assign n79011 = ~n79009 & n79010;
  assign n79012 = n78993 & ~n79011;
  assign n79013 = ~n78675 & n78684;
  assign n79014 = ~n78685 & ~n79013;
  assign n79015 = n78701 & ~n79014;
  assign n79016 = ~n78675 & ~n78684;
  assign n79017 = ~n78701 & n79016;
  assign n79018 = n78684 & n78702;
  assign n79019 = ~n79015 & ~n79017;
  assign n79020 = ~n79018 & n79019;
  assign n79021 = ~n78993 & n79011;
  assign n79022 = n79020 & ~n79021;
  assign n79023 = ~n79012 & ~n79022;
  assign n79024 = n78992 & ~n79023;
  assign n79025 = ~n78671 & n78672;
  assign n79026 = n78671 & ~n78672;
  assign n79027 = ~n79025 & ~n79026;
  assign n79028 = n78705 & ~n79027;
  assign n79029 = ~n78673 & ~n78674;
  assign n79030 = ~n78705 & ~n79029;
  assign n79031 = ~n79028 & ~n79030;
  assign n79032 = n78992 & ~n79031;
  assign n79033 = ~n79023 & ~n79031;
  assign n79034 = ~n79024 & ~n79032;
  assign n79035 = ~n79033 & n79034;
  assign n79036 = ~n78991 & ~n79035;
  assign n79037 = ~n78990 & ~n79036;
  assign n79038 = n78980 & ~n79037;
  assign n79039 = ~n78659 & n78660;
  assign n79040 = n78659 & ~n78660;
  assign n79041 = ~n79039 & ~n79040;
  assign n79042 = n78719 & ~n79041;
  assign n79043 = ~n78661 & ~n78662;
  assign n79044 = ~n78719 & ~n79043;
  assign n79045 = ~n79042 & ~n79044;
  assign n79046 = n78980 & ~n79045;
  assign n79047 = ~n79037 & ~n79045;
  assign n79048 = ~n79038 & ~n79046;
  assign n79049 = ~n79047 & n79048;
  assign n79050 = ~n78979 & ~n79049;
  assign n79051 = ~n78978 & ~n79050;
  assign n79052 = n78968 & ~n79051;
  assign n79053 = ~n78647 & n78648;
  assign n79054 = n78647 & ~n78648;
  assign n79055 = ~n79053 & ~n79054;
  assign n79056 = n78733 & ~n79055;
  assign n79057 = ~n78649 & ~n78650;
  assign n79058 = ~n78733 & ~n79057;
  assign n79059 = ~n79056 & ~n79058;
  assign n79060 = n78968 & ~n79059;
  assign n79061 = ~n79051 & ~n79059;
  assign n79062 = ~n79052 & ~n79060;
  assign n79063 = ~n79061 & n79062;
  assign n79064 = ~n78967 & ~n79063;
  assign n79065 = ~n78966 & ~n79064;
  assign n79066 = n78956 & ~n79065;
  assign n79067 = ~n78740 & ~n78749;
  assign n79068 = ~n78748 & n79067;
  assign n79069 = n78748 & ~n79067;
  assign n79070 = ~n79068 & ~n79069;
  assign n79071 = n78956 & ~n79070;
  assign n79072 = ~n79065 & ~n79070;
  assign n79073 = ~n79066 & ~n79071;
  assign n79074 = ~n79072 & n79073;
  assign n79075 = ~n78955 & ~n79074;
  assign n79076 = ~n78954 & ~n79075;
  assign n79077 = ~n78944 & ~n79076;
  assign n79078 = ~n78943 & ~n79077;
  assign n79079 = ~n78936 & ~n78937;
  assign n79080 = n79078 & n79079;
  assign n79081 = ~n79078 & ~n79079;
  assign n79082 = ~n79080 & ~n79081;
  assign n79083 = n77715 & ~n79082;
  assign n79084 = ~n77715 & n79082;
  assign n79085 = P3_DATAO_REG_2_ & n78934;
  assign n79086 = n78938 & n78942;
  assign n79087 = ~n78938 & ~n78942;
  assign n79088 = ~n79086 & ~n79087;
  assign n79089 = ~n79076 & ~n79088;
  assign n79090 = n79076 & n79088;
  assign n79091 = ~n79089 & ~n79090;
  assign n79092 = n79085 & n79091;
  assign n79093 = ~n79085 & ~n79091;
  assign n79094 = P3_DATAO_REG_2_ & n77716;
  assign n79095 = ~n78952 & n78953;
  assign n79096 = n78952 & ~n78953;
  assign n79097 = ~n79095 & ~n79096;
  assign n79098 = n79074 & ~n79097;
  assign n79099 = ~n78954 & ~n78955;
  assign n79100 = ~n79074 & ~n79099;
  assign n79101 = ~n79098 & ~n79100;
  assign n79102 = n79094 & ~n79101;
  assign n79103 = ~n78956 & n79070;
  assign n79104 = ~n79071 & ~n79103;
  assign n79105 = n79065 & ~n79104;
  assign n79106 = ~n78956 & ~n79070;
  assign n79107 = ~n79065 & n79106;
  assign n79108 = n79066 & n79070;
  assign n79109 = ~n79105 & ~n79107;
  assign n79110 = ~n79108 & n79109;
  assign n79111 = P3_DATAO_REG_2_ & n77718;
  assign n79112 = n79110 & n79111;
  assign n79113 = ~n79110 & ~n79111;
  assign n79114 = P3_DATAO_REG_2_ & n77720;
  assign n79115 = ~n78968 & n79059;
  assign n79116 = ~n79060 & ~n79115;
  assign n79117 = n79051 & ~n79116;
  assign n79118 = ~n78968 & ~n79059;
  assign n79119 = ~n79051 & n79118;
  assign n79120 = n79052 & n79059;
  assign n79121 = ~n79117 & ~n79119;
  assign n79122 = ~n79120 & n79121;
  assign n79123 = P3_DATAO_REG_2_ & n77722;
  assign n79124 = n79122 & n79123;
  assign n79125 = ~n79122 & ~n79123;
  assign n79126 = P3_DATAO_REG_2_ & n77724;
  assign n79127 = ~n78980 & n79045;
  assign n79128 = ~n79046 & ~n79127;
  assign n79129 = n79037 & ~n79128;
  assign n79130 = ~n78980 & ~n79045;
  assign n79131 = ~n79037 & n79130;
  assign n79132 = n79038 & n79045;
  assign n79133 = ~n79129 & ~n79131;
  assign n79134 = ~n79132 & n79133;
  assign n79135 = P3_DATAO_REG_2_ & n77726;
  assign n79136 = n79134 & n79135;
  assign n79137 = ~n79134 & ~n79135;
  assign n79138 = P3_DATAO_REG_2_ & n78036;
  assign n79139 = ~n78992 & n79031;
  assign n79140 = ~n79032 & ~n79139;
  assign n79141 = n79023 & ~n79140;
  assign n79142 = ~n78992 & ~n79031;
  assign n79143 = ~n79023 & n79142;
  assign n79144 = n79024 & n79031;
  assign n79145 = ~n79141 & ~n79143;
  assign n79146 = ~n79144 & n79145;
  assign n79147 = P3_DATAO_REG_2_ & n77955;
  assign n79148 = n79146 & n79147;
  assign n79149 = ~n79146 & ~n79147;
  assign n79150 = P3_DATAO_REG_2_ & n77688;
  assign n79151 = ~n78994 & n79003;
  assign n79152 = ~n79004 & ~n79151;
  assign n79153 = n79007 & ~n79152;
  assign n79154 = ~n78994 & ~n79003;
  assign n79155 = ~n79007 & n79154;
  assign n79156 = n79003 & n79008;
  assign n79157 = ~n79153 & ~n79155;
  assign n79158 = ~n79156 & n79157;
  assign n79159 = P3_DATAO_REG_2_ & n77434;
  assign n79160 = n79158 & n79159;
  assign n79161 = ~n79158 & ~n79159;
  assign n79162 = ~n77622 & ~n77668;
  assign n79163 = ~n77669 & ~n77675;
  assign n79164 = ~n79162 & n79163;
  assign n79165 = ~n79161 & ~n79164;
  assign n79166 = ~n79160 & ~n79165;
  assign n79167 = n79150 & ~n79166;
  assign n79168 = n78993 & ~n79020;
  assign n79169 = ~n78993 & n79020;
  assign n79170 = ~n79168 & ~n79169;
  assign n79171 = n79011 & ~n79170;
  assign n79172 = ~n78993 & ~n79020;
  assign n79173 = ~n79011 & n79172;
  assign n79174 = n79012 & n79020;
  assign n79175 = ~n79171 & ~n79173;
  assign n79176 = ~n79174 & n79175;
  assign n79177 = n79150 & ~n79176;
  assign n79178 = ~n79166 & ~n79176;
  assign n79179 = ~n79167 & ~n79177;
  assign n79180 = ~n79178 & n79179;
  assign n79181 = ~n79149 & ~n79180;
  assign n79182 = ~n79148 & ~n79181;
  assign n79183 = n79138 & ~n79182;
  assign n79184 = ~n78988 & n78989;
  assign n79185 = n78988 & ~n78989;
  assign n79186 = ~n79184 & ~n79185;
  assign n79187 = n79035 & ~n79186;
  assign n79188 = ~n78990 & ~n78991;
  assign n79189 = ~n79035 & ~n79188;
  assign n79190 = ~n79187 & ~n79189;
  assign n79191 = n79138 & ~n79190;
  assign n79192 = ~n79182 & ~n79190;
  assign n79193 = ~n79183 & ~n79191;
  assign n79194 = ~n79192 & n79193;
  assign n79195 = ~n79137 & ~n79194;
  assign n79196 = ~n79136 & ~n79195;
  assign n79197 = n79126 & ~n79196;
  assign n79198 = ~n78976 & n78977;
  assign n79199 = n78976 & ~n78977;
  assign n79200 = ~n79198 & ~n79199;
  assign n79201 = n79049 & ~n79200;
  assign n79202 = ~n78978 & ~n78979;
  assign n79203 = ~n79049 & ~n79202;
  assign n79204 = ~n79201 & ~n79203;
  assign n79205 = n79126 & ~n79204;
  assign n79206 = ~n79196 & ~n79204;
  assign n79207 = ~n79197 & ~n79205;
  assign n79208 = ~n79206 & n79207;
  assign n79209 = ~n79125 & ~n79208;
  assign n79210 = ~n79124 & ~n79209;
  assign n79211 = n79114 & ~n79210;
  assign n79212 = ~n78964 & n78965;
  assign n79213 = n78964 & ~n78965;
  assign n79214 = ~n79212 & ~n79213;
  assign n79215 = n79063 & ~n79214;
  assign n79216 = ~n78966 & ~n78967;
  assign n79217 = ~n79063 & ~n79216;
  assign n79218 = ~n79215 & ~n79217;
  assign n79219 = n79114 & ~n79218;
  assign n79220 = ~n79210 & ~n79218;
  assign n79221 = ~n79211 & ~n79219;
  assign n79222 = ~n79220 & n79221;
  assign n79223 = ~n79113 & ~n79222;
  assign n79224 = ~n79112 & ~n79223;
  assign n79225 = n79094 & ~n79224;
  assign n79226 = ~n79101 & ~n79224;
  assign n79227 = ~n79102 & ~n79225;
  assign n79228 = ~n79226 & n79227;
  assign n79229 = ~n79093 & ~n79228;
  assign n79230 = ~n79092 & ~n79229;
  assign n79231 = ~n79084 & ~n79230;
  assign n79232 = ~n79083 & ~n79231;
  assign n79233 = n77713 & ~n79232;
  assign n79234 = ~n77713 & n79232;
  assign n79235 = ~n79233 & ~n79234;
  assign n79236 = ~n78936 & ~n79078;
  assign n79237 = ~n78937 & ~n79236;
  assign n79238 = P3_DATAO_REG_3_ & n77714;
  assign n79239 = n77717 & ~n78930;
  assign n79240 = ~n77717 & n78930;
  assign n79241 = ~n78762 & ~n79240;
  assign n79242 = ~n79239 & ~n79241;
  assign n79243 = P3_DATAO_REG_4_ & n78934;
  assign n79244 = ~n78769 & ~n78927;
  assign n79245 = ~n78926 & ~n79244;
  assign n79246 = P3_DATAO_REG_5_ & n77716;
  assign n79247 = ~n78772 & ~n78911;
  assign n79248 = ~n78912 & ~n78918;
  assign n79249 = ~n79247 & n79248;
  assign n79250 = P3_DATAO_REG_6_ & n77718;
  assign n79251 = n78885 & ~n78889;
  assign n79252 = ~n78885 & n78889;
  assign n79253 = n78884 & ~n79252;
  assign n79254 = ~n79251 & ~n79253;
  assign n79255 = P3_DATAO_REG_9_ & n77724;
  assign n79256 = n78782 & ~n78881;
  assign n79257 = ~n78782 & n78881;
  assign n79258 = ~n78784 & ~n79257;
  assign n79259 = ~n79256 & ~n79258;
  assign n79260 = P3_DATAO_REG_10_ & n77726;
  assign n79261 = ~n78796 & ~n78868;
  assign n79262 = ~n78869 & ~n78875;
  assign n79263 = ~n79261 & n79262;
  assign n79264 = P3_DATAO_REG_12_ & n77955;
  assign n79265 = P3_DATAO_REG_14_ & n77434;
  assign n79266 = ~n78845 & ~n78848;
  assign n79267 = ~n78851 & ~n78856;
  assign n79268 = ~n79266 & n79267;
  assign n79269 = n79265 & ~n79268;
  assign n79270 = ~n79265 & n79268;
  assign n79271 = ~n79269 & ~n79270;
  assign n79272 = ~n78805 & ~n78842;
  assign n79273 = ~n78841 & ~n79272;
  assign n79274 = P3_DATAO_REG_15_ & n77436;
  assign n79275 = ~n78823 & n78824;
  assign n79276 = ~n78823 & ~n78826;
  assign n79277 = ~n78833 & ~n79275;
  assign n79278 = ~n79276 & n79277;
  assign n79279 = P3_DATAO_REG_16_ & n77475;
  assign n79280 = P3_DATAO_REG_18_ & n77440;
  assign n79281 = P3_DATAO_REG_19_ & n77442;
  assign n79282 = P3_DATAO_REG_20_ & n77444;
  assign n79283 = n79281 & ~n79282;
  assign n79284 = ~n79281 & n79282;
  assign n79285 = ~n79283 & ~n79284;
  assign n79286 = n79280 & ~n79285;
  assign n79287 = ~n79280 & n79285;
  assign n79288 = P3_DATAO_REG_18_ & P3_DATAO_REG_19_;
  assign n79289 = n77451 & n79288;
  assign n79290 = ~n79286 & ~n79287;
  assign n79291 = ~n79289 & n79290;
  assign n79292 = ~n79280 & ~n79283;
  assign n79293 = ~n79286 & ~n79292;
  assign n79294 = n79289 & ~n79293;
  assign n79295 = ~n79291 & ~n79294;
  assign n79296 = P3_DATAO_REG_17_ & n77438;
  assign n79297 = ~n78814 & n78816;
  assign n79298 = ~n78813 & ~n79297;
  assign n79299 = ~n79295 & ~n79296;
  assign n79300 = ~n79298 & n79299;
  assign n79301 = ~n79295 & n79296;
  assign n79302 = n79295 & ~n79296;
  assign n79303 = ~n79301 & ~n79302;
  assign n79304 = n79298 & ~n79303;
  assign n79305 = ~n79300 & ~n79304;
  assign n79306 = n79296 & ~n79298;
  assign n79307 = n79295 & n79306;
  assign n79308 = n79305 & ~n79307;
  assign n79309 = n79279 & ~n79308;
  assign n79310 = ~n79279 & n79308;
  assign n79311 = ~n79309 & ~n79310;
  assign n79312 = n79278 & ~n79311;
  assign n79313 = n79279 & ~n79307;
  assign n79314 = n79305 & n79313;
  assign n79315 = ~n79279 & ~n79308;
  assign n79316 = ~n79314 & ~n79315;
  assign n79317 = ~n79278 & ~n79316;
  assign n79318 = ~n79312 & ~n79317;
  assign n79319 = n79274 & ~n79318;
  assign n79320 = ~n79274 & n79318;
  assign n79321 = ~n79319 & ~n79320;
  assign n79322 = n79273 & ~n79321;
  assign n79323 = ~n79274 & ~n79318;
  assign n79324 = ~n79273 & n79323;
  assign n79325 = ~n79273 & n79274;
  assign n79326 = n79318 & n79325;
  assign n79327 = ~n79322 & ~n79324;
  assign n79328 = ~n79326 & n79327;
  assign n79329 = n79271 & ~n79328;
  assign n79330 = ~n79271 & n79328;
  assign n79331 = ~n79329 & ~n79330;
  assign n79332 = P3_DATAO_REG_13_ & n77688;
  assign n79333 = ~n78800 & n78801;
  assign n79334 = ~n78864 & ~n79333;
  assign n79335 = ~n78800 & n78858;
  assign n79336 = n79334 & ~n79335;
  assign n79337 = ~n79331 & ~n79332;
  assign n79338 = ~n79336 & n79337;
  assign n79339 = n79331 & n79332;
  assign n79340 = ~n79337 & ~n79339;
  assign n79341 = n79336 & n79340;
  assign n79342 = ~n79338 & ~n79341;
  assign n79343 = n79332 & ~n79336;
  assign n79344 = n79331 & n79343;
  assign n79345 = n79342 & ~n79344;
  assign n79346 = n79264 & ~n79345;
  assign n79347 = ~n79264 & n79345;
  assign n79348 = ~n79346 & ~n79347;
  assign n79349 = n79263 & ~n79348;
  assign n79350 = n79264 & ~n79344;
  assign n79351 = n79342 & n79350;
  assign n79352 = ~n79264 & ~n79345;
  assign n79353 = ~n79351 & ~n79352;
  assign n79354 = ~n79263 & ~n79353;
  assign n79355 = ~n79349 & ~n79354;
  assign n79356 = P3_DATAO_REG_11_ & n78036;
  assign n79357 = ~n78793 & n78878;
  assign n79358 = ~n78792 & ~n79357;
  assign n79359 = ~n79355 & ~n79356;
  assign n79360 = ~n79358 & n79359;
  assign n79361 = ~n79355 & n79356;
  assign n79362 = n79355 & ~n79356;
  assign n79363 = ~n79361 & ~n79362;
  assign n79364 = n79358 & ~n79363;
  assign n79365 = ~n79360 & ~n79364;
  assign n79366 = n79356 & ~n79358;
  assign n79367 = n79355 & n79366;
  assign n79368 = n79365 & ~n79367;
  assign n79369 = n79260 & ~n79368;
  assign n79370 = ~n79260 & n79368;
  assign n79371 = ~n79369 & ~n79370;
  assign n79372 = n79259 & ~n79371;
  assign n79373 = n79260 & ~n79367;
  assign n79374 = n79365 & n79373;
  assign n79375 = ~n79260 & ~n79368;
  assign n79376 = ~n79374 & ~n79375;
  assign n79377 = ~n79259 & ~n79376;
  assign n79378 = ~n79372 & ~n79377;
  assign n79379 = n79255 & ~n79378;
  assign n79380 = ~n79255 & n79378;
  assign n79381 = ~n79379 & ~n79380;
  assign n79382 = n79254 & ~n79381;
  assign n79383 = ~n79254 & n79381;
  assign n79384 = ~n79382 & ~n79383;
  assign n79385 = P3_DATAO_REG_8_ & n77722;
  assign n79386 = ~n79384 & ~n79385;
  assign n79387 = n79384 & n79385;
  assign n79388 = ~n78780 & ~n78892;
  assign n79389 = ~n78893 & ~n78899;
  assign n79390 = ~n79388 & n79389;
  assign n79391 = ~n79386 & ~n79387;
  assign n79392 = n79390 & n79391;
  assign n79393 = ~n79390 & ~n79391;
  assign n79394 = ~n79392 & ~n79393;
  assign n79395 = ~n78776 & n78777;
  assign n79396 = ~n78776 & n78902;
  assign n79397 = ~n78907 & ~n79395;
  assign n79398 = ~n79396 & n79397;
  assign n79399 = P3_DATAO_REG_7_ & n77720;
  assign n79400 = ~n79394 & ~n79398;
  assign n79401 = ~n79399 & n79400;
  assign n79402 = ~n79394 & n79398;
  assign n79403 = n79399 & n79402;
  assign n79404 = ~n79398 & n79399;
  assign n79405 = n79398 & ~n79399;
  assign n79406 = ~n79404 & ~n79405;
  assign n79407 = n79394 & ~n79406;
  assign n79408 = ~n79401 & ~n79403;
  assign n79409 = ~n79407 & n79408;
  assign n79410 = n79250 & ~n79409;
  assign n79411 = ~n79250 & n79409;
  assign n79412 = ~n79410 & ~n79411;
  assign n79413 = n79249 & ~n79412;
  assign n79414 = n79250 & n79409;
  assign n79415 = ~n79250 & ~n79409;
  assign n79416 = ~n79414 & ~n79415;
  assign n79417 = ~n79249 & ~n79416;
  assign n79418 = ~n79413 & ~n79417;
  assign n79419 = n79246 & ~n79418;
  assign n79420 = ~n79246 & n79418;
  assign n79421 = ~n79419 & ~n79420;
  assign n79422 = n79245 & ~n79421;
  assign n79423 = ~n79246 & ~n79418;
  assign n79424 = ~n79245 & n79423;
  assign n79425 = ~n79245 & n79246;
  assign n79426 = n79418 & n79425;
  assign n79427 = ~n79422 & ~n79424;
  assign n79428 = ~n79426 & n79427;
  assign n79429 = n79243 & ~n79428;
  assign n79430 = ~n79243 & n79428;
  assign n79431 = ~n79429 & ~n79430;
  assign n79432 = n79242 & ~n79431;
  assign n79433 = n79243 & n79428;
  assign n79434 = ~n79243 & ~n79428;
  assign n79435 = ~n79433 & ~n79434;
  assign n79436 = ~n79242 & ~n79435;
  assign n79437 = ~n79432 & ~n79436;
  assign n79438 = n79238 & ~n79437;
  assign n79439 = ~n79238 & n79437;
  assign n79440 = ~n79438 & ~n79439;
  assign n79441 = n79237 & ~n79440;
  assign n79442 = ~n79238 & ~n79437;
  assign n79443 = ~n79237 & n79442;
  assign n79444 = ~n79237 & n79238;
  assign n79445 = n79437 & n79444;
  assign n79446 = ~n79441 & ~n79443;
  assign n79447 = ~n79445 & n79446;
  assign n79448 = n79235 & ~n79447;
  assign n79449 = ~n79235 & n79447;
  assign n79450 = ~n79448 & ~n79449;
  assign n79451 = n77711 & ~n79450;
  assign n79452 = ~n77711 & n79450;
  assign n79453 = P3_DATAO_REG_1_ & n77712;
  assign n79454 = n77715 & n79082;
  assign n79455 = ~n77715 & ~n79082;
  assign n79456 = ~n79454 & ~n79455;
  assign n79457 = ~n79230 & ~n79456;
  assign n79458 = n79230 & n79456;
  assign n79459 = ~n79457 & ~n79458;
  assign n79460 = n79453 & n79459;
  assign n79461 = ~n79453 & ~n79459;
  assign n79462 = P3_DATAO_REG_1_ & n77714;
  assign n79463 = ~n79094 & n79224;
  assign n79464 = ~n79225 & ~n79463;
  assign n79465 = n79101 & ~n79464;
  assign n79466 = ~n79094 & ~n79224;
  assign n79467 = ~n79101 & n79466;
  assign n79468 = n79102 & n79224;
  assign n79469 = ~n79465 & ~n79467;
  assign n79470 = ~n79468 & n79469;
  assign n79471 = P3_DATAO_REG_1_ & n78934;
  assign n79472 = n79470 & n79471;
  assign n79473 = ~n79470 & ~n79471;
  assign n79474 = P3_DATAO_REG_1_ & n77716;
  assign n79475 = P3_DATAO_REG_1_ & n77718;
  assign n79476 = P3_DATAO_REG_1_ & n77720;
  assign n79477 = ~n79122 & n79123;
  assign n79478 = n79122 & ~n79123;
  assign n79479 = ~n79477 & ~n79478;
  assign n79480 = n79208 & ~n79479;
  assign n79481 = ~n79124 & ~n79125;
  assign n79482 = ~n79208 & ~n79481;
  assign n79483 = ~n79480 & ~n79482;
  assign n79484 = n79476 & ~n79483;
  assign n79485 = ~n79126 & n79204;
  assign n79486 = ~n79205 & ~n79485;
  assign n79487 = n79196 & ~n79486;
  assign n79488 = ~n79126 & ~n79204;
  assign n79489 = ~n79196 & n79488;
  assign n79490 = n79197 & n79204;
  assign n79491 = ~n79487 & ~n79489;
  assign n79492 = ~n79490 & n79491;
  assign n79493 = P3_DATAO_REG_1_ & n77722;
  assign n79494 = n79492 & n79493;
  assign n79495 = ~n79492 & ~n79493;
  assign n79496 = P3_DATAO_REG_1_ & n77724;
  assign n79497 = ~n79134 & n79135;
  assign n79498 = n79134 & ~n79135;
  assign n79499 = ~n79497 & ~n79498;
  assign n79500 = n79194 & ~n79499;
  assign n79501 = ~n79136 & ~n79137;
  assign n79502 = ~n79194 & ~n79501;
  assign n79503 = ~n79500 & ~n79502;
  assign n79504 = n79496 & ~n79503;
  assign n79505 = ~n79496 & n79503;
  assign n79506 = P3_DATAO_REG_1_ & n77726;
  assign n79507 = P3_DATAO_REG_1_ & n78036;
  assign n79508 = ~n79150 & n79166;
  assign n79509 = ~n79167 & ~n79508;
  assign n79510 = n79176 & ~n79509;
  assign n79511 = ~n79150 & ~n79166;
  assign n79512 = ~n79176 & n79511;
  assign n79513 = n79166 & n79177;
  assign n79514 = ~n79510 & ~n79512;
  assign n79515 = ~n79513 & n79514;
  assign n79516 = P3_DATAO_REG_1_ & n77955;
  assign n79517 = n79515 & n79516;
  assign n79518 = ~n79515 & ~n79516;
  assign n79519 = P3_DATAO_REG_1_ & n77688;
  assign n79520 = n79159 & ~n79164;
  assign n79521 = ~n79159 & n79164;
  assign n79522 = ~n79520 & ~n79521;
  assign n79523 = ~n79158 & n79522;
  assign n79524 = n79158 & n79521;
  assign n79525 = ~n79523 & ~n79524;
  assign n79526 = n79160 & ~n79164;
  assign n79527 = n79525 & ~n79526;
  assign n79528 = n79519 & ~n79527;
  assign n79529 = ~n79519 & n79527;
  assign n79530 = ~n77618 & ~n77684;
  assign n79531 = ~n77683 & ~n79530;
  assign n79532 = ~n79529 & ~n79531;
  assign n79533 = ~n79528 & ~n79532;
  assign n79534 = ~n79518 & ~n79533;
  assign n79535 = ~n79517 & ~n79534;
  assign n79536 = n79507 & ~n79535;
  assign n79537 = ~n79146 & n79147;
  assign n79538 = n79146 & ~n79147;
  assign n79539 = ~n79537 & ~n79538;
  assign n79540 = n79180 & ~n79539;
  assign n79541 = ~n79148 & ~n79149;
  assign n79542 = ~n79180 & ~n79541;
  assign n79543 = ~n79540 & ~n79542;
  assign n79544 = n79507 & ~n79543;
  assign n79545 = ~n79535 & ~n79543;
  assign n79546 = ~n79536 & ~n79544;
  assign n79547 = ~n79545 & n79546;
  assign n79548 = n79506 & ~n79547;
  assign n79549 = ~n79138 & n79190;
  assign n79550 = ~n79191 & ~n79549;
  assign n79551 = n79182 & ~n79550;
  assign n79552 = ~n79138 & ~n79190;
  assign n79553 = ~n79182 & n79552;
  assign n79554 = n79183 & n79190;
  assign n79555 = ~n79551 & ~n79553;
  assign n79556 = ~n79554 & n79555;
  assign n79557 = ~n79506 & n79547;
  assign n79558 = n79556 & ~n79557;
  assign n79559 = ~n79548 & ~n79558;
  assign n79560 = ~n79505 & ~n79559;
  assign n79561 = ~n79504 & ~n79560;
  assign n79562 = ~n79495 & ~n79561;
  assign n79563 = ~n79494 & ~n79562;
  assign n79564 = n79476 & ~n79563;
  assign n79565 = ~n79483 & ~n79563;
  assign n79566 = ~n79484 & ~n79564;
  assign n79567 = ~n79565 & n79566;
  assign n79568 = n79475 & ~n79567;
  assign n79569 = ~n79114 & n79218;
  assign n79570 = ~n79219 & ~n79569;
  assign n79571 = n79210 & ~n79570;
  assign n79572 = ~n79114 & ~n79218;
  assign n79573 = ~n79210 & n79572;
  assign n79574 = n79211 & n79218;
  assign n79575 = ~n79571 & ~n79573;
  assign n79576 = ~n79574 & n79575;
  assign n79577 = ~n79475 & n79567;
  assign n79578 = n79576 & ~n79577;
  assign n79579 = ~n79568 & ~n79578;
  assign n79580 = n79474 & ~n79579;
  assign n79581 = ~n79110 & n79111;
  assign n79582 = n79110 & ~n79111;
  assign n79583 = ~n79581 & ~n79582;
  assign n79584 = n79222 & ~n79583;
  assign n79585 = ~n79112 & ~n79113;
  assign n79586 = ~n79222 & ~n79585;
  assign n79587 = ~n79584 & ~n79586;
  assign n79588 = n79474 & ~n79587;
  assign n79589 = ~n79579 & ~n79587;
  assign n79590 = ~n79580 & ~n79588;
  assign n79591 = ~n79589 & n79590;
  assign n79592 = ~n79473 & ~n79591;
  assign n79593 = ~n79472 & ~n79592;
  assign n79594 = n79462 & ~n79593;
  assign n79595 = ~n79092 & ~n79093;
  assign n79596 = n79228 & n79595;
  assign n79597 = ~n79228 & ~n79595;
  assign n79598 = ~n79596 & ~n79597;
  assign n79599 = n79462 & ~n79598;
  assign n79600 = ~n79593 & ~n79598;
  assign n79601 = ~n79594 & ~n79599;
  assign n79602 = ~n79600 & n79601;
  assign n79603 = ~n79461 & ~n79602;
  assign n79604 = ~n79460 & ~n79603;
  assign n79605 = ~n79452 & ~n79604;
  assign n79606 = ~n79451 & ~n79605;
  assign n79607 = n77709 & ~n79606;
  assign n79608 = P3_DATAO_REG_2_ & n77710;
  assign n79609 = ~n79234 & n79447;
  assign n79610 = ~n79233 & ~n79609;
  assign n79611 = n79608 & ~n79610;
  assign n79612 = ~n79237 & ~n79437;
  assign n79613 = ~n79438 & ~n79444;
  assign n79614 = ~n79612 & n79613;
  assign n79615 = P3_DATAO_REG_3_ & n77712;
  assign n79616 = ~n79394 & n79399;
  assign n79617 = ~n79404 & ~n79616;
  assign n79618 = ~n79400 & n79617;
  assign n79619 = P3_DATAO_REG_7_ & n77718;
  assign n79620 = P3_DATAO_REG_10_ & n77724;
  assign n79621 = ~n79259 & ~n79375;
  assign n79622 = ~n79374 & ~n79621;
  assign n79623 = n79620 & ~n79622;
  assign n79624 = ~n79620 & n79622;
  assign n79625 = ~n79623 & ~n79624;
  assign n79626 = ~n79355 & ~n79358;
  assign n79627 = ~n79361 & ~n79366;
  assign n79628 = ~n79626 & n79627;
  assign n79629 = P3_DATAO_REG_11_ & n77726;
  assign n79630 = P3_DATAO_REG_13_ & n77955;
  assign n79631 = ~n79331 & n79332;
  assign n79632 = ~n79331 & ~n79336;
  assign n79633 = ~n79343 & ~n79631;
  assign n79634 = ~n79632 & n79633;
  assign n79635 = n79630 & ~n79634;
  assign n79636 = ~n79630 & n79634;
  assign n79637 = ~n79635 & ~n79636;
  assign n79638 = ~n79273 & ~n79318;
  assign n79639 = ~n79319 & ~n79325;
  assign n79640 = ~n79638 & n79639;
  assign n79641 = P3_DATAO_REG_15_ & n77434;
  assign n79642 = ~n79295 & ~n79298;
  assign n79643 = ~n79301 & ~n79306;
  assign n79644 = ~n79642 & n79643;
  assign n79645 = P3_DATAO_REG_17_ & n77475;
  assign n79646 = P3_DATAO_REG_19_ & n77440;
  assign n79647 = P3_DATAO_REG_20_ & n77442;
  assign n79648 = P3_DATAO_REG_21_ & n77444;
  assign n79649 = n79647 & ~n79648;
  assign n79650 = ~n79647 & n79648;
  assign n79651 = ~n79649 & ~n79650;
  assign n79652 = n79646 & ~n79651;
  assign n79653 = ~n79646 & n79651;
  assign n79654 = P3_DATAO_REG_19_ & P3_DATAO_REG_20_;
  assign n79655 = n77451 & n79654;
  assign n79656 = ~n79652 & ~n79653;
  assign n79657 = ~n79655 & n79656;
  assign n79658 = n79646 & ~n79649;
  assign n79659 = ~n79646 & n79649;
  assign n79660 = ~n79658 & ~n79659;
  assign n79661 = n79655 & n79660;
  assign n79662 = ~n79657 & ~n79661;
  assign n79663 = P3_DATAO_REG_18_ & n77438;
  assign n79664 = ~n79287 & n79289;
  assign n79665 = ~n79286 & ~n79664;
  assign n79666 = ~n79662 & ~n79663;
  assign n79667 = ~n79665 & n79666;
  assign n79668 = n79662 & n79663;
  assign n79669 = ~n79666 & ~n79668;
  assign n79670 = n79665 & n79669;
  assign n79671 = ~n79667 & ~n79670;
  assign n79672 = n79663 & ~n79665;
  assign n79673 = n79662 & n79672;
  assign n79674 = n79671 & ~n79673;
  assign n79675 = n79645 & ~n79674;
  assign n79676 = ~n79645 & n79674;
  assign n79677 = ~n79675 & ~n79676;
  assign n79678 = n79644 & ~n79677;
  assign n79679 = ~n79645 & n79673;
  assign n79680 = ~n79645 & ~n79671;
  assign n79681 = n79645 & n79671;
  assign n79682 = ~n79673 & n79681;
  assign n79683 = ~n79679 & ~n79680;
  assign n79684 = ~n79682 & n79683;
  assign n79685 = ~n79644 & ~n79684;
  assign n79686 = ~n79678 & ~n79685;
  assign n79687 = P3_DATAO_REG_16_ & n77436;
  assign n79688 = ~n79278 & ~n79315;
  assign n79689 = ~n79314 & ~n79688;
  assign n79690 = ~n79686 & ~n79687;
  assign n79691 = ~n79689 & n79690;
  assign n79692 = n79686 & n79687;
  assign n79693 = ~n79690 & ~n79692;
  assign n79694 = n79689 & n79693;
  assign n79695 = ~n79691 & ~n79694;
  assign n79696 = n79687 & ~n79689;
  assign n79697 = n79686 & n79696;
  assign n79698 = n79695 & ~n79697;
  assign n79699 = n79641 & ~n79698;
  assign n79700 = ~n79641 & n79698;
  assign n79701 = ~n79699 & ~n79700;
  assign n79702 = n79640 & ~n79701;
  assign n79703 = ~n79641 & n79697;
  assign n79704 = ~n79641 & ~n79695;
  assign n79705 = n79641 & ~n79697;
  assign n79706 = n79695 & n79705;
  assign n79707 = ~n79703 & ~n79704;
  assign n79708 = ~n79706 & n79707;
  assign n79709 = ~n79640 & ~n79708;
  assign n79710 = ~n79702 & ~n79709;
  assign n79711 = P3_DATAO_REG_14_ & n77688;
  assign n79712 = ~n79270 & n79328;
  assign n79713 = ~n79269 & ~n79712;
  assign n79714 = ~n79710 & ~n79711;
  assign n79715 = ~n79713 & n79714;
  assign n79716 = ~n79710 & n79711;
  assign n79717 = n79710 & ~n79711;
  assign n79718 = ~n79716 & ~n79717;
  assign n79719 = n79713 & ~n79718;
  assign n79720 = ~n79715 & ~n79719;
  assign n79721 = n79711 & ~n79713;
  assign n79722 = n79710 & n79721;
  assign n79723 = n79720 & ~n79722;
  assign n79724 = n79637 & ~n79723;
  assign n79725 = ~n79630 & ~n79632;
  assign n79726 = ~n79343 & n79725;
  assign n79727 = ~n79631 & n79726;
  assign n79728 = ~n79635 & ~n79727;
  assign n79729 = n79723 & ~n79728;
  assign n79730 = ~n79724 & ~n79729;
  assign n79731 = P3_DATAO_REG_12_ & n78036;
  assign n79732 = ~n79263 & ~n79352;
  assign n79733 = ~n79351 & ~n79732;
  assign n79734 = ~n79730 & ~n79731;
  assign n79735 = ~n79733 & n79734;
  assign n79736 = ~n79730 & n79731;
  assign n79737 = n79730 & ~n79731;
  assign n79738 = ~n79736 & ~n79737;
  assign n79739 = n79733 & ~n79738;
  assign n79740 = ~n79735 & ~n79739;
  assign n79741 = n79731 & ~n79733;
  assign n79742 = n79730 & n79741;
  assign n79743 = n79740 & ~n79742;
  assign n79744 = n79629 & ~n79743;
  assign n79745 = ~n79629 & n79743;
  assign n79746 = ~n79744 & ~n79745;
  assign n79747 = n79628 & ~n79746;
  assign n79748 = n79629 & ~n79742;
  assign n79749 = n79740 & n79748;
  assign n79750 = ~n79629 & ~n79743;
  assign n79751 = ~n79749 & ~n79750;
  assign n79752 = ~n79628 & ~n79751;
  assign n79753 = ~n79747 & ~n79752;
  assign n79754 = ~n79625 & n79753;
  assign n79755 = n79625 & ~n79753;
  assign n79756 = ~n79754 & ~n79755;
  assign n79757 = P3_DATAO_REG_9_ & n77722;
  assign n79758 = ~n79756 & ~n79757;
  assign n79759 = n79756 & n79757;
  assign n79760 = ~n77724 & n79378;
  assign n79761 = ~n79254 & ~n79760;
  assign n79762 = ~n79379 & ~n79761;
  assign n79763 = ~n79758 & ~n79759;
  assign n79764 = n79762 & n79763;
  assign n79765 = ~n79762 & ~n79763;
  assign n79766 = ~n79764 & ~n79765;
  assign n79767 = P3_DATAO_REG_8_ & n77720;
  assign n79768 = n79385 & ~n79390;
  assign n79769 = n79384 & ~n79390;
  assign n79770 = ~n79387 & ~n79768;
  assign n79771 = ~n79769 & n79770;
  assign n79772 = ~n79766 & ~n79767;
  assign n79773 = ~n79771 & n79772;
  assign n79774 = ~n79766 & n79767;
  assign n79775 = n79766 & ~n79767;
  assign n79776 = ~n79774 & ~n79775;
  assign n79777 = n79771 & ~n79776;
  assign n79778 = ~n79773 & ~n79777;
  assign n79779 = n79767 & ~n79771;
  assign n79780 = n79766 & n79779;
  assign n79781 = n79778 & ~n79780;
  assign n79782 = n79619 & ~n79781;
  assign n79783 = ~n79619 & n79781;
  assign n79784 = ~n79782 & ~n79783;
  assign n79785 = n79618 & ~n79784;
  assign n79786 = n79619 & n79778;
  assign n79787 = ~n79780 & n79786;
  assign n79788 = ~n79619 & ~n79781;
  assign n79789 = ~n79787 & ~n79788;
  assign n79790 = ~n79618 & ~n79789;
  assign n79791 = ~n79785 & ~n79790;
  assign n79792 = P3_DATAO_REG_6_ & n77716;
  assign n79793 = ~n79791 & ~n79792;
  assign n79794 = n79791 & n79792;
  assign n79795 = ~n79793 & ~n79794;
  assign n79796 = ~n79249 & ~n79415;
  assign n79797 = ~n79414 & ~n79796;
  assign n79798 = ~n79795 & ~n79797;
  assign n79799 = ~n79791 & n79792;
  assign n79800 = n79791 & ~n79792;
  assign n79801 = ~n79799 & ~n79800;
  assign n79802 = n79797 & ~n79801;
  assign n79803 = ~n79798 & ~n79802;
  assign n79804 = P3_DATAO_REG_5_ & n78934;
  assign n79805 = ~n79803 & ~n79804;
  assign n79806 = n79803 & n79804;
  assign n79807 = ~n79245 & ~n79418;
  assign n79808 = ~n79419 & ~n79425;
  assign n79809 = ~n79807 & n79808;
  assign n79810 = ~n79805 & ~n79806;
  assign n79811 = n79809 & n79810;
  assign n79812 = ~n79809 & ~n79810;
  assign n79813 = ~n79811 & ~n79812;
  assign n79814 = P3_DATAO_REG_4_ & n77714;
  assign n79815 = ~n79242 & ~n79434;
  assign n79816 = ~n79433 & ~n79815;
  assign n79817 = ~n79813 & ~n79814;
  assign n79818 = ~n79816 & n79817;
  assign n79819 = ~n79813 & n79814;
  assign n79820 = n79813 & ~n79814;
  assign n79821 = ~n79819 & ~n79820;
  assign n79822 = n79816 & ~n79821;
  assign n79823 = ~n79818 & ~n79822;
  assign n79824 = n79814 & ~n79816;
  assign n79825 = n79813 & n79824;
  assign n79826 = n79823 & ~n79825;
  assign n79827 = n79615 & ~n79826;
  assign n79828 = ~n79615 & n79826;
  assign n79829 = ~n79827 & ~n79828;
  assign n79830 = n79614 & ~n79829;
  assign n79831 = n79615 & n79826;
  assign n79832 = ~n79615 & ~n79826;
  assign n79833 = ~n79831 & ~n79832;
  assign n79834 = ~n79614 & ~n79833;
  assign n79835 = ~n79830 & ~n79834;
  assign n79836 = n79611 & n79835;
  assign n79837 = ~n79608 & ~n79835;
  assign n79838 = ~n79610 & n79837;
  assign n79839 = n79608 & ~n79835;
  assign n79840 = ~n79608 & n79835;
  assign n79841 = ~n79839 & ~n79840;
  assign n79842 = n79610 & ~n79841;
  assign n79843 = ~n79838 & ~n79842;
  assign n79844 = ~n77709 & n79606;
  assign n79845 = ~n79836 & n79843;
  assign n79846 = ~n79844 & n79845;
  assign n79847 = ~n79607 & ~n79846;
  assign n79848 = n77707 & ~n79847;
  assign n79849 = ~n79610 & ~n79835;
  assign n79850 = ~n79611 & ~n79839;
  assign n79851 = ~n79849 & n79850;
  assign n79852 = P3_DATAO_REG_2_ & n77708;
  assign n79853 = ~n79614 & ~n79832;
  assign n79854 = ~n79831 & ~n79853;
  assign n79855 = P3_DATAO_REG_3_ & n77710;
  assign n79856 = P3_DATAO_REG_5_ & n77714;
  assign n79857 = ~n79805 & ~n79809;
  assign n79858 = ~n79806 & ~n79857;
  assign n79859 = n79856 & ~n79858;
  assign n79860 = ~n79856 & n79858;
  assign n79861 = ~n79859 & ~n79860;
  assign n79862 = ~n79797 & ~n79800;
  assign n79863 = ~n79799 & ~n79862;
  assign n79864 = P3_DATAO_REG_6_ & n78934;
  assign n79865 = ~n79618 & ~n79788;
  assign n79866 = ~n79787 & ~n79865;
  assign n79867 = P3_DATAO_REG_7_ & n77716;
  assign n79868 = P3_DATAO_REG_8_ & n77718;
  assign n79869 = ~n79766 & ~n79771;
  assign n79870 = ~n79774 & ~n79779;
  assign n79871 = ~n79869 & n79870;
  assign n79872 = n79868 & ~n79871;
  assign n79873 = ~n79868 & n79871;
  assign n79874 = n79620 & ~n79753;
  assign n79875 = ~n79620 & n79753;
  assign n79876 = ~n79622 & ~n79875;
  assign n79877 = ~n79874 & ~n79876;
  assign n79878 = P3_DATAO_REG_10_ & n77722;
  assign n79879 = P3_DATAO_REG_12_ & n77726;
  assign n79880 = ~n79730 & ~n79733;
  assign n79881 = ~n79736 & ~n79741;
  assign n79882 = ~n79880 & n79881;
  assign n79883 = n79879 & ~n79882;
  assign n79884 = ~n79879 & n79882;
  assign n79885 = ~n79883 & ~n79884;
  assign n79886 = P3_DATAO_REG_13_ & n78036;
  assign n79887 = ~n79636 & n79723;
  assign n79888 = ~n79635 & ~n79887;
  assign n79889 = ~n79886 & ~n79888;
  assign n79890 = ~n79710 & ~n79713;
  assign n79891 = ~n79716 & ~n79721;
  assign n79892 = ~n79890 & n79891;
  assign n79893 = P3_DATAO_REG_14_ & n77955;
  assign n79894 = ~n79641 & ~n79698;
  assign n79895 = ~n79640 & ~n79894;
  assign n79896 = ~n79706 & ~n79895;
  assign n79897 = ~n79686 & n79687;
  assign n79898 = ~n79686 & ~n79689;
  assign n79899 = ~n79696 & ~n79897;
  assign n79900 = ~n79898 & n79899;
  assign n79901 = P3_DATAO_REG_16_ & n77434;
  assign n79902 = ~n79662 & n79663;
  assign n79903 = ~n79662 & ~n79665;
  assign n79904 = ~n79672 & ~n79902;
  assign n79905 = ~n79903 & n79904;
  assign n79906 = P3_DATAO_REG_18_ & n77475;
  assign n79907 = P3_DATAO_REG_20_ & n77440;
  assign n79908 = P3_DATAO_REG_21_ & n77442;
  assign n79909 = P3_DATAO_REG_22_ & n77444;
  assign n79910 = n79908 & ~n79909;
  assign n79911 = ~n79908 & n79909;
  assign n79912 = ~n79910 & ~n79911;
  assign n79913 = n79907 & ~n79912;
  assign n79914 = ~n79907 & n79912;
  assign n79915 = P3_DATAO_REG_20_ & P3_DATAO_REG_21_;
  assign n79916 = n77451 & n79915;
  assign n79917 = ~n79913 & ~n79914;
  assign n79918 = ~n79916 & n79917;
  assign n79919 = ~n79907 & ~n79910;
  assign n79920 = n79907 & ~n79909;
  assign n79921 = ~n79919 & ~n79920;
  assign n79922 = n79916 & ~n79921;
  assign n79923 = ~n79918 & ~n79922;
  assign n79924 = P3_DATAO_REG_19_ & n77438;
  assign n79925 = ~n79653 & n79655;
  assign n79926 = ~n79652 & ~n79925;
  assign n79927 = ~n79923 & ~n79924;
  assign n79928 = ~n79926 & n79927;
  assign n79929 = n79923 & n79924;
  assign n79930 = ~n79927 & ~n79929;
  assign n79931 = n79926 & n79930;
  assign n79932 = ~n79928 & ~n79931;
  assign n79933 = n79924 & ~n79926;
  assign n79934 = n79923 & n79933;
  assign n79935 = n79932 & ~n79934;
  assign n79936 = n79906 & ~n79935;
  assign n79937 = ~n79906 & n79935;
  assign n79938 = ~n79936 & ~n79937;
  assign n79939 = n79905 & ~n79938;
  assign n79940 = ~n79906 & n79934;
  assign n79941 = ~n79906 & ~n79932;
  assign n79942 = n79906 & n79932;
  assign n79943 = ~n79934 & n79942;
  assign n79944 = ~n79940 & ~n79941;
  assign n79945 = ~n79943 & n79944;
  assign n79946 = ~n79905 & ~n79945;
  assign n79947 = ~n79939 & ~n79946;
  assign n79948 = P3_DATAO_REG_17_ & n77436;
  assign n79949 = ~n79645 & ~n79674;
  assign n79950 = ~n79644 & ~n79949;
  assign n79951 = ~n79682 & ~n79950;
  assign n79952 = ~n79947 & ~n79948;
  assign n79953 = ~n79951 & n79952;
  assign n79954 = n79947 & n79948;
  assign n79955 = ~n79952 & ~n79954;
  assign n79956 = n79951 & n79955;
  assign n79957 = ~n79953 & ~n79956;
  assign n79958 = n79948 & ~n79951;
  assign n79959 = n79947 & n79958;
  assign n79960 = n79957 & ~n79959;
  assign n79961 = n79901 & ~n79960;
  assign n79962 = ~n79901 & n79960;
  assign n79963 = ~n79961 & ~n79962;
  assign n79964 = n79900 & ~n79963;
  assign n79965 = n79901 & ~n79959;
  assign n79966 = n79957 & n79965;
  assign n79967 = ~n79901 & ~n79960;
  assign n79968 = ~n79966 & ~n79967;
  assign n79969 = ~n79900 & ~n79968;
  assign n79970 = ~n79964 & ~n79969;
  assign n79971 = P3_DATAO_REG_15_ & n77688;
  assign n79972 = n79896 & ~n79970;
  assign n79973 = n79971 & n79972;
  assign n79974 = n79896 & n79970;
  assign n79975 = ~n79971 & n79974;
  assign n79976 = ~n79973 & ~n79975;
  assign n79977 = ~n79896 & ~n79971;
  assign n79978 = ~n79970 & n79977;
  assign n79979 = ~n79896 & n79971;
  assign n79980 = n79970 & n79979;
  assign n79981 = ~n79978 & ~n79980;
  assign n79982 = n79976 & n79981;
  assign n79983 = n79893 & ~n79982;
  assign n79984 = ~n79893 & n79982;
  assign n79985 = ~n79983 & ~n79984;
  assign n79986 = n79892 & ~n79985;
  assign n79987 = n79893 & n79981;
  assign n79988 = n79976 & n79987;
  assign n79989 = ~n79893 & ~n79982;
  assign n79990 = ~n79988 & ~n79989;
  assign n79991 = ~n79892 & ~n79990;
  assign n79992 = ~n79986 & ~n79991;
  assign n79993 = n79889 & ~n79992;
  assign n79994 = n79886 & ~n79888;
  assign n79995 = ~n79635 & ~n79886;
  assign n79996 = ~n79887 & n79995;
  assign n79997 = ~n79994 & ~n79996;
  assign n79998 = n79992 & ~n79997;
  assign n79999 = ~n79993 & ~n79998;
  assign n80000 = n79886 & ~n79992;
  assign n80001 = n79888 & n80000;
  assign n80002 = n79999 & ~n80001;
  assign n80003 = n79885 & ~n80002;
  assign n80004 = ~n79879 & ~n79880;
  assign n80005 = ~n79741 & n80004;
  assign n80006 = ~n79736 & n80005;
  assign n80007 = ~n79883 & ~n80006;
  assign n80008 = n80002 & ~n80007;
  assign n80009 = ~n80003 & ~n80008;
  assign n80010 = P3_DATAO_REG_11_ & n77724;
  assign n80011 = ~n80009 & ~n80010;
  assign n80012 = ~n79628 & ~n79750;
  assign n80013 = ~n79749 & ~n80012;
  assign n80014 = n80011 & ~n80013;
  assign n80015 = ~n80009 & n80010;
  assign n80016 = n80009 & ~n80010;
  assign n80017 = ~n80015 & ~n80016;
  assign n80018 = n80013 & ~n80017;
  assign n80019 = ~n80014 & ~n80018;
  assign n80020 = n80010 & ~n80013;
  assign n80021 = n80009 & n80020;
  assign n80022 = n80019 & ~n80021;
  assign n80023 = n79878 & ~n80022;
  assign n80024 = ~n79878 & n80022;
  assign n80025 = ~n80023 & ~n80024;
  assign n80026 = n79877 & ~n80025;
  assign n80027 = n79878 & ~n80021;
  assign n80028 = n80019 & n80027;
  assign n80029 = ~n79878 & ~n80022;
  assign n80030 = ~n80028 & ~n80029;
  assign n80031 = ~n79877 & ~n80030;
  assign n80032 = ~n80026 & ~n80031;
  assign n80033 = P3_DATAO_REG_9_ & n77720;
  assign n80034 = ~n79758 & ~n79762;
  assign n80035 = ~n79759 & ~n80034;
  assign n80036 = ~n80032 & ~n80033;
  assign n80037 = ~n80035 & n80036;
  assign n80038 = ~n80032 & n80033;
  assign n80039 = n80032 & ~n80033;
  assign n80040 = ~n80038 & ~n80039;
  assign n80041 = n80035 & ~n80040;
  assign n80042 = ~n80037 & ~n80041;
  assign n80043 = n80033 & ~n80035;
  assign n80044 = n80032 & n80043;
  assign n80045 = n80042 & ~n80044;
  assign n80046 = ~n79872 & ~n79873;
  assign n80047 = ~n80045 & n80046;
  assign n80048 = ~n79868 & ~n79869;
  assign n80049 = ~n79779 & n80048;
  assign n80050 = ~n79774 & n80049;
  assign n80051 = ~n79872 & ~n80050;
  assign n80052 = n80045 & ~n80051;
  assign n80053 = ~n80047 & ~n80052;
  assign n80054 = n79867 & ~n80053;
  assign n80055 = ~n79867 & n80053;
  assign n80056 = ~n80054 & ~n80055;
  assign n80057 = n79866 & ~n80056;
  assign n80058 = ~n79867 & ~n80053;
  assign n80059 = ~n79866 & n80058;
  assign n80060 = ~n79866 & n79867;
  assign n80061 = n80053 & n80060;
  assign n80062 = ~n80057 & ~n80059;
  assign n80063 = ~n80061 & n80062;
  assign n80064 = n79864 & ~n80063;
  assign n80065 = ~n79864 & n80063;
  assign n80066 = ~n80064 & ~n80065;
  assign n80067 = n79863 & ~n80066;
  assign n80068 = n79864 & n80063;
  assign n80069 = ~n79864 & ~n80063;
  assign n80070 = ~n80068 & ~n80069;
  assign n80071 = ~n79863 & ~n80070;
  assign n80072 = ~n80067 & ~n80071;
  assign n80073 = ~n79861 & n80072;
  assign n80074 = n79861 & ~n80072;
  assign n80075 = ~n80073 & ~n80074;
  assign n80076 = P3_DATAO_REG_4_ & n77712;
  assign n80077 = ~n80075 & ~n80076;
  assign n80078 = n80075 & n80076;
  assign n80079 = ~n79813 & ~n79816;
  assign n80080 = ~n79819 & ~n79824;
  assign n80081 = ~n80079 & n80080;
  assign n80082 = ~n80077 & ~n80078;
  assign n80083 = n80081 & n80082;
  assign n80084 = ~n80081 & ~n80082;
  assign n80085 = ~n80083 & ~n80084;
  assign n80086 = n79855 & ~n80085;
  assign n80087 = ~n79855 & n80085;
  assign n80088 = ~n80086 & ~n80087;
  assign n80089 = n79854 & ~n80088;
  assign n80090 = ~n79855 & ~n80085;
  assign n80091 = ~n79854 & n80090;
  assign n80092 = n79855 & n80085;
  assign n80093 = ~n79854 & n80092;
  assign n80094 = ~n80089 & ~n80091;
  assign n80095 = ~n80093 & n80094;
  assign n80096 = n79852 & ~n80095;
  assign n80097 = ~n79852 & n80095;
  assign n80098 = ~n80096 & ~n80097;
  assign n80099 = n79851 & ~n80098;
  assign n80100 = n79852 & n80095;
  assign n80101 = ~n79852 & ~n80095;
  assign n80102 = ~n80100 & ~n80101;
  assign n80103 = ~n79851 & ~n80102;
  assign n80104 = ~n80099 & ~n80103;
  assign n80105 = n77707 & ~n80104;
  assign n80106 = ~n79847 & ~n80104;
  assign n80107 = ~n79848 & ~n80105;
  assign n80108 = ~n80106 & n80107;
  assign n80109 = ~SEL & DIN_22_;
  assign n80110 = P3_DATAO_REG_1_ & n80109;
  assign n80111 = n80108 & ~n80110;
  assign n80112 = ~n80108 & n80110;
  assign n80113 = P3_DATAO_REG_4_ & n77710;
  assign n80114 = ~n80077 & ~n80081;
  assign n80115 = ~n80078 & ~n80114;
  assign n80116 = n80113 & ~n80115;
  assign n80117 = ~n80113 & n80115;
  assign n80118 = ~n80116 & ~n80117;
  assign n80119 = n79856 & ~n80072;
  assign n80120 = ~n79856 & n80072;
  assign n80121 = ~n79858 & ~n80120;
  assign n80122 = ~n80119 & ~n80121;
  assign n80123 = P3_DATAO_REG_5_ & n77712;
  assign n80124 = P3_DATAO_REG_6_ & n77714;
  assign n80125 = ~n79863 & n79864;
  assign n80126 = ~n79863 & n80063;
  assign n80127 = ~n80068 & ~n80125;
  assign n80128 = ~n80126 & n80127;
  assign n80129 = ~n80124 & ~n80128;
  assign n80130 = ~n79866 & ~n80053;
  assign n80131 = ~n80054 & ~n80060;
  assign n80132 = ~n80130 & n80131;
  assign n80133 = P3_DATAO_REG_7_ & n78934;
  assign n80134 = ~n80032 & ~n80035;
  assign n80135 = ~n80038 & ~n80043;
  assign n80136 = ~n80134 & n80135;
  assign n80137 = P3_DATAO_REG_9_ & n77718;
  assign n80138 = ~n80009 & ~n80013;
  assign n80139 = ~n80015 & ~n80020;
  assign n80140 = ~n80138 & n80139;
  assign n80141 = P3_DATAO_REG_11_ & n77722;
  assign n80142 = ~n79888 & ~n79992;
  assign n80143 = ~n79994 & ~n80000;
  assign n80144 = ~n80142 & n80143;
  assign n80145 = P3_DATAO_REG_13_ & n77726;
  assign n80146 = ~n79892 & n79893;
  assign n80147 = ~n79892 & n79982;
  assign n80148 = ~n79988 & ~n80146;
  assign n80149 = ~n80147 & n80148;
  assign n80150 = P3_DATAO_REG_14_ & n78036;
  assign n80151 = n80149 & ~n80150;
  assign n80152 = ~n79970 & n79971;
  assign n80153 = ~n79896 & ~n79970;
  assign n80154 = ~n79979 & ~n80152;
  assign n80155 = ~n80153 & n80154;
  assign n80156 = P3_DATAO_REG_15_ & n77955;
  assign n80157 = P3_DATAO_REG_16_ & n77688;
  assign n80158 = ~n79947 & n79948;
  assign n80159 = ~n79947 & ~n79951;
  assign n80160 = ~n79958 & ~n80158;
  assign n80161 = ~n80159 & n80160;
  assign n80162 = P3_DATAO_REG_17_ & n77434;
  assign n80163 = ~n79923 & n79924;
  assign n80164 = ~n79923 & ~n79926;
  assign n80165 = ~n79933 & ~n80163;
  assign n80166 = ~n80164 & n80165;
  assign n80167 = P3_DATAO_REG_19_ & n77475;
  assign n80168 = P3_DATAO_REG_21_ & n77440;
  assign n80169 = P3_DATAO_REG_22_ & n77442;
  assign n80170 = P3_DATAO_REG_23_ & n77444;
  assign n80171 = n80169 & ~n80170;
  assign n80172 = ~n80169 & n80170;
  assign n80173 = ~n80171 & ~n80172;
  assign n80174 = n80168 & ~n80173;
  assign n80175 = ~n80168 & n80173;
  assign n80176 = P3_DATAO_REG_21_ & P3_DATAO_REG_22_;
  assign n80177 = n77451 & n80176;
  assign n80178 = ~n80174 & ~n80175;
  assign n80179 = ~n80177 & n80178;
  assign n80180 = ~n80168 & ~n80171;
  assign n80181 = n80168 & ~n80170;
  assign n80182 = ~n80180 & ~n80181;
  assign n80183 = n80177 & ~n80182;
  assign n80184 = ~n80179 & ~n80183;
  assign n80185 = P3_DATAO_REG_20_ & n77438;
  assign n80186 = ~n79914 & n79916;
  assign n80187 = ~n79913 & ~n80186;
  assign n80188 = ~n80184 & ~n80185;
  assign n80189 = ~n80187 & n80188;
  assign n80190 = n80184 & n80185;
  assign n80191 = ~n80188 & ~n80190;
  assign n80192 = n80187 & n80191;
  assign n80193 = ~n80189 & ~n80192;
  assign n80194 = n80185 & ~n80187;
  assign n80195 = n80184 & n80194;
  assign n80196 = n80193 & ~n80195;
  assign n80197 = n80167 & ~n80196;
  assign n80198 = ~n80167 & n80196;
  assign n80199 = ~n80197 & ~n80198;
  assign n80200 = n80166 & ~n80199;
  assign n80201 = ~n80167 & n80195;
  assign n80202 = ~n80167 & ~n80193;
  assign n80203 = n80167 & n80193;
  assign n80204 = ~n80195 & n80203;
  assign n80205 = ~n80201 & ~n80202;
  assign n80206 = ~n80204 & n80205;
  assign n80207 = ~n80166 & ~n80206;
  assign n80208 = ~n80200 & ~n80207;
  assign n80209 = P3_DATAO_REG_18_ & n77436;
  assign n80210 = ~n79906 & ~n79935;
  assign n80211 = ~n79905 & ~n80210;
  assign n80212 = ~n79943 & ~n80211;
  assign n80213 = ~n80208 & ~n80209;
  assign n80214 = ~n80212 & n80213;
  assign n80215 = n80208 & n80209;
  assign n80216 = ~n80213 & ~n80215;
  assign n80217 = n80212 & n80216;
  assign n80218 = ~n80214 & ~n80217;
  assign n80219 = n80209 & ~n80212;
  assign n80220 = n80208 & n80219;
  assign n80221 = n80218 & ~n80220;
  assign n80222 = n80162 & ~n80221;
  assign n80223 = ~n80162 & n80221;
  assign n80224 = ~n80222 & ~n80223;
  assign n80225 = n80161 & ~n80224;
  assign n80226 = ~n80162 & n80220;
  assign n80227 = n80162 & ~n80220;
  assign n80228 = n80218 & n80227;
  assign n80229 = ~n80162 & ~n80218;
  assign n80230 = ~n80226 & ~n80228;
  assign n80231 = ~n80229 & n80230;
  assign n80232 = ~n80161 & ~n80231;
  assign n80233 = ~n80225 & ~n80232;
  assign n80234 = n80157 & ~n80233;
  assign n80235 = ~n79901 & n79959;
  assign n80236 = ~n79900 & ~n80235;
  assign n80237 = ~n79901 & ~n79957;
  assign n80238 = n80236 & ~n80237;
  assign n80239 = ~n79966 & ~n80238;
  assign n80240 = n80234 & n80239;
  assign n80241 = ~n80157 & ~n80233;
  assign n80242 = ~n80239 & n80241;
  assign n80243 = ~n80240 & ~n80242;
  assign n80244 = n80157 & ~n80239;
  assign n80245 = ~n79966 & ~n80157;
  assign n80246 = ~n80238 & n80245;
  assign n80247 = ~n80244 & ~n80246;
  assign n80248 = n80233 & ~n80247;
  assign n80249 = n80243 & ~n80248;
  assign n80250 = n80156 & ~n80249;
  assign n80251 = ~n80156 & n80249;
  assign n80252 = ~n80250 & ~n80251;
  assign n80253 = n80155 & ~n80252;
  assign n80254 = ~n80156 & n80233;
  assign n80255 = ~n80247 & n80254;
  assign n80256 = ~n80156 & ~n80243;
  assign n80257 = n80156 & ~n80248;
  assign n80258 = n80243 & n80257;
  assign n80259 = ~n80255 & ~n80256;
  assign n80260 = ~n80258 & n80259;
  assign n80261 = ~n80155 & ~n80260;
  assign n80262 = ~n80253 & ~n80261;
  assign n80263 = n80151 & n80262;
  assign n80264 = ~n80149 & n80150;
  assign n80265 = n80262 & n80264;
  assign n80266 = ~n80263 & ~n80265;
  assign n80267 = n80150 & ~n80262;
  assign n80268 = n80149 & n80267;
  assign n80269 = ~n80150 & ~n80262;
  assign n80270 = ~n80149 & n80269;
  assign n80271 = ~n80268 & ~n80270;
  assign n80272 = n80266 & n80271;
  assign n80273 = n80145 & ~n80272;
  assign n80274 = ~n80145 & n80272;
  assign n80275 = ~n80273 & ~n80274;
  assign n80276 = n80144 & ~n80275;
  assign n80277 = ~n80145 & ~n80271;
  assign n80278 = ~n80145 & ~n80266;
  assign n80279 = n80145 & n80271;
  assign n80280 = n80266 & n80279;
  assign n80281 = ~n80277 & ~n80278;
  assign n80282 = ~n80280 & n80281;
  assign n80283 = ~n80144 & ~n80282;
  assign n80284 = ~n80276 & ~n80283;
  assign n80285 = P3_DATAO_REG_12_ & n77724;
  assign n80286 = ~n80001 & ~n80006;
  assign n80287 = n79999 & n80286;
  assign n80288 = ~n79883 & ~n80287;
  assign n80289 = ~n80284 & ~n80285;
  assign n80290 = ~n80288 & n80289;
  assign n80291 = n80284 & n80285;
  assign n80292 = ~n80289 & ~n80291;
  assign n80293 = n80288 & n80292;
  assign n80294 = ~n80290 & ~n80293;
  assign n80295 = n80285 & ~n80288;
  assign n80296 = n80284 & n80295;
  assign n80297 = n80294 & ~n80296;
  assign n80298 = n80141 & ~n80297;
  assign n80299 = ~n80141 & n80297;
  assign n80300 = ~n80298 & ~n80299;
  assign n80301 = n80140 & ~n80300;
  assign n80302 = ~n80141 & n80296;
  assign n80303 = n80141 & ~n80296;
  assign n80304 = n80294 & n80303;
  assign n80305 = ~n80141 & ~n80294;
  assign n80306 = ~n80302 & ~n80304;
  assign n80307 = ~n80305 & n80306;
  assign n80308 = ~n80140 & ~n80307;
  assign n80309 = ~n80301 & ~n80308;
  assign n80310 = P3_DATAO_REG_10_ & n77720;
  assign n80311 = ~n79877 & ~n80029;
  assign n80312 = ~n80028 & ~n80311;
  assign n80313 = ~n80309 & ~n80310;
  assign n80314 = ~n80312 & n80313;
  assign n80315 = n80309 & n80310;
  assign n80316 = ~n80313 & ~n80315;
  assign n80317 = n80312 & n80316;
  assign n80318 = ~n80314 & ~n80317;
  assign n80319 = n80310 & ~n80312;
  assign n80320 = n80309 & n80319;
  assign n80321 = n80318 & ~n80320;
  assign n80322 = n80137 & ~n80321;
  assign n80323 = ~n80137 & n80321;
  assign n80324 = ~n80322 & ~n80323;
  assign n80325 = n80136 & ~n80324;
  assign n80326 = ~n80137 & n80320;
  assign n80327 = n80137 & ~n80320;
  assign n80328 = n80318 & n80327;
  assign n80329 = ~n80137 & ~n80318;
  assign n80330 = ~n80326 & ~n80328;
  assign n80331 = ~n80329 & n80330;
  assign n80332 = ~n80136 & ~n80331;
  assign n80333 = ~n80325 & ~n80332;
  assign n80334 = P3_DATAO_REG_8_ & n77716;
  assign n80335 = ~n79873 & n80045;
  assign n80336 = ~n79872 & ~n80335;
  assign n80337 = ~n80333 & ~n80334;
  assign n80338 = ~n80336 & n80337;
  assign n80339 = ~n80333 & n80334;
  assign n80340 = n80333 & ~n80334;
  assign n80341 = ~n80339 & ~n80340;
  assign n80342 = n80336 & ~n80341;
  assign n80343 = ~n80338 & ~n80342;
  assign n80344 = n80334 & ~n80336;
  assign n80345 = n80333 & n80344;
  assign n80346 = n80343 & ~n80345;
  assign n80347 = n80133 & ~n80346;
  assign n80348 = ~n80133 & n80346;
  assign n80349 = ~n80347 & ~n80348;
  assign n80350 = n80132 & ~n80349;
  assign n80351 = n80133 & ~n80345;
  assign n80352 = n80343 & n80351;
  assign n80353 = ~n80133 & ~n80346;
  assign n80354 = ~n80352 & ~n80353;
  assign n80355 = ~n80132 & ~n80354;
  assign n80356 = ~n80350 & ~n80355;
  assign n80357 = n80129 & ~n80356;
  assign n80358 = n80124 & ~n80128;
  assign n80359 = ~n80124 & n80128;
  assign n80360 = ~n80358 & ~n80359;
  assign n80361 = n80356 & ~n80360;
  assign n80362 = ~n80357 & ~n80361;
  assign n80363 = n80124 & ~n80356;
  assign n80364 = n80128 & n80363;
  assign n80365 = n80362 & ~n80364;
  assign n80366 = n80123 & ~n80365;
  assign n80367 = ~n80123 & n80365;
  assign n80368 = ~n80366 & ~n80367;
  assign n80369 = n80122 & ~n80368;
  assign n80370 = n80123 & n80362;
  assign n80371 = ~n80364 & n80370;
  assign n80372 = ~n80123 & ~n80365;
  assign n80373 = ~n80371 & ~n80372;
  assign n80374 = ~n80122 & ~n80373;
  assign n80375 = ~n80369 & ~n80374;
  assign n80376 = ~n80118 & n80375;
  assign n80377 = n80118 & ~n80375;
  assign n80378 = ~n80376 & ~n80377;
  assign n80379 = P3_DATAO_REG_3_ & n77708;
  assign n80380 = ~n80378 & ~n80379;
  assign n80381 = n80378 & n80379;
  assign n80382 = ~n79854 & n79855;
  assign n80383 = ~n79854 & ~n80085;
  assign n80384 = ~n80086 & ~n80382;
  assign n80385 = ~n80383 & n80384;
  assign n80386 = ~n80380 & ~n80381;
  assign n80387 = n80385 & n80386;
  assign n80388 = ~n80385 & ~n80386;
  assign n80389 = ~n80387 & ~n80388;
  assign n80390 = P3_DATAO_REG_2_ & n77706;
  assign n80391 = ~n79851 & ~n80101;
  assign n80392 = ~n80100 & ~n80391;
  assign n80393 = ~n80389 & ~n80390;
  assign n80394 = ~n80392 & n80393;
  assign n80395 = ~n80389 & n80390;
  assign n80396 = n80389 & ~n80390;
  assign n80397 = ~n80395 & ~n80396;
  assign n80398 = n80392 & ~n80397;
  assign n80399 = ~n80394 & ~n80398;
  assign n80400 = n80390 & ~n80392;
  assign n80401 = n80389 & n80400;
  assign n80402 = n80399 & ~n80401;
  assign n80403 = ~n80111 & ~n80112;
  assign n80404 = ~n80402 & n80403;
  assign n80405 = n80111 & n80402;
  assign n80406 = n80110 & ~n80401;
  assign n80407 = n80399 & n80406;
  assign n80408 = ~n80108 & n80407;
  assign n80409 = ~n80404 & ~n80405;
  assign n80410 = ~n80408 & n80409;
  assign n80411 = n77705 & ~n80410;
  assign n80412 = ~n77705 & n80410;
  assign n80413 = P3_DATAO_REG_0_ & n80109;
  assign n80414 = P3_DATAO_REG_0_ & n77706;
  assign n80415 = ~n79607 & ~n79844;
  assign n80416 = ~n79845 & n80415;
  assign n80417 = n79845 & ~n80415;
  assign n80418 = ~n80416 & ~n80417;
  assign n80419 = n80414 & ~n80418;
  assign n80420 = ~n80414 & n80418;
  assign n80421 = P3_DATAO_REG_0_ & n77708;
  assign n80422 = P3_DATAO_REG_0_ & n77710;
  assign n80423 = ~n79460 & ~n79461;
  assign n80424 = n79602 & n80423;
  assign n80425 = ~n79602 & ~n80423;
  assign n80426 = ~n80424 & ~n80425;
  assign n80427 = n80422 & ~n80426;
  assign n80428 = ~n80422 & n80426;
  assign n80429 = P3_DATAO_REG_0_ & n77712;
  assign n80430 = P3_DATAO_REG_0_ & n77714;
  assign n80431 = ~n79474 & n79587;
  assign n80432 = ~n79588 & ~n80431;
  assign n80433 = n79579 & ~n80432;
  assign n80434 = ~n79474 & ~n79587;
  assign n80435 = ~n79579 & n80434;
  assign n80436 = n79580 & n79587;
  assign n80437 = ~n80433 & ~n80435;
  assign n80438 = ~n80436 & n80437;
  assign n80439 = P3_DATAO_REG_0_ & n78934;
  assign n80440 = n80438 & n80439;
  assign n80441 = ~n80438 & ~n80439;
  assign n80442 = P3_DATAO_REG_0_ & n77716;
  assign n80443 = ~n79568 & ~n79577;
  assign n80444 = ~n79576 & n80443;
  assign n80445 = n79576 & ~n80443;
  assign n80446 = ~n80444 & ~n80445;
  assign n80447 = n80442 & ~n80446;
  assign n80448 = ~n80442 & n80446;
  assign n80449 = ~n79476 & n79563;
  assign n80450 = ~n79564 & ~n80449;
  assign n80451 = n79483 & ~n80450;
  assign n80452 = ~n79476 & ~n79563;
  assign n80453 = ~n79483 & n80452;
  assign n80454 = n79484 & n79563;
  assign n80455 = ~n80451 & ~n80453;
  assign n80456 = ~n80454 & n80455;
  assign n80457 = P3_DATAO_REG_0_ & n77718;
  assign n80458 = n80456 & n80457;
  assign n80459 = ~n80456 & ~n80457;
  assign n80460 = P3_DATAO_REG_0_ & n77720;
  assign n80461 = ~n79492 & n79493;
  assign n80462 = n79492 & ~n79493;
  assign n80463 = ~n80461 & ~n80462;
  assign n80464 = n79561 & ~n80463;
  assign n80465 = ~n79494 & ~n79495;
  assign n80466 = ~n79561 & ~n80465;
  assign n80467 = ~n80464 & ~n80466;
  assign n80468 = n80460 & ~n80467;
  assign n80469 = ~n80460 & n80467;
  assign n80470 = P3_DATAO_REG_0_ & n77722;
  assign n80471 = n79496 & ~n79559;
  assign n80472 = ~n79496 & n79559;
  assign n80473 = ~n80471 & ~n80472;
  assign n80474 = n79503 & ~n80473;
  assign n80475 = ~n79503 & n80473;
  assign n80476 = ~n80474 & ~n80475;
  assign n80477 = n80470 & n80476;
  assign n80478 = ~n80470 & ~n80476;
  assign n80479 = P3_DATAO_REG_0_ & n77724;
  assign n80480 = ~n79548 & ~n79557;
  assign n80481 = ~n79556 & n80480;
  assign n80482 = n79556 & ~n80480;
  assign n80483 = ~n80481 & ~n80482;
  assign n80484 = n80479 & ~n80483;
  assign n80485 = ~n80479 & n80483;
  assign n80486 = ~n79507 & n79543;
  assign n80487 = ~n79544 & ~n80486;
  assign n80488 = n79535 & ~n80487;
  assign n80489 = ~n79507 & ~n79543;
  assign n80490 = ~n79535 & n80489;
  assign n80491 = n79536 & n79543;
  assign n80492 = ~n80488 & ~n80490;
  assign n80493 = ~n80491 & n80492;
  assign n80494 = P3_DATAO_REG_0_ & n77726;
  assign n80495 = n80493 & n80494;
  assign n80496 = ~n80493 & ~n80494;
  assign n80497 = P3_DATAO_REG_0_ & n78036;
  assign n80498 = n79516 & ~n79533;
  assign n80499 = ~n79516 & n79533;
  assign n80500 = ~n80498 & ~n80499;
  assign n80501 = ~n79515 & n80500;
  assign n80502 = n79515 & n80499;
  assign n80503 = n79517 & ~n79533;
  assign n80504 = ~n80501 & ~n80502;
  assign n80505 = ~n80503 & n80504;
  assign n80506 = n80497 & ~n80505;
  assign n80507 = ~n80497 & n80505;
  assign n80508 = P3_DATAO_REG_0_ & n77955;
  assign n80509 = ~n77615 & ~n77694;
  assign n80510 = ~n77695 & ~n80509;
  assign n80511 = n80508 & ~n80510;
  assign n80512 = n79519 & ~n79531;
  assign n80513 = ~n79519 & n79531;
  assign n80514 = ~n80512 & ~n80513;
  assign n80515 = ~n79527 & ~n80514;
  assign n80516 = n79527 & n80514;
  assign n80517 = ~n80515 & ~n80516;
  assign n80518 = ~n80508 & n80510;
  assign n80519 = ~n80517 & ~n80518;
  assign n80520 = ~n80511 & ~n80519;
  assign n80521 = ~n80507 & ~n80520;
  assign n80522 = ~n80506 & ~n80521;
  assign n80523 = ~n80496 & ~n80522;
  assign n80524 = ~n80495 & ~n80523;
  assign n80525 = ~n80485 & ~n80524;
  assign n80526 = ~n80484 & ~n80525;
  assign n80527 = ~n80478 & ~n80526;
  assign n80528 = ~n80477 & ~n80527;
  assign n80529 = ~n80469 & ~n80528;
  assign n80530 = ~n80468 & ~n80529;
  assign n80531 = ~n80459 & ~n80530;
  assign n80532 = ~n80458 & ~n80531;
  assign n80533 = ~n80448 & ~n80532;
  assign n80534 = ~n80447 & ~n80533;
  assign n80535 = ~n80441 & ~n80534;
  assign n80536 = ~n80440 & ~n80535;
  assign n80537 = n80430 & ~n80536;
  assign n80538 = ~n79470 & n79471;
  assign n80539 = n79470 & ~n79471;
  assign n80540 = ~n80538 & ~n80539;
  assign n80541 = n79591 & ~n80540;
  assign n80542 = ~n79472 & ~n79473;
  assign n80543 = ~n79591 & ~n80542;
  assign n80544 = ~n80541 & ~n80543;
  assign n80545 = ~n80430 & n80536;
  assign n80546 = ~n80544 & ~n80545;
  assign n80547 = ~n80537 & ~n80546;
  assign n80548 = n80429 & ~n80547;
  assign n80549 = ~n79462 & n79598;
  assign n80550 = ~n79599 & ~n80549;
  assign n80551 = n79593 & ~n80550;
  assign n80552 = ~n79462 & ~n79598;
  assign n80553 = ~n79593 & n80552;
  assign n80554 = n79594 & n79598;
  assign n80555 = ~n80551 & ~n80553;
  assign n80556 = ~n80554 & n80555;
  assign n80557 = ~n80429 & n80547;
  assign n80558 = n80556 & ~n80557;
  assign n80559 = ~n80548 & ~n80558;
  assign n80560 = ~n80428 & ~n80559;
  assign n80561 = ~n80427 & ~n80560;
  assign n80562 = n80421 & ~n80561;
  assign n80563 = n77711 & ~n79604;
  assign n80564 = ~n77711 & n79604;
  assign n80565 = ~n80563 & ~n80564;
  assign n80566 = n79450 & ~n80565;
  assign n80567 = ~n79450 & n80565;
  assign n80568 = ~n80566 & ~n80567;
  assign n80569 = ~n80421 & n80561;
  assign n80570 = n80568 & ~n80569;
  assign n80571 = ~n80562 & ~n80570;
  assign n80572 = ~n80420 & ~n80571;
  assign n80573 = ~n80419 & ~n80572;
  assign n80574 = n80413 & ~n80573;
  assign n80575 = ~n77707 & n80104;
  assign n80576 = ~n80105 & ~n80575;
  assign n80577 = n79847 & ~n80576;
  assign n80578 = ~n77707 & ~n80104;
  assign n80579 = ~n79847 & n80578;
  assign n80580 = n79848 & n80104;
  assign n80581 = ~n80577 & ~n80579;
  assign n80582 = ~n80580 & n80581;
  assign n80583 = ~n80413 & n80573;
  assign n80584 = n80582 & ~n80583;
  assign n80585 = ~n80574 & ~n80584;
  assign n80586 = ~n80411 & ~n80412;
  assign n80587 = n80585 & n80586;
  assign n80588 = ~n80585 & ~n80586;
  assign n80589 = ~n80587 & ~n80588;
  assign n80590 = ~n12802 & ~n80589;
  assign n80591 = ~n77703 & ~n80590;
  assign n80592 = n77374 & n77429;
  assign n80593 = ~n80591 & n80592;
  assign n80594 = n77420 & n80593;
  assign n80595 = ~n77425 & ~n77428;
  assign n80596 = ~n77702 & n80595;
  assign n80597 = ~n80594 & n80596;
  assign n80598 = P2_BUF1_REG_31_ & n12802;
  assign n80599 = ~SEL & DIN_29_;
  assign n80600 = P3_DATAO_REG_1_ & n80599;
  assign n80601 = ~SEL & DIN_28_;
  assign n80602 = P3_DATAO_REG_1_ & n80601;
  assign n80603 = ~SEL & DIN_27_;
  assign n80604 = P3_DATAO_REG_2_ & n80603;
  assign n80605 = ~SEL & DIN_26_;
  assign n80606 = P3_DATAO_REG_2_ & n80605;
  assign n80607 = ~SEL & DIN_25_;
  assign n80608 = P3_DATAO_REG_2_ & n80607;
  assign n80609 = ~SEL & DIN_24_;
  assign n80610 = P3_DATAO_REG_2_ & n80609;
  assign n80611 = P3_DATAO_REG_4_ & n77706;
  assign n80612 = P3_DATAO_REG_4_ & n77708;
  assign n80613 = P3_DATAO_REG_5_ & n77710;
  assign n80614 = ~n80122 & ~n80372;
  assign n80615 = ~n80371 & ~n80614;
  assign n80616 = n80613 & ~n80615;
  assign n80617 = ~n80128 & ~n80356;
  assign n80618 = ~n80358 & ~n80363;
  assign n80619 = ~n80617 & n80618;
  assign n80620 = P3_DATAO_REG_6_ & n77712;
  assign n80621 = ~n80333 & ~n80336;
  assign n80622 = ~n80339 & ~n80344;
  assign n80623 = ~n80621 & n80622;
  assign n80624 = P3_DATAO_REG_8_ & n78934;
  assign n80625 = P3_DATAO_REG_12_ & n77722;
  assign n80626 = ~n80284 & n80285;
  assign n80627 = ~n80284 & ~n80288;
  assign n80628 = ~n80295 & ~n80626;
  assign n80629 = ~n80627 & n80628;
  assign n80630 = n80625 & ~n80629;
  assign n80631 = ~n80625 & n80629;
  assign n80632 = P3_DATAO_REG_14_ & n77726;
  assign n80633 = ~n80149 & ~n80262;
  assign n80634 = ~n80264 & ~n80267;
  assign n80635 = ~n80633 & n80634;
  assign n80636 = n80632 & ~n80635;
  assign n80637 = ~n80632 & n80635;
  assign n80638 = ~n80636 & ~n80637;
  assign n80639 = ~n80233 & ~n80239;
  assign n80640 = ~n80234 & ~n80244;
  assign n80641 = ~n80639 & n80640;
  assign n80642 = P3_DATAO_REG_16_ & n77955;
  assign n80643 = ~n80208 & n80209;
  assign n80644 = ~n80208 & ~n80212;
  assign n80645 = ~n80219 & ~n80643;
  assign n80646 = ~n80644 & n80645;
  assign n80647 = P3_DATAO_REG_18_ & n77434;
  assign n80648 = ~n80184 & n80185;
  assign n80649 = ~n80184 & ~n80187;
  assign n80650 = ~n80194 & ~n80648;
  assign n80651 = ~n80649 & n80650;
  assign n80652 = P3_DATAO_REG_20_ & n77475;
  assign n80653 = P3_DATAO_REG_22_ & n77440;
  assign n80654 = P3_DATAO_REG_23_ & n77442;
  assign n80655 = P3_DATAO_REG_24_ & n77444;
  assign n80656 = n80654 & ~n80655;
  assign n80657 = ~n80654 & n80655;
  assign n80658 = ~n80656 & ~n80657;
  assign n80659 = n80653 & ~n80658;
  assign n80660 = ~n80653 & n80658;
  assign n80661 = P3_DATAO_REG_22_ & P3_DATAO_REG_23_;
  assign n80662 = n77451 & n80661;
  assign n80663 = ~n80659 & ~n80660;
  assign n80664 = ~n80662 & n80663;
  assign n80665 = n80653 & ~n80656;
  assign n80666 = ~n80653 & n80656;
  assign n80667 = ~n80665 & ~n80666;
  assign n80668 = n80662 & n80667;
  assign n80669 = ~n80664 & ~n80668;
  assign n80670 = P3_DATAO_REG_21_ & n77438;
  assign n80671 = ~n80175 & n80177;
  assign n80672 = ~n80174 & ~n80671;
  assign n80673 = ~n80669 & ~n80670;
  assign n80674 = ~n80672 & n80673;
  assign n80675 = n80669 & n80670;
  assign n80676 = ~n80673 & ~n80675;
  assign n80677 = n80672 & n80676;
  assign n80678 = ~n80674 & ~n80677;
  assign n80679 = n80670 & ~n80672;
  assign n80680 = n80669 & n80679;
  assign n80681 = n80678 & ~n80680;
  assign n80682 = n80652 & ~n80681;
  assign n80683 = ~n80652 & n80681;
  assign n80684 = ~n80682 & ~n80683;
  assign n80685 = n80651 & ~n80684;
  assign n80686 = ~n80652 & n80680;
  assign n80687 = ~n80652 & ~n80678;
  assign n80688 = n80652 & n80678;
  assign n80689 = ~n80680 & n80688;
  assign n80690 = ~n80686 & ~n80687;
  assign n80691 = ~n80689 & n80690;
  assign n80692 = ~n80651 & ~n80691;
  assign n80693 = ~n80685 & ~n80692;
  assign n80694 = P3_DATAO_REG_19_ & n77436;
  assign n80695 = ~n80167 & ~n80196;
  assign n80696 = ~n80166 & ~n80695;
  assign n80697 = ~n80204 & ~n80696;
  assign n80698 = ~n80693 & ~n80694;
  assign n80699 = ~n80697 & n80698;
  assign n80700 = n80693 & n80694;
  assign n80701 = ~n80698 & ~n80700;
  assign n80702 = n80697 & n80701;
  assign n80703 = ~n80699 & ~n80702;
  assign n80704 = n80694 & ~n80697;
  assign n80705 = n80693 & n80704;
  assign n80706 = n80703 & ~n80705;
  assign n80707 = n80647 & ~n80706;
  assign n80708 = ~n80647 & n80706;
  assign n80709 = ~n80707 & ~n80708;
  assign n80710 = n80646 & ~n80709;
  assign n80711 = ~n80647 & n80705;
  assign n80712 = n80647 & ~n80705;
  assign n80713 = n80703 & n80712;
  assign n80714 = ~n80647 & ~n80703;
  assign n80715 = ~n80711 & ~n80713;
  assign n80716 = ~n80714 & n80715;
  assign n80717 = ~n80646 & ~n80716;
  assign n80718 = ~n80710 & ~n80717;
  assign n80719 = P3_DATAO_REG_17_ & n77688;
  assign n80720 = ~n80162 & ~n80221;
  assign n80721 = ~n80161 & ~n80720;
  assign n80722 = ~n80228 & ~n80721;
  assign n80723 = ~n80718 & ~n80719;
  assign n80724 = ~n80722 & n80723;
  assign n80725 = n80718 & n80719;
  assign n80726 = ~n80723 & ~n80725;
  assign n80727 = n80722 & n80726;
  assign n80728 = ~n80724 & ~n80727;
  assign n80729 = n80719 & ~n80722;
  assign n80730 = n80718 & n80729;
  assign n80731 = n80728 & ~n80730;
  assign n80732 = n80642 & ~n80731;
  assign n80733 = ~n80642 & n80731;
  assign n80734 = ~n80732 & ~n80733;
  assign n80735 = n80641 & ~n80734;
  assign n80736 = ~n80642 & n80730;
  assign n80737 = n80642 & ~n80730;
  assign n80738 = n80728 & n80737;
  assign n80739 = ~n80642 & ~n80728;
  assign n80740 = ~n80736 & ~n80738;
  assign n80741 = ~n80739 & n80740;
  assign n80742 = ~n80641 & ~n80741;
  assign n80743 = ~n80735 & ~n80742;
  assign n80744 = P3_DATAO_REG_15_ & n78036;
  assign n80745 = ~n80156 & ~n80249;
  assign n80746 = ~n80155 & ~n80745;
  assign n80747 = ~n80258 & ~n80746;
  assign n80748 = ~n80743 & ~n80744;
  assign n80749 = ~n80747 & n80748;
  assign n80750 = ~n80743 & n80744;
  assign n80751 = n80743 & ~n80744;
  assign n80752 = ~n80750 & ~n80751;
  assign n80753 = n80747 & ~n80752;
  assign n80754 = ~n80749 & ~n80753;
  assign n80755 = n80744 & ~n80747;
  assign n80756 = n80743 & n80755;
  assign n80757 = n80754 & ~n80756;
  assign n80758 = n80638 & ~n80757;
  assign n80759 = ~n80632 & ~n80633;
  assign n80760 = ~n80264 & n80759;
  assign n80761 = ~n80267 & n80760;
  assign n80762 = ~n80636 & ~n80761;
  assign n80763 = n80757 & ~n80762;
  assign n80764 = ~n80758 & ~n80763;
  assign n80765 = P3_DATAO_REG_13_ & n77724;
  assign n80766 = ~n80144 & n80145;
  assign n80767 = ~n80144 & n80272;
  assign n80768 = ~n80280 & ~n80766;
  assign n80769 = ~n80767 & n80768;
  assign n80770 = ~n80764 & ~n80765;
  assign n80771 = ~n80769 & n80770;
  assign n80772 = n80764 & n80765;
  assign n80773 = ~n80770 & ~n80772;
  assign n80774 = n80769 & n80773;
  assign n80775 = ~n80771 & ~n80774;
  assign n80776 = n80765 & ~n80769;
  assign n80777 = n80764 & n80776;
  assign n80778 = n80775 & ~n80777;
  assign n80779 = ~n80630 & ~n80631;
  assign n80780 = ~n80778 & n80779;
  assign n80781 = ~n80625 & ~n80627;
  assign n80782 = ~n80295 & n80781;
  assign n80783 = ~n80626 & n80782;
  assign n80784 = ~n80630 & ~n80783;
  assign n80785 = n80778 & ~n80784;
  assign n80786 = ~n80780 & ~n80785;
  assign n80787 = P3_DATAO_REG_11_ & n77720;
  assign n80788 = ~n80786 & ~n80787;
  assign n80789 = ~n80141 & ~n80297;
  assign n80790 = ~n80140 & ~n80789;
  assign n80791 = ~n80304 & ~n80790;
  assign n80792 = n80788 & ~n80791;
  assign n80793 = ~n80786 & n80787;
  assign n80794 = n80786 & ~n80787;
  assign n80795 = ~n80793 & ~n80794;
  assign n80796 = n80791 & ~n80795;
  assign n80797 = ~n80792 & ~n80796;
  assign n80798 = n80787 & ~n80791;
  assign n80799 = n80786 & n80798;
  assign n80800 = n80797 & ~n80799;
  assign n80801 = ~n80309 & n80310;
  assign n80802 = ~n80309 & ~n80312;
  assign n80803 = P3_DATAO_REG_10_ & n77718;
  assign n80804 = ~n80319 & ~n80801;
  assign n80805 = ~n80802 & n80804;
  assign n80806 = ~n80803 & n80805;
  assign n80807 = n80803 & ~n80805;
  assign n80808 = ~n80806 & ~n80807;
  assign n80809 = n80800 & ~n80808;
  assign n80810 = ~n80800 & n80808;
  assign n80811 = ~n80809 & ~n80810;
  assign n80812 = P3_DATAO_REG_9_ & n77716;
  assign n80813 = ~n80811 & ~n80812;
  assign n80814 = ~n80137 & ~n80321;
  assign n80815 = ~n80136 & ~n80814;
  assign n80816 = ~n80328 & ~n80815;
  assign n80817 = n80813 & ~n80816;
  assign n80818 = n80811 & n80812;
  assign n80819 = ~n80813 & ~n80818;
  assign n80820 = n80816 & n80819;
  assign n80821 = ~n80817 & ~n80820;
  assign n80822 = n80812 & ~n80816;
  assign n80823 = n80811 & n80822;
  assign n80824 = n80821 & ~n80823;
  assign n80825 = n80624 & ~n80824;
  assign n80826 = ~n80624 & n80824;
  assign n80827 = ~n80825 & ~n80826;
  assign n80828 = n80623 & ~n80827;
  assign n80829 = ~n80624 & n80823;
  assign n80830 = ~n80624 & ~n80821;
  assign n80831 = n80624 & ~n80823;
  assign n80832 = n80821 & n80831;
  assign n80833 = ~n80829 & ~n80830;
  assign n80834 = ~n80832 & n80833;
  assign n80835 = ~n80623 & ~n80834;
  assign n80836 = ~n80828 & ~n80835;
  assign n80837 = P3_DATAO_REG_7_ & n77714;
  assign n80838 = ~n80132 & n80133;
  assign n80839 = ~n80132 & ~n80345;
  assign n80840 = n80343 & n80839;
  assign n80841 = ~n80352 & ~n80838;
  assign n80842 = ~n80840 & n80841;
  assign n80843 = ~n80836 & ~n80837;
  assign n80844 = ~n80842 & n80843;
  assign n80845 = n80836 & n80837;
  assign n80846 = ~n80843 & ~n80845;
  assign n80847 = n80842 & n80846;
  assign n80848 = ~n80844 & ~n80847;
  assign n80849 = ~n80842 & n80845;
  assign n80850 = n80848 & ~n80849;
  assign n80851 = n80620 & ~n80850;
  assign n80852 = ~n80620 & n80850;
  assign n80853 = ~n80851 & ~n80852;
  assign n80854 = n80619 & ~n80853;
  assign n80855 = n80620 & ~n80849;
  assign n80856 = n80848 & n80855;
  assign n80857 = ~n80620 & ~n80850;
  assign n80858 = ~n80856 & ~n80857;
  assign n80859 = ~n80619 & ~n80858;
  assign n80860 = ~n80854 & ~n80859;
  assign n80861 = n80616 & n80860;
  assign n80862 = n80612 & ~n80861;
  assign n80863 = ~n80613 & ~n80860;
  assign n80864 = ~n80615 & n80863;
  assign n80865 = n80613 & ~n80860;
  assign n80866 = ~n80613 & n80860;
  assign n80867 = ~n80865 & ~n80866;
  assign n80868 = n80615 & ~n80867;
  assign n80869 = ~n80864 & ~n80868;
  assign n80870 = n80862 & n80869;
  assign n80871 = ~n80861 & n80869;
  assign n80872 = ~n80612 & ~n80871;
  assign n80873 = n80113 & ~n80375;
  assign n80874 = ~n80113 & n80375;
  assign n80875 = ~n80115 & ~n80874;
  assign n80876 = ~n80873 & ~n80875;
  assign n80877 = ~n80872 & ~n80876;
  assign n80878 = ~n80870 & ~n80877;
  assign n80879 = n80611 & ~n80878;
  assign n80880 = P3_DATAO_REG_5_ & n77708;
  assign n80881 = n80837 & ~n80842;
  assign n80882 = ~n80836 & n80837;
  assign n80883 = ~n80836 & ~n80842;
  assign n80884 = ~n80881 & ~n80882;
  assign n80885 = ~n80883 & n80884;
  assign n80886 = P3_DATAO_REG_7_ & n77712;
  assign n80887 = P3_DATAO_REG_8_ & n77714;
  assign n80888 = ~n80623 & n80833;
  assign n80889 = ~n80832 & ~n80888;
  assign n80890 = ~n80887 & ~n80889;
  assign n80891 = ~n80811 & n80812;
  assign n80892 = ~n80811 & ~n80816;
  assign n80893 = ~n80822 & ~n80891;
  assign n80894 = ~n80892 & n80893;
  assign n80895 = P3_DATAO_REG_9_ & n78934;
  assign n80896 = ~n80786 & ~n80791;
  assign n80897 = ~n80793 & ~n80798;
  assign n80898 = ~n80896 & n80897;
  assign n80899 = P3_DATAO_REG_11_ & n77718;
  assign n80900 = P3_DATAO_REG_14_ & n77724;
  assign n80901 = ~n80637 & n80757;
  assign n80902 = ~n80636 & ~n80901;
  assign n80903 = ~n80743 & ~n80747;
  assign n80904 = ~n80750 & ~n80755;
  assign n80905 = ~n80903 & n80904;
  assign n80906 = P3_DATAO_REG_15_ & n77726;
  assign n80907 = P3_DATAO_REG_16_ & n78036;
  assign n80908 = ~n80642 & ~n80731;
  assign n80909 = ~n80641 & ~n80908;
  assign n80910 = ~n80738 & ~n80909;
  assign n80911 = ~n80718 & n80719;
  assign n80912 = ~n80718 & ~n80722;
  assign n80913 = ~n80729 & ~n80911;
  assign n80914 = ~n80912 & n80913;
  assign n80915 = P3_DATAO_REG_17_ & n77955;
  assign n80916 = P3_DATAO_REG_18_ & n77688;
  assign n80917 = ~n80646 & ~n80711;
  assign n80918 = ~n80714 & n80917;
  assign n80919 = ~n80713 & ~n80918;
  assign n80920 = ~n80916 & ~n80919;
  assign n80921 = ~n80693 & n80694;
  assign n80922 = ~n80693 & ~n80697;
  assign n80923 = ~n80704 & ~n80921;
  assign n80924 = ~n80922 & n80923;
  assign n80925 = P3_DATAO_REG_19_ & n77434;
  assign n80926 = P3_DATAO_REG_20_ & n77436;
  assign n80927 = ~n80669 & n80670;
  assign n80928 = ~n80669 & ~n80672;
  assign n80929 = ~n80679 & ~n80927;
  assign n80930 = ~n80928 & n80929;
  assign n80931 = P3_DATAO_REG_21_ & n77475;
  assign n80932 = P3_DATAO_REG_23_ & n77440;
  assign n80933 = P3_DATAO_REG_24_ & n77442;
  assign n80934 = P3_DATAO_REG_25_ & n77444;
  assign n80935 = n80933 & ~n80934;
  assign n80936 = ~n80933 & n80934;
  assign n80937 = ~n80935 & ~n80936;
  assign n80938 = n80932 & ~n80937;
  assign n80939 = ~n80932 & n80937;
  assign n80940 = P3_DATAO_REG_23_ & P3_DATAO_REG_24_;
  assign n80941 = n77451 & n80940;
  assign n80942 = ~n80938 & ~n80939;
  assign n80943 = ~n80941 & n80942;
  assign n80944 = n80932 & ~n80935;
  assign n80945 = ~n80932 & n80935;
  assign n80946 = ~n80944 & ~n80945;
  assign n80947 = n80941 & n80946;
  assign n80948 = ~n80943 & ~n80947;
  assign n80949 = P3_DATAO_REG_22_ & n77438;
  assign n80950 = ~n80660 & n80662;
  assign n80951 = ~n80659 & ~n80950;
  assign n80952 = ~n80948 & ~n80949;
  assign n80953 = ~n80951 & n80952;
  assign n80954 = n80948 & n80949;
  assign n80955 = ~n80952 & ~n80954;
  assign n80956 = n80951 & n80955;
  assign n80957 = ~n80953 & ~n80956;
  assign n80958 = n80949 & ~n80951;
  assign n80959 = n80948 & n80958;
  assign n80960 = n80957 & ~n80959;
  assign n80961 = n80931 & ~n80960;
  assign n80962 = ~n80931 & n80960;
  assign n80963 = ~n80961 & ~n80962;
  assign n80964 = n80930 & ~n80963;
  assign n80965 = ~n80931 & n80959;
  assign n80966 = ~n80931 & ~n80957;
  assign n80967 = n80931 & n80957;
  assign n80968 = ~n80959 & n80967;
  assign n80969 = ~n80965 & ~n80966;
  assign n80970 = ~n80968 & n80969;
  assign n80971 = ~n80930 & ~n80970;
  assign n80972 = ~n80964 & ~n80971;
  assign n80973 = n80926 & ~n80972;
  assign n80974 = ~n80652 & ~n80681;
  assign n80975 = ~n80651 & ~n80974;
  assign n80976 = ~n80689 & ~n80975;
  assign n80977 = n80973 & n80976;
  assign n80978 = ~n80926 & ~n80972;
  assign n80979 = ~n80976 & n80978;
  assign n80980 = ~n80977 & ~n80979;
  assign n80981 = n80926 & ~n80976;
  assign n80982 = ~n80926 & n80976;
  assign n80983 = ~n80981 & ~n80982;
  assign n80984 = n80972 & ~n80983;
  assign n80985 = n80980 & ~n80984;
  assign n80986 = n80925 & ~n80985;
  assign n80987 = ~n80925 & n80985;
  assign n80988 = ~n80986 & ~n80987;
  assign n80989 = n80924 & ~n80988;
  assign n80990 = n80925 & ~n80984;
  assign n80991 = n80980 & n80990;
  assign n80992 = ~n80925 & ~n80985;
  assign n80993 = ~n80991 & ~n80992;
  assign n80994 = ~n80924 & ~n80993;
  assign n80995 = ~n80989 & ~n80994;
  assign n80996 = n80920 & ~n80995;
  assign n80997 = ~n80916 & n80919;
  assign n80998 = n80916 & ~n80919;
  assign n80999 = ~n80997 & ~n80998;
  assign n81000 = n80995 & ~n80999;
  assign n81001 = ~n80996 & ~n81000;
  assign n81002 = n80916 & n80919;
  assign n81003 = ~n80995 & n81002;
  assign n81004 = n81001 & ~n81003;
  assign n81005 = n80915 & ~n81004;
  assign n81006 = ~n80915 & n81004;
  assign n81007 = ~n81005 & ~n81006;
  assign n81008 = n80914 & ~n81007;
  assign n81009 = n80915 & ~n81003;
  assign n81010 = n81001 & n81009;
  assign n81011 = ~n80915 & ~n81004;
  assign n81012 = ~n81010 & ~n81011;
  assign n81013 = ~n80914 & ~n81012;
  assign n81014 = ~n81008 & ~n81013;
  assign n81015 = ~n80907 & ~n80910;
  assign n81016 = ~n81014 & n81015;
  assign n81017 = n80907 & ~n80910;
  assign n81018 = n81014 & n81017;
  assign n81019 = ~n81016 & ~n81018;
  assign n81020 = ~n80907 & ~n81014;
  assign n81021 = n80907 & n81014;
  assign n81022 = ~n81020 & ~n81021;
  assign n81023 = n80910 & n81022;
  assign n81024 = n81019 & ~n81023;
  assign n81025 = n80906 & ~n81024;
  assign n81026 = ~n80906 & n81024;
  assign n81027 = ~n81025 & ~n81026;
  assign n81028 = n80905 & ~n81027;
  assign n81029 = n80906 & n81019;
  assign n81030 = ~n81023 & n81029;
  assign n81031 = ~n80906 & ~n81024;
  assign n81032 = ~n81030 & ~n81031;
  assign n81033 = ~n80905 & ~n81032;
  assign n81034 = ~n81028 & ~n81033;
  assign n81035 = ~n80900 & ~n80902;
  assign n81036 = ~n81034 & n81035;
  assign n81037 = n80900 & ~n80902;
  assign n81038 = ~n80636 & ~n80900;
  assign n81039 = ~n80901 & n81038;
  assign n81040 = ~n81037 & ~n81039;
  assign n81041 = n81034 & ~n81040;
  assign n81042 = ~n81036 & ~n81041;
  assign n81043 = n80900 & ~n81034;
  assign n81044 = n80902 & n81043;
  assign n81045 = n81042 & ~n81044;
  assign n81046 = ~n80764 & n80765;
  assign n81047 = ~n80764 & ~n80769;
  assign n81048 = P3_DATAO_REG_13_ & n77722;
  assign n81049 = ~n80776 & ~n81046;
  assign n81050 = ~n81047 & n81049;
  assign n81051 = ~n81048 & n81050;
  assign n81052 = n81048 & ~n81050;
  assign n81053 = ~n81051 & ~n81052;
  assign n81054 = n81045 & ~n81053;
  assign n81055 = ~n81045 & n81053;
  assign n81056 = ~n81054 & ~n81055;
  assign n81057 = P3_DATAO_REG_12_ & n77720;
  assign n81058 = n80625 & ~n80777;
  assign n81059 = n80775 & n81058;
  assign n81060 = ~n80629 & n80778;
  assign n81061 = ~n80630 & ~n81059;
  assign n81062 = ~n81060 & n81061;
  assign n81063 = ~n81056 & ~n81057;
  assign n81064 = ~n81062 & n81063;
  assign n81065 = n81056 & n81057;
  assign n81066 = ~n81063 & ~n81065;
  assign n81067 = n81062 & n81066;
  assign n81068 = ~n81064 & ~n81067;
  assign n81069 = n81057 & ~n81062;
  assign n81070 = n81056 & n81069;
  assign n81071 = n81068 & ~n81070;
  assign n81072 = n80899 & ~n81071;
  assign n81073 = ~n80899 & n81071;
  assign n81074 = ~n81072 & ~n81073;
  assign n81075 = n80898 & ~n81074;
  assign n81076 = ~n80899 & ~n81068;
  assign n81077 = n80899 & n81068;
  assign n81078 = ~n81070 & n81077;
  assign n81079 = ~n80899 & n81070;
  assign n81080 = ~n81076 & ~n81078;
  assign n81081 = ~n81079 & n81080;
  assign n81082 = ~n80898 & ~n81081;
  assign n81083 = ~n81075 & ~n81082;
  assign n81084 = P3_DATAO_REG_10_ & n77716;
  assign n81085 = ~n80802 & ~n80803;
  assign n81086 = ~n80319 & n81085;
  assign n81087 = ~n80801 & n81086;
  assign n81088 = ~n80799 & ~n81087;
  assign n81089 = n80797 & n81088;
  assign n81090 = ~n80807 & ~n81089;
  assign n81091 = ~n81083 & ~n81084;
  assign n81092 = ~n81090 & n81091;
  assign n81093 = n81083 & n81084;
  assign n81094 = ~n81091 & ~n81093;
  assign n81095 = n81090 & n81094;
  assign n81096 = ~n81092 & ~n81095;
  assign n81097 = n81084 & ~n81090;
  assign n81098 = n81083 & n81097;
  assign n81099 = n81096 & ~n81098;
  assign n81100 = n80895 & ~n81099;
  assign n81101 = ~n80895 & n81099;
  assign n81102 = ~n81100 & ~n81101;
  assign n81103 = n80894 & ~n81102;
  assign n81104 = ~n80895 & n81098;
  assign n81105 = ~n80895 & ~n81096;
  assign n81106 = n80895 & ~n81098;
  assign n81107 = n81096 & n81106;
  assign n81108 = ~n81104 & ~n81105;
  assign n81109 = ~n81107 & n81108;
  assign n81110 = ~n80894 & ~n81109;
  assign n81111 = ~n81103 & ~n81110;
  assign n81112 = n80890 & ~n81111;
  assign n81113 = n80832 & n80887;
  assign n81114 = ~n80887 & ~n80888;
  assign n81115 = ~n80832 & n81114;
  assign n81116 = n80887 & n80888;
  assign n81117 = ~n81113 & ~n81115;
  assign n81118 = ~n81116 & n81117;
  assign n81119 = n81111 & ~n81118;
  assign n81120 = ~n81112 & ~n81119;
  assign n81121 = n80887 & n80889;
  assign n81122 = ~n81111 & n81121;
  assign n81123 = n81120 & ~n81122;
  assign n81124 = n80886 & ~n81123;
  assign n81125 = ~n80886 & n81123;
  assign n81126 = ~n81124 & ~n81125;
  assign n81127 = n80885 & ~n81126;
  assign n81128 = ~n80886 & n81122;
  assign n81129 = n80886 & ~n81122;
  assign n81130 = n81120 & n81129;
  assign n81131 = ~n80886 & ~n81120;
  assign n81132 = ~n81128 & ~n81130;
  assign n81133 = ~n81131 & n81132;
  assign n81134 = ~n80885 & ~n81133;
  assign n81135 = ~n81127 & ~n81134;
  assign n81136 = P3_DATAO_REG_6_ & n77710;
  assign n81137 = ~n80619 & ~n80857;
  assign n81138 = ~n80856 & ~n81137;
  assign n81139 = ~n81135 & ~n81136;
  assign n81140 = ~n81138 & n81139;
  assign n81141 = n81135 & n81136;
  assign n81142 = ~n81139 & ~n81141;
  assign n81143 = n81138 & n81142;
  assign n81144 = ~n81140 & ~n81143;
  assign n81145 = n81136 & ~n81138;
  assign n81146 = n81135 & n81145;
  assign n81147 = n81144 & ~n81146;
  assign n81148 = n80880 & ~n81147;
  assign n81149 = ~n80880 & n81147;
  assign n81150 = ~n81148 & ~n81149;
  assign n81151 = ~n80615 & ~n80860;
  assign n81152 = ~n80616 & ~n80865;
  assign n81153 = ~n81151 & n81152;
  assign n81154 = ~n81150 & n81153;
  assign n81155 = ~n80880 & n81146;
  assign n81156 = n80880 & ~n81146;
  assign n81157 = n81144 & n81156;
  assign n81158 = ~n80880 & ~n81144;
  assign n81159 = ~n81155 & ~n81157;
  assign n81160 = ~n81158 & n81159;
  assign n81161 = ~n81153 & ~n81160;
  assign n81162 = ~n81154 & ~n81161;
  assign n81163 = n80611 & ~n81162;
  assign n81164 = ~n80878 & ~n81162;
  assign n81165 = ~n80879 & ~n81163;
  assign n81166 = ~n81164 & n81165;
  assign n81167 = P3_DATAO_REG_4_ & n80109;
  assign n81168 = P3_DATAO_REG_7_ & n77710;
  assign n81169 = ~n80885 & n80886;
  assign n81170 = ~n80885 & n81123;
  assign n81171 = ~n81130 & ~n81169;
  assign n81172 = ~n81170 & n81171;
  assign n81173 = n81168 & ~n81172;
  assign n81174 = ~n81168 & n81172;
  assign n81175 = ~n81173 & ~n81174;
  assign n81176 = n80887 & ~n81111;
  assign n81177 = n80887 & ~n80889;
  assign n81178 = ~n80889 & ~n81111;
  assign n81179 = ~n81176 & ~n81177;
  assign n81180 = ~n81178 & n81179;
  assign n81181 = P3_DATAO_REG_8_ & n77712;
  assign n81182 = ~n81083 & n81084;
  assign n81183 = ~n81083 & ~n81090;
  assign n81184 = ~n81097 & ~n81182;
  assign n81185 = ~n81183 & n81184;
  assign n81186 = P3_DATAO_REG_10_ & n78934;
  assign n81187 = P3_DATAO_REG_11_ & n77716;
  assign n81188 = ~n80898 & n80899;
  assign n81189 = ~n80898 & n81071;
  assign n81190 = ~n81078 & ~n81188;
  assign n81191 = ~n81189 & n81190;
  assign n81192 = P3_DATAO_REG_14_ & n77722;
  assign n81193 = ~n80902 & ~n81034;
  assign n81194 = ~n81037 & ~n81043;
  assign n81195 = ~n81193 & n81194;
  assign n81196 = n81192 & ~n81195;
  assign n81197 = ~n81192 & n81195;
  assign n81198 = ~n81196 & ~n81197;
  assign n81199 = ~n80905 & ~n81031;
  assign n81200 = ~n81030 & ~n81199;
  assign n81201 = n80907 & ~n81014;
  assign n81202 = ~n80910 & ~n81014;
  assign n81203 = ~n81017 & ~n81201;
  assign n81204 = ~n81202 & n81203;
  assign n81205 = P3_DATAO_REG_16_ & n77726;
  assign n81206 = n80916 & ~n80995;
  assign n81207 = ~n80919 & ~n80995;
  assign n81208 = ~n80998 & ~n81206;
  assign n81209 = ~n81207 & n81208;
  assign n81210 = P3_DATAO_REG_18_ & n77955;
  assign n81211 = ~n80972 & ~n80976;
  assign n81212 = ~n80973 & ~n80981;
  assign n81213 = ~n81211 & n81212;
  assign n81214 = P3_DATAO_REG_20_ & n77434;
  assign n81215 = ~n80948 & n80949;
  assign n81216 = ~n80948 & ~n80951;
  assign n81217 = ~n80958 & ~n81215;
  assign n81218 = ~n81216 & n81217;
  assign n81219 = P3_DATAO_REG_22_ & n77475;
  assign n81220 = P3_DATAO_REG_24_ & n77440;
  assign n81221 = P3_DATAO_REG_25_ & n77442;
  assign n81222 = P3_DATAO_REG_26_ & n77444;
  assign n81223 = n81221 & ~n81222;
  assign n81224 = ~n81221 & n81222;
  assign n81225 = ~n81223 & ~n81224;
  assign n81226 = n81220 & ~n81225;
  assign n81227 = ~n81220 & n81225;
  assign n81228 = P3_DATAO_REG_24_ & P3_DATAO_REG_25_;
  assign n81229 = n77451 & n81228;
  assign n81230 = ~n81226 & ~n81227;
  assign n81231 = ~n81229 & n81230;
  assign n81232 = ~n81220 & ~n81223;
  assign n81233 = n81220 & ~n81222;
  assign n81234 = ~n81232 & ~n81233;
  assign n81235 = n81229 & ~n81234;
  assign n81236 = ~n81231 & ~n81235;
  assign n81237 = P3_DATAO_REG_23_ & n77438;
  assign n81238 = ~n80939 & n80941;
  assign n81239 = ~n80938 & ~n81238;
  assign n81240 = ~n81236 & ~n81237;
  assign n81241 = ~n81239 & n81240;
  assign n81242 = n81236 & n81237;
  assign n81243 = ~n81240 & ~n81242;
  assign n81244 = n81239 & n81243;
  assign n81245 = ~n81241 & ~n81244;
  assign n81246 = n81237 & ~n81239;
  assign n81247 = n81236 & n81246;
  assign n81248 = n81245 & ~n81247;
  assign n81249 = n81219 & ~n81248;
  assign n81250 = ~n81219 & n81248;
  assign n81251 = ~n81249 & ~n81250;
  assign n81252 = n81218 & ~n81251;
  assign n81253 = ~n81219 & n81247;
  assign n81254 = ~n81219 & ~n81245;
  assign n81255 = n81219 & n81245;
  assign n81256 = ~n81247 & n81255;
  assign n81257 = ~n81253 & ~n81254;
  assign n81258 = ~n81256 & n81257;
  assign n81259 = ~n81218 & ~n81258;
  assign n81260 = ~n81252 & ~n81259;
  assign n81261 = P3_DATAO_REG_21_ & n77436;
  assign n81262 = ~n80930 & n80931;
  assign n81263 = ~n80930 & n80960;
  assign n81264 = ~n80968 & ~n81262;
  assign n81265 = ~n81263 & n81264;
  assign n81266 = ~n81260 & ~n81261;
  assign n81267 = ~n81265 & n81266;
  assign n81268 = n81260 & n81261;
  assign n81269 = ~n81266 & ~n81268;
  assign n81270 = n81265 & n81269;
  assign n81271 = ~n81267 & ~n81270;
  assign n81272 = n81261 & ~n81265;
  assign n81273 = n81260 & n81272;
  assign n81274 = n81271 & ~n81273;
  assign n81275 = n81214 & ~n81274;
  assign n81276 = ~n81214 & n81274;
  assign n81277 = ~n81275 & ~n81276;
  assign n81278 = n81213 & ~n81277;
  assign n81279 = ~n81214 & n81273;
  assign n81280 = n81214 & ~n81273;
  assign n81281 = n81271 & n81280;
  assign n81282 = ~n81214 & ~n81271;
  assign n81283 = ~n81279 & ~n81281;
  assign n81284 = ~n81282 & n81283;
  assign n81285 = ~n81213 & ~n81284;
  assign n81286 = ~n81278 & ~n81285;
  assign n81287 = P3_DATAO_REG_19_ & n77688;
  assign n81288 = ~n80924 & ~n80992;
  assign n81289 = ~n80991 & ~n81288;
  assign n81290 = ~n81286 & ~n81287;
  assign n81291 = ~n81289 & n81290;
  assign n81292 = n81286 & n81287;
  assign n81293 = ~n81290 & ~n81292;
  assign n81294 = n81289 & n81293;
  assign n81295 = ~n81291 & ~n81294;
  assign n81296 = n81287 & ~n81289;
  assign n81297 = n81286 & n81296;
  assign n81298 = n81295 & ~n81297;
  assign n81299 = n81210 & ~n81298;
  assign n81300 = ~n81210 & n81298;
  assign n81301 = ~n81299 & ~n81300;
  assign n81302 = n81209 & ~n81301;
  assign n81303 = ~n81210 & n81297;
  assign n81304 = n81210 & ~n81297;
  assign n81305 = n81295 & n81304;
  assign n81306 = ~n81210 & ~n81295;
  assign n81307 = ~n81303 & ~n81305;
  assign n81308 = ~n81306 & n81307;
  assign n81309 = ~n81209 & ~n81308;
  assign n81310 = ~n81302 & ~n81309;
  assign n81311 = P3_DATAO_REG_17_ & n78036;
  assign n81312 = ~n80914 & ~n81011;
  assign n81313 = ~n81010 & ~n81312;
  assign n81314 = ~n81310 & ~n81311;
  assign n81315 = ~n81313 & n81314;
  assign n81316 = n81310 & n81311;
  assign n81317 = ~n81314 & ~n81316;
  assign n81318 = n81313 & n81317;
  assign n81319 = ~n81315 & ~n81318;
  assign n81320 = n81311 & ~n81313;
  assign n81321 = n81310 & n81320;
  assign n81322 = n81319 & ~n81321;
  assign n81323 = n81205 & ~n81322;
  assign n81324 = ~n81205 & n81322;
  assign n81325 = ~n81323 & ~n81324;
  assign n81326 = n81204 & ~n81325;
  assign n81327 = ~n81205 & n81321;
  assign n81328 = n81205 & ~n81321;
  assign n81329 = n81319 & n81328;
  assign n81330 = ~n81205 & ~n81319;
  assign n81331 = ~n81327 & ~n81329;
  assign n81332 = ~n81330 & n81331;
  assign n81333 = ~n81204 & ~n81332;
  assign n81334 = ~n81326 & ~n81333;
  assign n81335 = P3_DATAO_REG_15_ & n77724;
  assign n81336 = n81200 & ~n81334;
  assign n81337 = n81335 & n81336;
  assign n81338 = n81200 & n81334;
  assign n81339 = ~n81335 & n81338;
  assign n81340 = ~n81337 & ~n81339;
  assign n81341 = ~n81200 & ~n81335;
  assign n81342 = ~n81334 & n81341;
  assign n81343 = ~n81200 & n81335;
  assign n81344 = n81334 & n81343;
  assign n81345 = ~n81342 & ~n81344;
  assign n81346 = n81340 & n81345;
  assign n81347 = n81198 & ~n81346;
  assign n81348 = ~n81192 & ~n81193;
  assign n81349 = ~n81043 & n81348;
  assign n81350 = ~n81037 & n81349;
  assign n81351 = ~n81196 & ~n81350;
  assign n81352 = n81346 & ~n81351;
  assign n81353 = ~n81347 & ~n81352;
  assign n81354 = P3_DATAO_REG_13_ & n77720;
  assign n81355 = n81045 & ~n81051;
  assign n81356 = ~n81052 & ~n81355;
  assign n81357 = ~n81353 & ~n81354;
  assign n81358 = ~n81356 & n81357;
  assign n81359 = n81353 & n81354;
  assign n81360 = ~n81357 & ~n81359;
  assign n81361 = n81356 & n81360;
  assign n81362 = ~n81358 & ~n81361;
  assign n81363 = n81354 & ~n81356;
  assign n81364 = n81353 & n81363;
  assign n81365 = n81362 & ~n81364;
  assign n81366 = ~n81056 & n81057;
  assign n81367 = ~n81056 & ~n81062;
  assign n81368 = P3_DATAO_REG_12_ & n77718;
  assign n81369 = ~n81069 & ~n81366;
  assign n81370 = ~n81367 & n81369;
  assign n81371 = ~n81368 & n81370;
  assign n81372 = n81368 & ~n81370;
  assign n81373 = ~n81371 & ~n81372;
  assign n81374 = n81365 & ~n81373;
  assign n81375 = ~n81365 & n81373;
  assign n81376 = ~n81374 & ~n81375;
  assign n81377 = ~n81187 & ~n81191;
  assign n81378 = ~n81376 & n81377;
  assign n81379 = n81187 & ~n81191;
  assign n81380 = n81376 & n81379;
  assign n81381 = ~n81378 & ~n81380;
  assign n81382 = n81191 & ~n81376;
  assign n81383 = n81187 & n81382;
  assign n81384 = ~n81189 & n81376;
  assign n81385 = n81190 & n81384;
  assign n81386 = ~n81187 & n81385;
  assign n81387 = ~n81383 & ~n81386;
  assign n81388 = n81381 & n81387;
  assign n81389 = n81186 & ~n81388;
  assign n81390 = ~n81186 & n81388;
  assign n81391 = ~n81389 & ~n81390;
  assign n81392 = n81185 & ~n81391;
  assign n81393 = ~n81186 & ~n81387;
  assign n81394 = ~n81186 & ~n81381;
  assign n81395 = n81186 & n81381;
  assign n81396 = n81387 & n81395;
  assign n81397 = ~n81393 & ~n81394;
  assign n81398 = ~n81396 & n81397;
  assign n81399 = ~n81185 & ~n81398;
  assign n81400 = ~n81392 & ~n81399;
  assign n81401 = P3_DATAO_REG_9_ & n77714;
  assign n81402 = ~n81400 & ~n81401;
  assign n81403 = ~n80895 & ~n81099;
  assign n81404 = ~n80894 & ~n81403;
  assign n81405 = ~n81107 & ~n81404;
  assign n81406 = n81402 & ~n81405;
  assign n81407 = n81400 & n81401;
  assign n81408 = ~n81402 & ~n81407;
  assign n81409 = n81405 & n81408;
  assign n81410 = ~n81406 & ~n81409;
  assign n81411 = n81401 & ~n81405;
  assign n81412 = n81400 & n81411;
  assign n81413 = n81410 & ~n81412;
  assign n81414 = n81181 & ~n81413;
  assign n81415 = ~n81181 & n81413;
  assign n81416 = ~n81414 & ~n81415;
  assign n81417 = n81180 & ~n81416;
  assign n81418 = ~n81181 & n81412;
  assign n81419 = n81181 & ~n81412;
  assign n81420 = n81410 & n81419;
  assign n81421 = ~n81181 & ~n81410;
  assign n81422 = ~n81418 & ~n81420;
  assign n81423 = ~n81421 & n81422;
  assign n81424 = ~n81180 & ~n81423;
  assign n81425 = ~n81417 & ~n81424;
  assign n81426 = ~n81175 & n81425;
  assign n81427 = n81175 & ~n81425;
  assign n81428 = ~n81426 & ~n81427;
  assign n81429 = P3_DATAO_REG_6_ & n77708;
  assign n81430 = ~n81428 & ~n81429;
  assign n81431 = n81428 & n81429;
  assign n81432 = ~n81135 & n81136;
  assign n81433 = ~n81135 & ~n81138;
  assign n81434 = ~n81145 & ~n81432;
  assign n81435 = ~n81433 & n81434;
  assign n81436 = ~n81430 & ~n81431;
  assign n81437 = n81435 & n81436;
  assign n81438 = ~n81435 & ~n81436;
  assign n81439 = ~n81437 & ~n81438;
  assign n81440 = P3_DATAO_REG_5_ & n77706;
  assign n81441 = ~n81439 & ~n81440;
  assign n81442 = n81439 & n81440;
  assign n81443 = ~n80880 & ~n81147;
  assign n81444 = ~n81153 & ~n81443;
  assign n81445 = ~n81157 & ~n81444;
  assign n81446 = ~n81441 & ~n81442;
  assign n81447 = n81445 & n81446;
  assign n81448 = n81441 & ~n81445;
  assign n81449 = n81440 & ~n81445;
  assign n81450 = n81439 & n81449;
  assign n81451 = ~n81447 & ~n81448;
  assign n81452 = ~n81450 & n81451;
  assign n81453 = n81167 & ~n81452;
  assign n81454 = ~n81167 & n81452;
  assign n81455 = ~n81453 & ~n81454;
  assign n81456 = n81166 & ~n81455;
  assign n81457 = n81167 & n81452;
  assign n81458 = ~n81167 & ~n81452;
  assign n81459 = ~n81457 & ~n81458;
  assign n81460 = ~n81166 & ~n81459;
  assign n81461 = ~n81456 & ~n81460;
  assign n81462 = P3_DATAO_REG_3_ & n77704;
  assign n81463 = n81461 & n81462;
  assign n81464 = ~n81461 & ~n81462;
  assign n81465 = ~n81463 & ~n81464;
  assign n81466 = P3_DATAO_REG_3_ & n80109;
  assign n81467 = P3_DATAO_REG_3_ & n77706;
  assign n81468 = ~n80380 & ~n80385;
  assign n81469 = ~n80381 & ~n81468;
  assign n81470 = n81467 & ~n81469;
  assign n81471 = n80612 & ~n80871;
  assign n81472 = ~n80612 & n80871;
  assign n81473 = ~n81471 & ~n81472;
  assign n81474 = n80876 & ~n81473;
  assign n81475 = ~n80870 & ~n80872;
  assign n81476 = ~n80876 & ~n81475;
  assign n81477 = ~n81474 & ~n81476;
  assign n81478 = n81467 & ~n81477;
  assign n81479 = ~n81469 & ~n81477;
  assign n81480 = ~n81470 & ~n81478;
  assign n81481 = ~n81479 & n81480;
  assign n81482 = n81466 & ~n81481;
  assign n81483 = n80879 & n81162;
  assign n81484 = n81466 & ~n81483;
  assign n81485 = ~n80611 & ~n81162;
  assign n81486 = ~n80878 & n81485;
  assign n81487 = n80611 & n81162;
  assign n81488 = ~n81485 & ~n81487;
  assign n81489 = n80878 & n81488;
  assign n81490 = ~n81486 & ~n81489;
  assign n81491 = n81484 & n81490;
  assign n81492 = ~n81483 & n81490;
  assign n81493 = ~n81481 & n81492;
  assign n81494 = ~n81482 & ~n81491;
  assign n81495 = ~n81493 & n81494;
  assign n81496 = ~n81465 & ~n81495;
  assign n81497 = n81465 & n81495;
  assign n81498 = ~n81496 & ~n81497;
  assign n81499 = n80610 & n81498;
  assign n81500 = ~n80610 & ~n81498;
  assign n81501 = P3_DATAO_REG_2_ & n77704;
  assign n81502 = P3_DATAO_REG_2_ & n80109;
  assign n81503 = ~n81467 & n81469;
  assign n81504 = ~n81470 & ~n81503;
  assign n81505 = n81477 & ~n81504;
  assign n81506 = ~n81477 & n81504;
  assign n81507 = ~n81505 & ~n81506;
  assign n81508 = n81502 & n81507;
  assign n81509 = ~n81502 & ~n81507;
  assign n81510 = ~n80389 & ~n80392;
  assign n81511 = ~n80395 & ~n80400;
  assign n81512 = ~n81510 & n81511;
  assign n81513 = ~n81509 & ~n81512;
  assign n81514 = ~n81508 & ~n81513;
  assign n81515 = n81501 & ~n81514;
  assign n81516 = n81466 & ~n81492;
  assign n81517 = ~n81466 & n81492;
  assign n81518 = ~n81516 & ~n81517;
  assign n81519 = n81481 & ~n81518;
  assign n81520 = ~n81466 & n81483;
  assign n81521 = ~n81466 & ~n81490;
  assign n81522 = ~n81491 & ~n81520;
  assign n81523 = ~n81521 & n81522;
  assign n81524 = ~n81481 & ~n81523;
  assign n81525 = ~n81519 & ~n81524;
  assign n81526 = n81501 & ~n81525;
  assign n81527 = ~n81514 & ~n81525;
  assign n81528 = ~n81515 & ~n81526;
  assign n81529 = ~n81527 & n81528;
  assign n81530 = ~n81500 & ~n81529;
  assign n81531 = ~n81499 & ~n81530;
  assign n81532 = n80608 & ~n81531;
  assign n81533 = ~n81461 & n81462;
  assign n81534 = n81461 & ~n81462;
  assign n81535 = ~n81495 & ~n81534;
  assign n81536 = ~n81533 & ~n81535;
  assign n81537 = P3_DATAO_REG_3_ & n80609;
  assign n81538 = P3_DATAO_REG_4_ & n77704;
  assign n81539 = ~n81166 & ~n81458;
  assign n81540 = ~n81457 & ~n81539;
  assign n81541 = ~n77706 & ~n77708;
  assign n81542 = ~n81147 & n81541;
  assign n81543 = n81153 & ~n81440;
  assign n81544 = ~n81157 & n81543;
  assign n81545 = ~n81439 & ~n81542;
  assign n81546 = ~n81544 & n81545;
  assign n81547 = ~n81449 & ~n81546;
  assign n81548 = P3_DATAO_REG_5_ & n80109;
  assign n81549 = n81168 & ~n81425;
  assign n81550 = ~n81172 & ~n81425;
  assign n81551 = ~n81173 & ~n81549;
  assign n81552 = ~n81550 & n81551;
  assign n81553 = P3_DATAO_REG_7_ & n77708;
  assign n81554 = ~n81400 & n81401;
  assign n81555 = ~n81400 & ~n81405;
  assign n81556 = ~n81411 & ~n81554;
  assign n81557 = ~n81555 & n81556;
  assign n81558 = P3_DATAO_REG_9_ & n77712;
  assign n81559 = P3_DATAO_REG_12_ & n77716;
  assign n81560 = ~n81367 & ~n81368;
  assign n81561 = ~n81069 & n81560;
  assign n81562 = ~n81366 & n81561;
  assign n81563 = n81365 & ~n81562;
  assign n81564 = ~n81372 & ~n81563;
  assign n81565 = P3_DATAO_REG_13_ & n77718;
  assign n81566 = ~n81353 & n81354;
  assign n81567 = ~n81353 & ~n81356;
  assign n81568 = ~n81363 & ~n81566;
  assign n81569 = ~n81567 & n81568;
  assign n81570 = n81565 & ~n81569;
  assign n81571 = ~n81565 & n81569;
  assign n81572 = ~n81570 & ~n81571;
  assign n81573 = ~n81334 & n81335;
  assign n81574 = ~n81200 & ~n81334;
  assign n81575 = ~n81343 & ~n81573;
  assign n81576 = ~n81574 & n81575;
  assign n81577 = P3_DATAO_REG_15_ & n77722;
  assign n81578 = ~n81310 & n81311;
  assign n81579 = ~n81310 & ~n81313;
  assign n81580 = ~n81320 & ~n81578;
  assign n81581 = ~n81579 & n81580;
  assign n81582 = P3_DATAO_REG_17_ & n77726;
  assign n81583 = ~n81260 & n81261;
  assign n81584 = ~n81260 & ~n81265;
  assign n81585 = ~n81272 & ~n81583;
  assign n81586 = ~n81584 & n81585;
  assign n81587 = P3_DATAO_REG_21_ & n77434;
  assign n81588 = P3_DATAO_REG_22_ & n77436;
  assign n81589 = ~n81218 & n81219;
  assign n81590 = ~n81218 & n81248;
  assign n81591 = ~n81256 & ~n81589;
  assign n81592 = ~n81590 & n81591;
  assign n81593 = ~n81588 & ~n81592;
  assign n81594 = ~n81236 & n81237;
  assign n81595 = ~n81236 & ~n81239;
  assign n81596 = ~n81246 & ~n81594;
  assign n81597 = ~n81595 & n81596;
  assign n81598 = P3_DATAO_REG_23_ & n77475;
  assign n81599 = P3_DATAO_REG_25_ & n77440;
  assign n81600 = P3_DATAO_REG_26_ & n77442;
  assign n81601 = P3_DATAO_REG_27_ & n77444;
  assign n81602 = n81600 & ~n81601;
  assign n81603 = ~n81600 & n81601;
  assign n81604 = ~n81602 & ~n81603;
  assign n81605 = n81599 & ~n81604;
  assign n81606 = ~n81599 & n81604;
  assign n81607 = P3_DATAO_REG_25_ & P3_DATAO_REG_26_;
  assign n81608 = n77451 & n81607;
  assign n81609 = ~n81605 & ~n81606;
  assign n81610 = ~n81608 & n81609;
  assign n81611 = n81599 & ~n81602;
  assign n81612 = ~n81599 & n81602;
  assign n81613 = ~n81611 & ~n81612;
  assign n81614 = n81608 & n81613;
  assign n81615 = ~n81610 & ~n81614;
  assign n81616 = P3_DATAO_REG_24_ & n77438;
  assign n81617 = ~n81227 & n81229;
  assign n81618 = ~n81226 & ~n81617;
  assign n81619 = ~n81615 & ~n81616;
  assign n81620 = ~n81618 & n81619;
  assign n81621 = n81615 & n81616;
  assign n81622 = ~n81619 & ~n81621;
  assign n81623 = n81618 & n81622;
  assign n81624 = ~n81620 & ~n81623;
  assign n81625 = n81616 & ~n81618;
  assign n81626 = n81615 & n81625;
  assign n81627 = n81624 & ~n81626;
  assign n81628 = n81598 & ~n81627;
  assign n81629 = ~n81598 & n81627;
  assign n81630 = ~n81628 & ~n81629;
  assign n81631 = n81597 & ~n81630;
  assign n81632 = ~n81598 & n81626;
  assign n81633 = ~n81598 & ~n81624;
  assign n81634 = n81598 & n81624;
  assign n81635 = ~n81626 & n81634;
  assign n81636 = ~n81632 & ~n81633;
  assign n81637 = ~n81635 & n81636;
  assign n81638 = ~n81597 & ~n81637;
  assign n81639 = ~n81631 & ~n81638;
  assign n81640 = n81593 & ~n81639;
  assign n81641 = n81588 & ~n81592;
  assign n81642 = n81639 & n81641;
  assign n81643 = ~n81640 & ~n81642;
  assign n81644 = n81592 & ~n81639;
  assign n81645 = n81588 & n81644;
  assign n81646 = n81592 & n81639;
  assign n81647 = ~n81588 & n81646;
  assign n81648 = ~n81645 & ~n81647;
  assign n81649 = n81643 & n81648;
  assign n81650 = n81587 & ~n81649;
  assign n81651 = ~n81587 & n81649;
  assign n81652 = ~n81650 & ~n81651;
  assign n81653 = n81586 & ~n81652;
  assign n81654 = ~n81587 & ~n81643;
  assign n81655 = n81587 & n81643;
  assign n81656 = n81648 & n81655;
  assign n81657 = ~n81587 & ~n81648;
  assign n81658 = ~n81654 & ~n81656;
  assign n81659 = ~n81657 & n81658;
  assign n81660 = ~n81586 & ~n81659;
  assign n81661 = ~n81653 & ~n81660;
  assign n81662 = P3_DATAO_REG_20_ & n77688;
  assign n81663 = ~n81214 & ~n81274;
  assign n81664 = ~n81213 & ~n81663;
  assign n81665 = ~n81281 & ~n81664;
  assign n81666 = ~n81661 & ~n81662;
  assign n81667 = ~n81665 & n81666;
  assign n81668 = n81661 & n81662;
  assign n81669 = ~n81666 & ~n81668;
  assign n81670 = n81665 & n81669;
  assign n81671 = ~n81667 & ~n81670;
  assign n81672 = n81662 & ~n81665;
  assign n81673 = n81661 & n81672;
  assign n81674 = n81671 & ~n81673;
  assign n81675 = ~n81286 & n81287;
  assign n81676 = ~n81286 & ~n81289;
  assign n81677 = P3_DATAO_REG_19_ & n77955;
  assign n81678 = ~n81296 & ~n81675;
  assign n81679 = ~n81676 & n81678;
  assign n81680 = ~n81677 & n81679;
  assign n81681 = n81677 & ~n81679;
  assign n81682 = ~n81680 & ~n81681;
  assign n81683 = n81674 & ~n81682;
  assign n81684 = ~n81674 & n81682;
  assign n81685 = ~n81683 & ~n81684;
  assign n81686 = P3_DATAO_REG_18_ & n78036;
  assign n81687 = ~n81685 & ~n81686;
  assign n81688 = ~n81210 & ~n81298;
  assign n81689 = ~n81209 & ~n81688;
  assign n81690 = ~n81305 & ~n81689;
  assign n81691 = n81687 & ~n81690;
  assign n81692 = n81685 & n81686;
  assign n81693 = ~n81687 & ~n81692;
  assign n81694 = n81690 & n81693;
  assign n81695 = ~n81691 & ~n81694;
  assign n81696 = n81686 & ~n81690;
  assign n81697 = n81685 & n81696;
  assign n81698 = n81695 & ~n81697;
  assign n81699 = n81582 & ~n81698;
  assign n81700 = ~n81582 & n81698;
  assign n81701 = ~n81699 & ~n81700;
  assign n81702 = n81581 & ~n81701;
  assign n81703 = n81582 & ~n81697;
  assign n81704 = n81695 & n81703;
  assign n81705 = ~n81582 & ~n81698;
  assign n81706 = ~n81704 & ~n81705;
  assign n81707 = ~n81581 & ~n81706;
  assign n81708 = ~n81702 & ~n81707;
  assign n81709 = P3_DATAO_REG_16_ & n77724;
  assign n81710 = ~n81708 & ~n81709;
  assign n81711 = ~n81205 & ~n81322;
  assign n81712 = ~n81204 & ~n81711;
  assign n81713 = ~n81329 & ~n81712;
  assign n81714 = n81710 & ~n81713;
  assign n81715 = ~n81708 & n81709;
  assign n81716 = n81708 & ~n81709;
  assign n81717 = ~n81715 & ~n81716;
  assign n81718 = n81713 & ~n81717;
  assign n81719 = ~n81714 & ~n81718;
  assign n81720 = n81709 & ~n81713;
  assign n81721 = n81708 & n81720;
  assign n81722 = n81719 & ~n81721;
  assign n81723 = n81577 & ~n81722;
  assign n81724 = ~n81577 & n81722;
  assign n81725 = ~n81723 & ~n81724;
  assign n81726 = n81576 & ~n81725;
  assign n81727 = n81577 & ~n81721;
  assign n81728 = n81719 & n81727;
  assign n81729 = ~n81577 & ~n81722;
  assign n81730 = ~n81728 & ~n81729;
  assign n81731 = ~n81576 & ~n81730;
  assign n81732 = ~n81726 & ~n81731;
  assign n81733 = ~n81197 & n81346;
  assign n81734 = ~n81196 & ~n81733;
  assign n81735 = P3_DATAO_REG_14_ & n77720;
  assign n81736 = ~n81732 & ~n81734;
  assign n81737 = ~n81735 & n81736;
  assign n81738 = ~n81732 & n81734;
  assign n81739 = n81735 & n81738;
  assign n81740 = ~n81734 & n81735;
  assign n81741 = n81734 & ~n81735;
  assign n81742 = ~n81740 & ~n81741;
  assign n81743 = n81732 & ~n81742;
  assign n81744 = ~n81737 & ~n81739;
  assign n81745 = ~n81743 & n81744;
  assign n81746 = n81572 & ~n81745;
  assign n81747 = ~n81572 & n81745;
  assign n81748 = ~n81746 & ~n81747;
  assign n81749 = ~n81559 & ~n81564;
  assign n81750 = ~n81748 & n81749;
  assign n81751 = n81559 & ~n81564;
  assign n81752 = ~n81559 & n81564;
  assign n81753 = ~n81751 & ~n81752;
  assign n81754 = n81748 & ~n81753;
  assign n81755 = ~n81750 & ~n81754;
  assign n81756 = n81559 & n81564;
  assign n81757 = ~n81748 & n81756;
  assign n81758 = n81755 & ~n81757;
  assign n81759 = n81187 & ~n81376;
  assign n81760 = ~n81191 & ~n81376;
  assign n81761 = P3_DATAO_REG_11_ & n78934;
  assign n81762 = ~n81379 & ~n81759;
  assign n81763 = ~n81760 & n81762;
  assign n81764 = ~n81761 & n81763;
  assign n81765 = n81761 & ~n81763;
  assign n81766 = ~n81764 & ~n81765;
  assign n81767 = n81758 & ~n81766;
  assign n81768 = ~n81758 & n81766;
  assign n81769 = ~n81767 & ~n81768;
  assign n81770 = P3_DATAO_REG_10_ & n77714;
  assign n81771 = ~n81185 & n81397;
  assign n81772 = ~n81396 & ~n81771;
  assign n81773 = ~n81769 & ~n81770;
  assign n81774 = ~n81772 & n81773;
  assign n81775 = n81769 & n81770;
  assign n81776 = ~n81773 & ~n81775;
  assign n81777 = n81772 & n81776;
  assign n81778 = ~n81774 & ~n81777;
  assign n81779 = ~n81772 & n81775;
  assign n81780 = n81778 & ~n81779;
  assign n81781 = n81558 & ~n81780;
  assign n81782 = ~n81558 & n81780;
  assign n81783 = ~n81781 & ~n81782;
  assign n81784 = n81557 & ~n81783;
  assign n81785 = ~n81558 & n81779;
  assign n81786 = ~n81558 & ~n81778;
  assign n81787 = n81558 & ~n81779;
  assign n81788 = n81778 & n81787;
  assign n81789 = ~n81785 & ~n81786;
  assign n81790 = ~n81788 & n81789;
  assign n81791 = ~n81557 & ~n81790;
  assign n81792 = ~n81784 & ~n81791;
  assign n81793 = P3_DATAO_REG_8_ & n77710;
  assign n81794 = ~n81181 & ~n81413;
  assign n81795 = ~n81180 & ~n81794;
  assign n81796 = ~n81420 & ~n81795;
  assign n81797 = ~n81792 & ~n81793;
  assign n81798 = ~n81796 & n81797;
  assign n81799 = n81792 & n81793;
  assign n81800 = ~n81797 & ~n81799;
  assign n81801 = n81796 & n81800;
  assign n81802 = ~n81798 & ~n81801;
  assign n81803 = n81793 & ~n81796;
  assign n81804 = n81792 & n81803;
  assign n81805 = n81802 & ~n81804;
  assign n81806 = n81553 & ~n81805;
  assign n81807 = ~n81553 & n81805;
  assign n81808 = ~n81806 & ~n81807;
  assign n81809 = n81552 & ~n81808;
  assign n81810 = ~n81553 & ~n81805;
  assign n81811 = n81553 & ~n81804;
  assign n81812 = n81802 & n81811;
  assign n81813 = ~n81810 & ~n81812;
  assign n81814 = ~n81552 & ~n81813;
  assign n81815 = ~n81809 & ~n81814;
  assign n81816 = P3_DATAO_REG_6_ & n77706;
  assign n81817 = ~n81430 & ~n81435;
  assign n81818 = ~n81431 & ~n81817;
  assign n81819 = ~n81815 & ~n81816;
  assign n81820 = ~n81818 & n81819;
  assign n81821 = n81815 & n81816;
  assign n81822 = ~n81819 & ~n81821;
  assign n81823 = n81818 & n81822;
  assign n81824 = ~n81820 & ~n81823;
  assign n81825 = n81816 & ~n81818;
  assign n81826 = n81815 & n81825;
  assign n81827 = n81824 & ~n81826;
  assign n81828 = n81548 & ~n81827;
  assign n81829 = ~n81548 & n81827;
  assign n81830 = ~n81828 & ~n81829;
  assign n81831 = n81547 & ~n81830;
  assign n81832 = n81548 & n81824;
  assign n81833 = ~n81826 & n81832;
  assign n81834 = ~n81548 & ~n81827;
  assign n81835 = ~n81833 & ~n81834;
  assign n81836 = ~n81547 & ~n81835;
  assign n81837 = ~n81831 & ~n81836;
  assign n81838 = ~n81538 & ~n81540;
  assign n81839 = ~n81837 & n81838;
  assign n81840 = n81538 & ~n81540;
  assign n81841 = n81837 & n81840;
  assign n81842 = ~n81839 & ~n81841;
  assign n81843 = n81540 & ~n81837;
  assign n81844 = n81538 & n81843;
  assign n81845 = n81540 & n81837;
  assign n81846 = ~n81538 & n81845;
  assign n81847 = ~n81844 & ~n81846;
  assign n81848 = n81842 & n81847;
  assign n81849 = n81537 & ~n81848;
  assign n81850 = ~n81537 & n81848;
  assign n81851 = ~n81849 & ~n81850;
  assign n81852 = n81536 & ~n81851;
  assign n81853 = ~n81537 & ~n81847;
  assign n81854 = ~n81537 & ~n81842;
  assign n81855 = n81537 & n81842;
  assign n81856 = n81847 & n81855;
  assign n81857 = ~n81853 & ~n81854;
  assign n81858 = ~n81856 & n81857;
  assign n81859 = ~n81536 & ~n81858;
  assign n81860 = ~n81852 & ~n81859;
  assign n81861 = n80608 & ~n81860;
  assign n81862 = ~n81531 & ~n81860;
  assign n81863 = ~n81532 & ~n81861;
  assign n81864 = ~n81862 & n81863;
  assign n81865 = n80606 & ~n81864;
  assign n81866 = P3_DATAO_REG_3_ & n80607;
  assign n81867 = ~n81537 & ~n81848;
  assign n81868 = ~n81536 & ~n81867;
  assign n81869 = ~n81856 & ~n81868;
  assign n81870 = n81866 & ~n81869;
  assign n81871 = n81538 & ~n81837;
  assign n81872 = ~n81540 & ~n81837;
  assign n81873 = ~n81840 & ~n81871;
  assign n81874 = ~n81872 & n81873;
  assign n81875 = P3_DATAO_REG_4_ & n80609;
  assign n81876 = ~n81815 & n81816;
  assign n81877 = ~n81815 & ~n81818;
  assign n81878 = ~n81825 & ~n81876;
  assign n81879 = ~n81877 & n81878;
  assign n81880 = P3_DATAO_REG_6_ & n80109;
  assign n81881 = P3_DATAO_REG_7_ & n77706;
  assign n81882 = ~n81552 & n81553;
  assign n81883 = ~n81552 & n81805;
  assign n81884 = ~n81812 & ~n81882;
  assign n81885 = ~n81883 & n81884;
  assign n81886 = ~n81881 & ~n81885;
  assign n81887 = ~n81792 & n81793;
  assign n81888 = ~n81792 & ~n81796;
  assign n81889 = ~n81803 & ~n81887;
  assign n81890 = ~n81888 & n81889;
  assign n81891 = P3_DATAO_REG_8_ & n77708;
  assign n81892 = ~n81760 & ~n81761;
  assign n81893 = ~n81379 & n81892;
  assign n81894 = ~n81759 & n81893;
  assign n81895 = n81758 & ~n81894;
  assign n81896 = ~n81765 & ~n81895;
  assign n81897 = P3_DATAO_REG_11_ & n77714;
  assign n81898 = n81896 & n81897;
  assign n81899 = P3_DATAO_REG_12_ & n78934;
  assign n81900 = n81559 & ~n81748;
  assign n81901 = ~n81564 & ~n81748;
  assign n81902 = ~n81751 & ~n81900;
  assign n81903 = ~n81901 & n81902;
  assign n81904 = n81899 & ~n81903;
  assign n81905 = ~n81899 & n81903;
  assign n81906 = ~n81904 & ~n81905;
  assign n81907 = ~n81732 & n81735;
  assign n81908 = ~n81740 & ~n81907;
  assign n81909 = ~n81736 & n81908;
  assign n81910 = P3_DATAO_REG_14_ & n77718;
  assign n81911 = ~n81708 & ~n81713;
  assign n81912 = ~n81715 & ~n81720;
  assign n81913 = ~n81911 & n81912;
  assign n81914 = P3_DATAO_REG_16_ & n77722;
  assign n81915 = ~n81685 & n81686;
  assign n81916 = ~n81685 & ~n81690;
  assign n81917 = ~n81696 & ~n81915;
  assign n81918 = ~n81916 & n81917;
  assign n81919 = P3_DATAO_REG_18_ & n77726;
  assign n81920 = ~n81661 & n81662;
  assign n81921 = ~n81661 & ~n81665;
  assign n81922 = ~n81672 & ~n81920;
  assign n81923 = ~n81921 & n81922;
  assign n81924 = P3_DATAO_REG_20_ & n77955;
  assign n81925 = P3_DATAO_REG_21_ & n77688;
  assign n81926 = ~n81586 & ~n81654;
  assign n81927 = ~n81657 & n81926;
  assign n81928 = ~n81656 & ~n81927;
  assign n81929 = ~n81925 & ~n81928;
  assign n81930 = n81588 & ~n81639;
  assign n81931 = ~n81592 & ~n81639;
  assign n81932 = ~n81641 & ~n81930;
  assign n81933 = ~n81931 & n81932;
  assign n81934 = P3_DATAO_REG_22_ & n77434;
  assign n81935 = P3_DATAO_REG_23_ & n77436;
  assign n81936 = ~n81615 & n81616;
  assign n81937 = ~n81615 & ~n81618;
  assign n81938 = ~n81625 & ~n81936;
  assign n81939 = ~n81937 & n81938;
  assign n81940 = P3_DATAO_REG_24_ & n77475;
  assign n81941 = P3_DATAO_REG_25_ & n77438;
  assign n81942 = ~n81606 & n81608;
  assign n81943 = ~n81605 & ~n81942;
  assign n81944 = ~n81941 & ~n81943;
  assign n81945 = P3_DATAO_REG_26_ & n77440;
  assign n81946 = P3_DATAO_REG_27_ & n77442;
  assign n81947 = P3_DATAO_REG_28_ & n77444;
  assign n81948 = n81946 & ~n81947;
  assign n81949 = ~n81946 & n81947;
  assign n81950 = ~n81948 & ~n81949;
  assign n81951 = n81945 & ~n81950;
  assign n81952 = ~n81945 & n81950;
  assign n81953 = P3_DATAO_REG_26_ & P3_DATAO_REG_27_;
  assign n81954 = n77451 & n81953;
  assign n81955 = ~n81951 & ~n81952;
  assign n81956 = ~n81954 & n81955;
  assign n81957 = ~n81945 & ~n81948;
  assign n81958 = ~n81951 & ~n81957;
  assign n81959 = n81954 & ~n81958;
  assign n81960 = ~n81956 & ~n81959;
  assign n81961 = n81944 & ~n81960;
  assign n81962 = n81941 & ~n81943;
  assign n81963 = n81960 & n81962;
  assign n81964 = n81943 & ~n81960;
  assign n81965 = n81941 & n81964;
  assign n81966 = n81943 & n81960;
  assign n81967 = ~n81941 & n81966;
  assign n81968 = ~n81961 & ~n81963;
  assign n81969 = ~n81965 & n81968;
  assign n81970 = ~n81967 & n81969;
  assign n81971 = n81940 & ~n81970;
  assign n81972 = ~n81940 & n81970;
  assign n81973 = ~n81971 & ~n81972;
  assign n81974 = n81939 & ~n81973;
  assign n81975 = n81940 & n81970;
  assign n81976 = ~n81940 & ~n81970;
  assign n81977 = ~n81975 & ~n81976;
  assign n81978 = ~n81939 & ~n81977;
  assign n81979 = ~n81974 & ~n81978;
  assign n81980 = n81935 & ~n81979;
  assign n81981 = ~n81598 & ~n81627;
  assign n81982 = ~n81597 & ~n81981;
  assign n81983 = ~n81635 & ~n81982;
  assign n81984 = n81980 & n81983;
  assign n81985 = ~n81935 & ~n81979;
  assign n81986 = ~n81983 & n81985;
  assign n81987 = ~n81984 & ~n81986;
  assign n81988 = n81935 & ~n81983;
  assign n81989 = ~n81635 & ~n81935;
  assign n81990 = ~n81982 & n81989;
  assign n81991 = ~n81988 & ~n81990;
  assign n81992 = n81979 & ~n81991;
  assign n81993 = n81987 & ~n81992;
  assign n81994 = n81934 & ~n81993;
  assign n81995 = ~n81934 & n81993;
  assign n81996 = ~n81994 & ~n81995;
  assign n81997 = n81933 & ~n81996;
  assign n81998 = n81934 & ~n81992;
  assign n81999 = n81987 & n81998;
  assign n82000 = ~n81934 & ~n81993;
  assign n82001 = ~n81999 & ~n82000;
  assign n82002 = ~n81933 & ~n82001;
  assign n82003 = ~n81997 & ~n82002;
  assign n82004 = n81929 & ~n82003;
  assign n82005 = n81925 & n81927;
  assign n82006 = ~n81925 & n81928;
  assign n82007 = n81656 & n81925;
  assign n82008 = ~n82005 & ~n82006;
  assign n82009 = ~n82007 & n82008;
  assign n82010 = n82003 & ~n82009;
  assign n82011 = ~n82004 & ~n82010;
  assign n82012 = n81925 & n81928;
  assign n82013 = ~n82003 & n82012;
  assign n82014 = n82011 & ~n82013;
  assign n82015 = n81924 & ~n82014;
  assign n82016 = ~n81924 & n82014;
  assign n82017 = ~n82015 & ~n82016;
  assign n82018 = n81923 & ~n82017;
  assign n82019 = ~n81924 & n82013;
  assign n82020 = n81924 & ~n82013;
  assign n82021 = n82011 & n82020;
  assign n82022 = ~n81924 & ~n82011;
  assign n82023 = ~n82019 & ~n82021;
  assign n82024 = ~n82022 & n82023;
  assign n82025 = ~n81923 & ~n82024;
  assign n82026 = ~n82018 & ~n82025;
  assign n82027 = P3_DATAO_REG_19_ & n78036;
  assign n82028 = n81674 & ~n81680;
  assign n82029 = ~n81681 & ~n82028;
  assign n82030 = ~n82026 & ~n82027;
  assign n82031 = ~n82029 & n82030;
  assign n82032 = n82026 & n82027;
  assign n82033 = ~n82030 & ~n82032;
  assign n82034 = n82029 & n82033;
  assign n82035 = ~n82031 & ~n82034;
  assign n82036 = n82027 & ~n82029;
  assign n82037 = n82026 & n82036;
  assign n82038 = n82035 & ~n82037;
  assign n82039 = n81919 & ~n82038;
  assign n82040 = ~n81919 & n82038;
  assign n82041 = ~n82039 & ~n82040;
  assign n82042 = n81918 & ~n82041;
  assign n82043 = ~n81919 & n82037;
  assign n82044 = n81919 & ~n82037;
  assign n82045 = n82035 & n82044;
  assign n82046 = ~n81919 & ~n82035;
  assign n82047 = ~n82043 & ~n82045;
  assign n82048 = ~n82046 & n82047;
  assign n82049 = ~n81918 & ~n82048;
  assign n82050 = ~n82042 & ~n82049;
  assign n82051 = P3_DATAO_REG_17_ & n77724;
  assign n82052 = ~n81581 & ~n81705;
  assign n82053 = ~n81704 & ~n82052;
  assign n82054 = ~n82050 & ~n82051;
  assign n82055 = ~n82053 & n82054;
  assign n82056 = n82050 & n82051;
  assign n82057 = ~n82054 & ~n82056;
  assign n82058 = n82053 & n82057;
  assign n82059 = ~n82055 & ~n82058;
  assign n82060 = n82051 & ~n82053;
  assign n82061 = n82050 & n82060;
  assign n82062 = n82059 & ~n82061;
  assign n82063 = n81914 & ~n82062;
  assign n82064 = ~n81914 & n82062;
  assign n82065 = ~n82063 & ~n82064;
  assign n82066 = n81913 & ~n82065;
  assign n82067 = ~n81914 & n82061;
  assign n82068 = n81914 & ~n82061;
  assign n82069 = n82059 & n82068;
  assign n82070 = ~n81914 & ~n82059;
  assign n82071 = ~n82067 & ~n82069;
  assign n82072 = ~n82070 & n82071;
  assign n82073 = ~n81913 & ~n82072;
  assign n82074 = ~n82066 & ~n82073;
  assign n82075 = P3_DATAO_REG_15_ & n77720;
  assign n82076 = ~n81576 & ~n81729;
  assign n82077 = ~n81728 & ~n82076;
  assign n82078 = ~n82074 & ~n82075;
  assign n82079 = ~n82077 & n82078;
  assign n82080 = n82074 & n82075;
  assign n82081 = ~n82078 & ~n82080;
  assign n82082 = n82077 & n82081;
  assign n82083 = ~n82079 & ~n82082;
  assign n82084 = n82075 & ~n82077;
  assign n82085 = n82074 & n82084;
  assign n82086 = n82083 & ~n82085;
  assign n82087 = n81910 & ~n82086;
  assign n82088 = ~n81910 & n82086;
  assign n82089 = ~n82087 & ~n82088;
  assign n82090 = n81909 & ~n82089;
  assign n82091 = ~n81910 & n82085;
  assign n82092 = n81910 & ~n82085;
  assign n82093 = n82083 & n82092;
  assign n82094 = ~n81910 & ~n82083;
  assign n82095 = ~n82091 & ~n82093;
  assign n82096 = ~n82094 & n82095;
  assign n82097 = ~n81909 & ~n82096;
  assign n82098 = ~n82090 & ~n82097;
  assign n82099 = P3_DATAO_REG_13_ & n77716;
  assign n82100 = ~n81571 & n81745;
  assign n82101 = ~n81570 & ~n82100;
  assign n82102 = ~n82098 & ~n82099;
  assign n82103 = ~n82101 & n82102;
  assign n82104 = n82098 & n82099;
  assign n82105 = ~n82102 & ~n82104;
  assign n82106 = n82101 & n82105;
  assign n82107 = ~n82103 & ~n82106;
  assign n82108 = n82099 & ~n82101;
  assign n82109 = n82098 & n82108;
  assign n82110 = n82107 & ~n82109;
  assign n82111 = n81906 & ~n82110;
  assign n82112 = ~n81899 & ~n81901;
  assign n82113 = ~n81900 & n82112;
  assign n82114 = ~n81751 & n82113;
  assign n82115 = ~n81904 & ~n82114;
  assign n82116 = n82110 & ~n82115;
  assign n82117 = ~n82111 & ~n82116;
  assign n82118 = n81898 & ~n82117;
  assign n82119 = ~n81896 & n81897;
  assign n82120 = n81896 & ~n81897;
  assign n82121 = ~n82119 & ~n82120;
  assign n82122 = n82117 & ~n82121;
  assign n82123 = ~n82118 & ~n82122;
  assign n82124 = ~n81896 & ~n81897;
  assign n82125 = ~n82117 & n82124;
  assign n82126 = n82123 & ~n82125;
  assign n82127 = n81770 & ~n81772;
  assign n82128 = ~n81769 & n81770;
  assign n82129 = ~n81769 & ~n81772;
  assign n82130 = P3_DATAO_REG_10_ & n77712;
  assign n82131 = ~n82127 & ~n82128;
  assign n82132 = ~n82129 & n82131;
  assign n82133 = ~n82130 & n82132;
  assign n82134 = n82130 & ~n82132;
  assign n82135 = ~n82133 & ~n82134;
  assign n82136 = n82126 & ~n82135;
  assign n82137 = ~n82126 & n82135;
  assign n82138 = ~n82136 & ~n82137;
  assign n82139 = P3_DATAO_REG_9_ & n77710;
  assign n82140 = ~n81558 & ~n81780;
  assign n82141 = ~n81557 & ~n82140;
  assign n82142 = ~n81788 & ~n82141;
  assign n82143 = ~n82138 & ~n82139;
  assign n82144 = ~n82142 & n82143;
  assign n82145 = n82138 & n82139;
  assign n82146 = ~n82143 & ~n82145;
  assign n82147 = n82142 & n82146;
  assign n82148 = ~n82144 & ~n82147;
  assign n82149 = ~n82142 & n82145;
  assign n82150 = n82148 & ~n82149;
  assign n82151 = n81891 & ~n82150;
  assign n82152 = ~n81891 & n82150;
  assign n82153 = ~n82151 & ~n82152;
  assign n82154 = n81890 & ~n82153;
  assign n82155 = ~n81891 & n82149;
  assign n82156 = ~n81891 & ~n82148;
  assign n82157 = n81891 & ~n82149;
  assign n82158 = n82148 & n82157;
  assign n82159 = ~n82155 & ~n82156;
  assign n82160 = ~n82158 & n82159;
  assign n82161 = ~n81890 & ~n82160;
  assign n82162 = ~n82154 & ~n82161;
  assign n82163 = n81886 & ~n82162;
  assign n82164 = n81881 & ~n81885;
  assign n82165 = n82162 & n82164;
  assign n82166 = ~n82163 & ~n82165;
  assign n82167 = n81885 & ~n82162;
  assign n82168 = n81881 & n82167;
  assign n82169 = ~n81883 & n82162;
  assign n82170 = n81884 & n82169;
  assign n82171 = ~n81881 & n82170;
  assign n82172 = ~n82168 & ~n82171;
  assign n82173 = n82166 & n82172;
  assign n82174 = n81880 & ~n82173;
  assign n82175 = ~n81880 & n82173;
  assign n82176 = ~n82174 & ~n82175;
  assign n82177 = n81879 & ~n82176;
  assign n82178 = ~n81880 & ~n82172;
  assign n82179 = ~n81880 & ~n82166;
  assign n82180 = n81880 & n82166;
  assign n82181 = n82172 & n82180;
  assign n82182 = ~n82178 & ~n82179;
  assign n82183 = ~n82181 & n82182;
  assign n82184 = ~n81879 & ~n82183;
  assign n82185 = ~n82177 & ~n82184;
  assign n82186 = P3_DATAO_REG_5_ & n77704;
  assign n82187 = ~n81547 & n81548;
  assign n82188 = ~n81547 & n81827;
  assign n82189 = ~n81833 & ~n82187;
  assign n82190 = ~n82188 & n82189;
  assign n82191 = ~n82185 & ~n82186;
  assign n82192 = ~n82190 & n82191;
  assign n82193 = n82185 & n82186;
  assign n82194 = ~n82191 & ~n82193;
  assign n82195 = n82190 & n82194;
  assign n82196 = ~n82192 & ~n82195;
  assign n82197 = n82186 & ~n82190;
  assign n82198 = n82185 & n82197;
  assign n82199 = n82196 & ~n82198;
  assign n82200 = n81875 & ~n82199;
  assign n82201 = ~n81875 & n82199;
  assign n82202 = ~n82200 & ~n82201;
  assign n82203 = n81874 & ~n82202;
  assign n82204 = n81875 & ~n82198;
  assign n82205 = n82196 & n82204;
  assign n82206 = ~n81875 & ~n82199;
  assign n82207 = ~n82205 & ~n82206;
  assign n82208 = ~n81874 & ~n82207;
  assign n82209 = ~n82203 & ~n82208;
  assign n82210 = n81870 & n82209;
  assign n82211 = n80606 & ~n82210;
  assign n82212 = ~n81866 & ~n82209;
  assign n82213 = ~n81869 & n82212;
  assign n82214 = n81866 & ~n82209;
  assign n82215 = ~n81866 & n82209;
  assign n82216 = ~n82214 & ~n82215;
  assign n82217 = n81869 & ~n82216;
  assign n82218 = ~n82213 & ~n82217;
  assign n82219 = n82211 & n82218;
  assign n82220 = ~n81864 & ~n82210;
  assign n82221 = n82218 & n82220;
  assign n82222 = ~n81865 & ~n82219;
  assign n82223 = ~n82221 & n82222;
  assign n82224 = n80604 & ~n82223;
  assign n82225 = ~n81869 & ~n82209;
  assign n82226 = ~n81870 & ~n82214;
  assign n82227 = ~n82225 & n82226;
  assign n82228 = P3_DATAO_REG_3_ & n80605;
  assign n82229 = ~n82185 & n82186;
  assign n82230 = ~n82185 & ~n82190;
  assign n82231 = ~n82197 & ~n82229;
  assign n82232 = ~n82230 & n82231;
  assign n82233 = P3_DATAO_REG_5_ & n80609;
  assign n82234 = P3_DATAO_REG_6_ & n77704;
  assign n82235 = ~n81880 & ~n82173;
  assign n82236 = ~n81879 & ~n82235;
  assign n82237 = ~n82181 & ~n82236;
  assign n82238 = ~n82234 & ~n82237;
  assign n82239 = n81881 & ~n82162;
  assign n82240 = ~n81885 & ~n82162;
  assign n82241 = ~n82164 & ~n82239;
  assign n82242 = ~n82240 & n82241;
  assign n82243 = P3_DATAO_REG_7_ & n80109;
  assign n82244 = n82139 & ~n82142;
  assign n82245 = ~n82138 & n82139;
  assign n82246 = ~n82138 & ~n82142;
  assign n82247 = ~n82244 & ~n82245;
  assign n82248 = ~n82246 & n82247;
  assign n82249 = P3_DATAO_REG_9_ & n77708;
  assign n82250 = P3_DATAO_REG_10_ & n77710;
  assign n82251 = ~n82129 & ~n82130;
  assign n82252 = ~n82127 & n82251;
  assign n82253 = ~n82128 & n82252;
  assign n82254 = n82126 & ~n82253;
  assign n82255 = ~n82134 & ~n82254;
  assign n82256 = ~n82250 & ~n82255;
  assign n82257 = P3_DATAO_REG_11_ & n77712;
  assign n82258 = n81897 & ~n82117;
  assign n82259 = ~n81896 & ~n82117;
  assign n82260 = ~n82119 & ~n82258;
  assign n82261 = ~n82259 & n82260;
  assign n82262 = n82257 & ~n82261;
  assign n82263 = ~n82257 & n82261;
  assign n82264 = ~n82098 & n82099;
  assign n82265 = ~n82098 & ~n82101;
  assign n82266 = ~n82108 & ~n82264;
  assign n82267 = ~n82265 & n82266;
  assign n82268 = P3_DATAO_REG_13_ & n78934;
  assign n82269 = ~n82074 & n82075;
  assign n82270 = ~n82074 & ~n82077;
  assign n82271 = ~n82084 & ~n82269;
  assign n82272 = ~n82270 & n82271;
  assign n82273 = P3_DATAO_REG_15_ & n77718;
  assign n82274 = ~n82050 & n82051;
  assign n82275 = ~n82050 & ~n82053;
  assign n82276 = ~n82060 & ~n82274;
  assign n82277 = ~n82275 & n82276;
  assign n82278 = P3_DATAO_REG_17_ & n77722;
  assign n82279 = P3_DATAO_REG_19_ & n77726;
  assign n82280 = ~n82026 & n82027;
  assign n82281 = ~n82026 & ~n82029;
  assign n82282 = ~n82036 & ~n82280;
  assign n82283 = ~n82281 & n82282;
  assign n82284 = n82279 & ~n82283;
  assign n82285 = ~n82279 & n82283;
  assign n82286 = ~n82284 & ~n82285;
  assign n82287 = P3_DATAO_REG_20_ & n78036;
  assign n82288 = ~n81924 & ~n82014;
  assign n82289 = ~n81923 & ~n82288;
  assign n82290 = ~n82021 & ~n82289;
  assign n82291 = ~n82287 & ~n82290;
  assign n82292 = n81925 & ~n82003;
  assign n82293 = n81925 & ~n81928;
  assign n82294 = ~n81928 & ~n82003;
  assign n82295 = ~n82292 & ~n82293;
  assign n82296 = ~n82294 & n82295;
  assign n82297 = P3_DATAO_REG_21_ & n77955;
  assign n82298 = ~n81979 & ~n81983;
  assign n82299 = ~n81980 & ~n81988;
  assign n82300 = ~n82298 & n82299;
  assign n82301 = P3_DATAO_REG_23_ & n77434;
  assign n82302 = n81941 & ~n81960;
  assign n82303 = ~n81943 & ~n81960;
  assign n82304 = ~n81962 & ~n82302;
  assign n82305 = ~n82303 & n82304;
  assign n82306 = P3_DATAO_REG_25_ & n77475;
  assign n82307 = P3_DATAO_REG_27_ & n77440;
  assign n82308 = P3_DATAO_REG_28_ & n77442;
  assign n82309 = P3_DATAO_REG_29_ & n77444;
  assign n82310 = n82308 & ~n82309;
  assign n82311 = ~n82308 & n82309;
  assign n82312 = ~n82310 & ~n82311;
  assign n82313 = n82307 & ~n82312;
  assign n82314 = ~n82307 & n82312;
  assign n82315 = P3_DATAO_REG_27_ & P3_DATAO_REG_28_;
  assign n82316 = n77451 & n82315;
  assign n82317 = ~n82313 & ~n82314;
  assign n82318 = ~n82316 & n82317;
  assign n82319 = n82307 & ~n82310;
  assign n82320 = ~n82307 & n82310;
  assign n82321 = ~n82319 & ~n82320;
  assign n82322 = n82316 & n82321;
  assign n82323 = ~n82318 & ~n82322;
  assign n82324 = P3_DATAO_REG_26_ & n77438;
  assign n82325 = ~n81952 & n81954;
  assign n82326 = ~n81951 & ~n82325;
  assign n82327 = ~n82323 & ~n82324;
  assign n82328 = ~n82326 & n82327;
  assign n82329 = n82323 & n82324;
  assign n82330 = ~n82327 & ~n82329;
  assign n82331 = n82326 & n82330;
  assign n82332 = ~n82328 & ~n82331;
  assign n82333 = n82324 & ~n82326;
  assign n82334 = n82323 & n82333;
  assign n82335 = n82332 & ~n82334;
  assign n82336 = n82306 & ~n82335;
  assign n82337 = ~n82306 & n82335;
  assign n82338 = ~n82336 & ~n82337;
  assign n82339 = n82305 & ~n82338;
  assign n82340 = ~n82306 & n82334;
  assign n82341 = ~n82306 & ~n82332;
  assign n82342 = n82306 & n82332;
  assign n82343 = ~n82334 & n82342;
  assign n82344 = ~n82340 & ~n82341;
  assign n82345 = ~n82343 & n82344;
  assign n82346 = ~n82305 & ~n82345;
  assign n82347 = ~n82339 & ~n82346;
  assign n82348 = P3_DATAO_REG_24_ & n77436;
  assign n82349 = ~n81939 & ~n81976;
  assign n82350 = ~n81975 & ~n82349;
  assign n82351 = ~n82347 & ~n82348;
  assign n82352 = ~n82350 & n82351;
  assign n82353 = n82347 & n82348;
  assign n82354 = ~n82351 & ~n82353;
  assign n82355 = n82350 & n82354;
  assign n82356 = ~n82352 & ~n82355;
  assign n82357 = n82348 & ~n82350;
  assign n82358 = n82347 & n82357;
  assign n82359 = n82356 & ~n82358;
  assign n82360 = n82301 & ~n82359;
  assign n82361 = ~n82301 & n82359;
  assign n82362 = ~n82360 & ~n82361;
  assign n82363 = n82300 & ~n82362;
  assign n82364 = ~n82301 & n82358;
  assign n82365 = n82301 & ~n82358;
  assign n82366 = n82356 & n82365;
  assign n82367 = ~n82301 & ~n82356;
  assign n82368 = ~n82364 & ~n82366;
  assign n82369 = ~n82367 & n82368;
  assign n82370 = ~n82300 & ~n82369;
  assign n82371 = ~n82363 & ~n82370;
  assign n82372 = P3_DATAO_REG_22_ & n77688;
  assign n82373 = ~n81933 & ~n82000;
  assign n82374 = ~n81999 & ~n82373;
  assign n82375 = ~n82371 & ~n82372;
  assign n82376 = ~n82374 & n82375;
  assign n82377 = ~n82371 & n82372;
  assign n82378 = n82371 & ~n82372;
  assign n82379 = ~n82377 & ~n82378;
  assign n82380 = n82374 & ~n82379;
  assign n82381 = ~n82376 & ~n82380;
  assign n82382 = n82372 & ~n82374;
  assign n82383 = n82371 & n82382;
  assign n82384 = n82381 & ~n82383;
  assign n82385 = n82297 & ~n82384;
  assign n82386 = ~n82297 & n82384;
  assign n82387 = ~n82385 & ~n82386;
  assign n82388 = n82296 & ~n82387;
  assign n82389 = n82297 & ~n82383;
  assign n82390 = n82381 & n82389;
  assign n82391 = ~n82297 & ~n82384;
  assign n82392 = ~n82390 & ~n82391;
  assign n82393 = ~n82296 & ~n82392;
  assign n82394 = ~n82388 & ~n82393;
  assign n82395 = n82291 & ~n82394;
  assign n82396 = n82287 & ~n82290;
  assign n82397 = n82394 & n82396;
  assign n82398 = n82290 & ~n82394;
  assign n82399 = n82287 & n82398;
  assign n82400 = n82290 & n82394;
  assign n82401 = ~n82287 & n82400;
  assign n82402 = ~n82395 & ~n82397;
  assign n82403 = ~n82399 & n82402;
  assign n82404 = ~n82401 & n82403;
  assign n82405 = n82286 & ~n82404;
  assign n82406 = ~n82279 & ~n82281;
  assign n82407 = ~n82036 & n82406;
  assign n82408 = ~n82280 & n82407;
  assign n82409 = ~n82284 & ~n82408;
  assign n82410 = n82404 & ~n82409;
  assign n82411 = ~n82405 & ~n82410;
  assign n82412 = P3_DATAO_REG_18_ & n77724;
  assign n82413 = ~n81919 & ~n82038;
  assign n82414 = ~n81918 & ~n82413;
  assign n82415 = ~n82045 & ~n82414;
  assign n82416 = ~n82411 & ~n82412;
  assign n82417 = ~n82415 & n82416;
  assign n82418 = n82411 & n82412;
  assign n82419 = ~n82416 & ~n82418;
  assign n82420 = n82415 & n82419;
  assign n82421 = ~n82417 & ~n82420;
  assign n82422 = n82412 & ~n82415;
  assign n82423 = n82411 & n82422;
  assign n82424 = n82421 & ~n82423;
  assign n82425 = n82278 & ~n82424;
  assign n82426 = ~n82278 & n82424;
  assign n82427 = ~n82425 & ~n82426;
  assign n82428 = n82277 & ~n82427;
  assign n82429 = ~n82278 & n82423;
  assign n82430 = n82278 & ~n82423;
  assign n82431 = n82421 & n82430;
  assign n82432 = ~n82278 & ~n82421;
  assign n82433 = ~n82429 & ~n82431;
  assign n82434 = ~n82432 & n82433;
  assign n82435 = ~n82277 & ~n82434;
  assign n82436 = ~n82428 & ~n82435;
  assign n82437 = P3_DATAO_REG_16_ & n77720;
  assign n82438 = ~n81914 & ~n82062;
  assign n82439 = ~n81913 & ~n82438;
  assign n82440 = ~n82069 & ~n82439;
  assign n82441 = ~n82436 & ~n82437;
  assign n82442 = ~n82440 & n82441;
  assign n82443 = n82436 & n82437;
  assign n82444 = ~n82441 & ~n82443;
  assign n82445 = n82440 & n82444;
  assign n82446 = ~n82442 & ~n82445;
  assign n82447 = n82437 & ~n82440;
  assign n82448 = n82436 & n82447;
  assign n82449 = n82446 & ~n82448;
  assign n82450 = n82273 & ~n82449;
  assign n82451 = ~n82273 & n82449;
  assign n82452 = ~n82450 & ~n82451;
  assign n82453 = n82272 & ~n82452;
  assign n82454 = ~n82273 & n82448;
  assign n82455 = n82273 & ~n82448;
  assign n82456 = n82446 & n82455;
  assign n82457 = ~n82273 & ~n82446;
  assign n82458 = ~n82454 & ~n82456;
  assign n82459 = ~n82457 & n82458;
  assign n82460 = ~n82272 & ~n82459;
  assign n82461 = ~n82453 & ~n82460;
  assign n82462 = P3_DATAO_REG_14_ & n77716;
  assign n82463 = ~n81910 & ~n82086;
  assign n82464 = ~n81909 & ~n82463;
  assign n82465 = ~n82093 & ~n82464;
  assign n82466 = ~n82461 & ~n82462;
  assign n82467 = ~n82465 & n82466;
  assign n82468 = n82461 & n82462;
  assign n82469 = ~n82466 & ~n82468;
  assign n82470 = n82465 & n82469;
  assign n82471 = ~n82467 & ~n82470;
  assign n82472 = n82462 & ~n82465;
  assign n82473 = n82461 & n82472;
  assign n82474 = n82471 & ~n82473;
  assign n82475 = n82268 & ~n82474;
  assign n82476 = ~n82268 & n82474;
  assign n82477 = ~n82475 & ~n82476;
  assign n82478 = n82267 & ~n82477;
  assign n82479 = ~n82268 & n82473;
  assign n82480 = n82268 & ~n82473;
  assign n82481 = n82471 & n82480;
  assign n82482 = ~n82268 & ~n82471;
  assign n82483 = ~n82479 & ~n82481;
  assign n82484 = ~n82482 & n82483;
  assign n82485 = ~n82267 & ~n82484;
  assign n82486 = ~n82478 & ~n82485;
  assign n82487 = ~n81905 & n82110;
  assign n82488 = ~n81904 & ~n82487;
  assign n82489 = P3_DATAO_REG_12_ & n77714;
  assign n82490 = ~n82486 & ~n82488;
  assign n82491 = ~n82489 & n82490;
  assign n82492 = ~n82486 & n82488;
  assign n82493 = n82489 & n82492;
  assign n82494 = ~n82488 & n82489;
  assign n82495 = n82488 & ~n82489;
  assign n82496 = ~n82494 & ~n82495;
  assign n82497 = n82486 & ~n82496;
  assign n82498 = ~n82491 & ~n82493;
  assign n82499 = ~n82497 & n82498;
  assign n82500 = ~n82262 & ~n82263;
  assign n82501 = ~n82499 & n82500;
  assign n82502 = ~n82257 & ~n82259;
  assign n82503 = ~n82258 & n82502;
  assign n82504 = ~n82119 & n82503;
  assign n82505 = ~n82262 & ~n82504;
  assign n82506 = n82499 & ~n82505;
  assign n82507 = ~n82501 & ~n82506;
  assign n82508 = n82256 & ~n82507;
  assign n82509 = n82250 & ~n82255;
  assign n82510 = ~n82250 & n82255;
  assign n82511 = ~n82509 & ~n82510;
  assign n82512 = n82507 & ~n82511;
  assign n82513 = ~n82508 & ~n82512;
  assign n82514 = n82250 & n82255;
  assign n82515 = ~n82507 & n82514;
  assign n82516 = n82513 & ~n82515;
  assign n82517 = n82249 & ~n82516;
  assign n82518 = ~n82249 & n82516;
  assign n82519 = ~n82517 & ~n82518;
  assign n82520 = n82248 & ~n82519;
  assign n82521 = ~n82249 & ~n82507;
  assign n82522 = n82514 & n82521;
  assign n82523 = n82249 & ~n82515;
  assign n82524 = n82513 & n82523;
  assign n82525 = ~n82249 & ~n82513;
  assign n82526 = ~n82522 & ~n82524;
  assign n82527 = ~n82525 & n82526;
  assign n82528 = ~n82248 & ~n82527;
  assign n82529 = ~n82520 & ~n82528;
  assign n82530 = P3_DATAO_REG_8_ & n77706;
  assign n82531 = ~n81891 & ~n82150;
  assign n82532 = ~n81890 & ~n82531;
  assign n82533 = ~n82158 & ~n82532;
  assign n82534 = ~n82529 & ~n82530;
  assign n82535 = ~n82533 & n82534;
  assign n82536 = n82529 & n82530;
  assign n82537 = ~n82534 & ~n82536;
  assign n82538 = n82533 & n82537;
  assign n82539 = ~n82535 & ~n82538;
  assign n82540 = n82530 & ~n82533;
  assign n82541 = n82529 & n82540;
  assign n82542 = n82539 & ~n82541;
  assign n82543 = n82243 & ~n82542;
  assign n82544 = ~n82243 & n82542;
  assign n82545 = ~n82543 & ~n82544;
  assign n82546 = n82242 & ~n82545;
  assign n82547 = ~n82243 & n82541;
  assign n82548 = n82243 & ~n82541;
  assign n82549 = n82539 & n82548;
  assign n82550 = ~n82243 & ~n82539;
  assign n82551 = ~n82547 & ~n82549;
  assign n82552 = ~n82550 & n82551;
  assign n82553 = ~n82242 & ~n82552;
  assign n82554 = ~n82546 & ~n82553;
  assign n82555 = n82238 & ~n82554;
  assign n82556 = n82234 & n82236;
  assign n82557 = ~n82234 & n82237;
  assign n82558 = n82181 & n82234;
  assign n82559 = ~n82556 & ~n82557;
  assign n82560 = ~n82558 & n82559;
  assign n82561 = n82554 & ~n82560;
  assign n82562 = ~n82555 & ~n82561;
  assign n82563 = n82234 & n82237;
  assign n82564 = ~n82554 & n82563;
  assign n82565 = n82562 & ~n82564;
  assign n82566 = n82233 & ~n82565;
  assign n82567 = ~n82233 & n82565;
  assign n82568 = ~n82566 & ~n82567;
  assign n82569 = n82232 & ~n82568;
  assign n82570 = ~n82233 & ~n82554;
  assign n82571 = n82563 & n82570;
  assign n82572 = n82233 & ~n82564;
  assign n82573 = n82562 & n82572;
  assign n82574 = ~n82233 & ~n82562;
  assign n82575 = ~n82571 & ~n82573;
  assign n82576 = ~n82574 & n82575;
  assign n82577 = ~n82232 & ~n82576;
  assign n82578 = ~n82569 & ~n82577;
  assign n82579 = P3_DATAO_REG_4_ & n80607;
  assign n82580 = ~n81874 & ~n82206;
  assign n82581 = ~n82205 & ~n82580;
  assign n82582 = ~n82578 & ~n82579;
  assign n82583 = ~n82581 & n82582;
  assign n82584 = n82578 & n82579;
  assign n82585 = ~n82582 & ~n82584;
  assign n82586 = n82581 & n82585;
  assign n82587 = ~n82583 & ~n82586;
  assign n82588 = n82579 & ~n82581;
  assign n82589 = n82578 & n82588;
  assign n82590 = n82587 & ~n82589;
  assign n82591 = n82228 & ~n82590;
  assign n82592 = ~n82228 & n82590;
  assign n82593 = ~n82591 & ~n82592;
  assign n82594 = n82227 & ~n82593;
  assign n82595 = ~n82228 & n82589;
  assign n82596 = n82228 & ~n82589;
  assign n82597 = n82587 & n82596;
  assign n82598 = ~n82228 & ~n82587;
  assign n82599 = ~n82595 & ~n82597;
  assign n82600 = ~n82598 & n82599;
  assign n82601 = ~n82227 & ~n82600;
  assign n82602 = ~n82594 & ~n82601;
  assign n82603 = n82224 & n82602;
  assign n82604 = n80602 & ~n82603;
  assign n82605 = ~n80604 & ~n82602;
  assign n82606 = ~n82223 & n82605;
  assign n82607 = n80604 & n82602;
  assign n82608 = ~n82605 & ~n82607;
  assign n82609 = n82223 & n82608;
  assign n82610 = ~n82606 & ~n82609;
  assign n82611 = n82604 & n82610;
  assign n82612 = ~n82603 & n82610;
  assign n82613 = ~n80602 & ~n82612;
  assign n82614 = P3_DATAO_REG_1_ & n80603;
  assign n82615 = P3_DATAO_REG_1_ & n80607;
  assign n82616 = P3_DATAO_REG_1_ & n80609;
  assign n82617 = ~n81508 & ~n81509;
  assign n82618 = ~n81512 & ~n82617;
  assign n82619 = n81512 & n82617;
  assign n82620 = ~n82618 & ~n82619;
  assign n82621 = ~n77704 & ~n80109;
  assign n82622 = ~n80402 & n82621;
  assign n82623 = P3_DATAO_REG_1_ & n77704;
  assign n82624 = ~n80407 & ~n82623;
  assign n82625 = n80108 & n82624;
  assign n82626 = ~n82620 & ~n82622;
  assign n82627 = ~n82625 & n82626;
  assign n82628 = ~n80110 & ~n80402;
  assign n82629 = ~n80108 & ~n82628;
  assign n82630 = ~n80407 & ~n82629;
  assign n82631 = n82623 & ~n82630;
  assign n82632 = ~n82627 & ~n82631;
  assign n82633 = n82616 & ~n82632;
  assign n82634 = ~n81501 & n81514;
  assign n82635 = ~n81515 & ~n82634;
  assign n82636 = n81525 & ~n82635;
  assign n82637 = ~n81525 & n82635;
  assign n82638 = ~n82636 & ~n82637;
  assign n82639 = ~n82616 & n82632;
  assign n82640 = n82638 & ~n82639;
  assign n82641 = ~n82633 & ~n82640;
  assign n82642 = n82615 & ~n82641;
  assign n82643 = ~n81499 & ~n81500;
  assign n82644 = n81529 & n82643;
  assign n82645 = ~n81529 & ~n82643;
  assign n82646 = ~n82644 & ~n82645;
  assign n82647 = n82615 & ~n82646;
  assign n82648 = ~n82641 & ~n82646;
  assign n82649 = ~n82642 & ~n82647;
  assign n82650 = ~n82648 & n82649;
  assign n82651 = n80608 & ~n81499;
  assign n82652 = ~n81530 & n82651;
  assign n82653 = ~n81860 & n82652;
  assign n82654 = n81532 & n81860;
  assign n82655 = ~n82653 & ~n82654;
  assign n82656 = ~n80608 & ~n81531;
  assign n82657 = ~n81860 & n82656;
  assign n82658 = ~n80608 & ~n81499;
  assign n82659 = ~n81530 & n82658;
  assign n82660 = n81860 & n82659;
  assign n82661 = ~n82657 & ~n82660;
  assign n82662 = n82655 & n82661;
  assign n82663 = P3_DATAO_REG_1_ & n80605;
  assign n82664 = n82662 & n82663;
  assign n82665 = ~n82614 & n82650;
  assign n82666 = ~n82664 & n82665;
  assign n82667 = ~n80603 & ~n80605;
  assign n82668 = ~n82662 & n82667;
  assign n82669 = ~n82666 & ~n82668;
  assign n82670 = ~n82210 & n82218;
  assign n82671 = n80606 & ~n82670;
  assign n82672 = ~n80606 & n82670;
  assign n82673 = ~n82671 & ~n82672;
  assign n82674 = n81864 & ~n82673;
  assign n82675 = ~n80606 & ~n82670;
  assign n82676 = ~n82219 & ~n82675;
  assign n82677 = ~n81864 & ~n82676;
  assign n82678 = ~n82674 & ~n82677;
  assign n82679 = n82669 & ~n82678;
  assign n82680 = ~n82655 & ~n82663;
  assign n82681 = ~n82661 & ~n82663;
  assign n82682 = ~n82650 & ~n82680;
  assign n82683 = ~n82681 & n82682;
  assign n82684 = ~n82664 & ~n82683;
  assign n82685 = n82614 & ~n82684;
  assign n82686 = ~n82679 & ~n82685;
  assign n82687 = ~n82613 & ~n82686;
  assign n82688 = ~n82611 & ~n82687;
  assign n82689 = n80600 & ~n82688;
  assign n82690 = n80604 & ~n82602;
  assign n82691 = ~n82223 & ~n82602;
  assign n82692 = ~n82224 & ~n82690;
  assign n82693 = ~n82691 & n82692;
  assign n82694 = P3_DATAO_REG_2_ & n80601;
  assign n82695 = ~n82578 & n82579;
  assign n82696 = ~n82578 & ~n82581;
  assign n82697 = ~n82588 & ~n82695;
  assign n82698 = ~n82696 & n82697;
  assign n82699 = P3_DATAO_REG_4_ & n80605;
  assign n82700 = P3_DATAO_REG_5_ & n80607;
  assign n82701 = ~n82571 & ~n82574;
  assign n82702 = ~n82232 & n82701;
  assign n82703 = ~n82573 & ~n82702;
  assign n82704 = ~n82700 & ~n82703;
  assign n82705 = P3_DATAO_REG_6_ & n80609;
  assign n82706 = n82234 & ~n82554;
  assign n82707 = n82234 & ~n82237;
  assign n82708 = ~n82237 & ~n82554;
  assign n82709 = ~n82706 & ~n82707;
  assign n82710 = ~n82708 & n82709;
  assign n82711 = n82705 & ~n82710;
  assign n82712 = ~n82705 & n82710;
  assign n82713 = ~n82711 & ~n82712;
  assign n82714 = P3_DATAO_REG_7_ & n77704;
  assign n82715 = ~n82243 & ~n82542;
  assign n82716 = ~n82242 & ~n82715;
  assign n82717 = ~n82549 & ~n82716;
  assign n82718 = ~n82714 & ~n82717;
  assign n82719 = P3_DATAO_REG_8_ & n80109;
  assign n82720 = ~n82529 & n82530;
  assign n82721 = ~n82529 & ~n82533;
  assign n82722 = ~n82540 & ~n82720;
  assign n82723 = ~n82721 & n82722;
  assign n82724 = n82719 & ~n82723;
  assign n82725 = ~n82719 & n82723;
  assign n82726 = ~n82724 & ~n82725;
  assign n82727 = ~n82249 & ~n82516;
  assign n82728 = ~n82248 & ~n82727;
  assign n82729 = ~n82524 & ~n82728;
  assign n82730 = P3_DATAO_REG_9_ & n77706;
  assign n82731 = n82729 & n82730;
  assign n82732 = n82250 & ~n82507;
  assign n82733 = ~n82255 & ~n82507;
  assign n82734 = ~n82509 & ~n82732;
  assign n82735 = ~n82733 & n82734;
  assign n82736 = P3_DATAO_REG_10_ & n77708;
  assign n82737 = ~n82486 & n82489;
  assign n82738 = ~n82494 & ~n82737;
  assign n82739 = ~n82490 & n82738;
  assign n82740 = P3_DATAO_REG_12_ & n77712;
  assign n82741 = ~n82461 & n82462;
  assign n82742 = ~n82461 & ~n82465;
  assign n82743 = ~n82472 & ~n82741;
  assign n82744 = ~n82742 & n82743;
  assign n82745 = P3_DATAO_REG_14_ & n78934;
  assign n82746 = ~n82436 & n82437;
  assign n82747 = ~n82436 & ~n82440;
  assign n82748 = ~n82447 & ~n82746;
  assign n82749 = ~n82747 & n82748;
  assign n82750 = P3_DATAO_REG_16_ & n77718;
  assign n82751 = ~n82411 & n82412;
  assign n82752 = ~n82411 & ~n82415;
  assign n82753 = ~n82422 & ~n82751;
  assign n82754 = ~n82752 & n82753;
  assign n82755 = P3_DATAO_REG_18_ & n77722;
  assign n82756 = n82287 & ~n82394;
  assign n82757 = ~n82290 & ~n82394;
  assign n82758 = ~n82396 & ~n82756;
  assign n82759 = ~n82757 & n82758;
  assign n82760 = P3_DATAO_REG_20_ & n77726;
  assign n82761 = ~n82371 & ~n82374;
  assign n82762 = ~n82377 & ~n82382;
  assign n82763 = ~n82761 & n82762;
  assign n82764 = P3_DATAO_REG_22_ & n77955;
  assign n82765 = ~n82347 & n82348;
  assign n82766 = ~n82347 & ~n82350;
  assign n82767 = ~n82357 & ~n82765;
  assign n82768 = ~n82766 & n82767;
  assign n82769 = P3_DATAO_REG_24_ & n77434;
  assign n82770 = ~n82323 & n82324;
  assign n82771 = ~n82323 & ~n82326;
  assign n82772 = ~n82333 & ~n82770;
  assign n82773 = ~n82771 & n82772;
  assign n82774 = P3_DATAO_REG_26_ & n77475;
  assign n82775 = P3_DATAO_REG_28_ & n77440;
  assign n82776 = P3_DATAO_REG_29_ & n77442;
  assign n82777 = P3_DATAO_REG_30_ & n77444;
  assign n82778 = n82776 & ~n82777;
  assign n82779 = ~n82776 & n82777;
  assign n82780 = ~n82778 & ~n82779;
  assign n82781 = n82775 & ~n82780;
  assign n82782 = ~n82775 & n82780;
  assign n82783 = P3_DATAO_REG_28_ & P3_DATAO_REG_29_;
  assign n82784 = n77451 & n82783;
  assign n82785 = ~n82781 & ~n82782;
  assign n82786 = ~n82784 & n82785;
  assign n82787 = ~n82775 & ~n82778;
  assign n82788 = n82775 & ~n82777;
  assign n82789 = ~n82787 & ~n82788;
  assign n82790 = n82784 & ~n82789;
  assign n82791 = ~n82786 & ~n82790;
  assign n82792 = P3_DATAO_REG_27_ & n77438;
  assign n82793 = ~n82314 & n82316;
  assign n82794 = ~n82313 & ~n82793;
  assign n82795 = ~n82791 & ~n82792;
  assign n82796 = ~n82794 & n82795;
  assign n82797 = n82791 & n82792;
  assign n82798 = ~n82795 & ~n82797;
  assign n82799 = n82794 & n82798;
  assign n82800 = ~n82796 & ~n82799;
  assign n82801 = n82792 & ~n82794;
  assign n82802 = n82791 & n82801;
  assign n82803 = n82800 & ~n82802;
  assign n82804 = n82774 & ~n82803;
  assign n82805 = ~n82774 & n82803;
  assign n82806 = ~n82804 & ~n82805;
  assign n82807 = n82773 & ~n82806;
  assign n82808 = ~n82774 & n82802;
  assign n82809 = ~n82774 & ~n82800;
  assign n82810 = n82774 & n82800;
  assign n82811 = ~n82802 & n82810;
  assign n82812 = ~n82808 & ~n82809;
  assign n82813 = ~n82811 & n82812;
  assign n82814 = ~n82773 & ~n82813;
  assign n82815 = ~n82807 & ~n82814;
  assign n82816 = P3_DATAO_REG_25_ & n77436;
  assign n82817 = ~n82306 & ~n82335;
  assign n82818 = ~n82305 & ~n82817;
  assign n82819 = ~n82343 & ~n82818;
  assign n82820 = ~n82815 & ~n82816;
  assign n82821 = ~n82819 & n82820;
  assign n82822 = n82815 & n82816;
  assign n82823 = ~n82820 & ~n82822;
  assign n82824 = n82819 & n82823;
  assign n82825 = ~n82821 & ~n82824;
  assign n82826 = n82816 & ~n82819;
  assign n82827 = n82815 & n82826;
  assign n82828 = n82825 & ~n82827;
  assign n82829 = n82769 & ~n82828;
  assign n82830 = ~n82769 & n82828;
  assign n82831 = ~n82829 & ~n82830;
  assign n82832 = n82768 & ~n82831;
  assign n82833 = ~n82769 & n82827;
  assign n82834 = n82769 & ~n82827;
  assign n82835 = n82825 & n82834;
  assign n82836 = ~n82769 & ~n82825;
  assign n82837 = ~n82833 & ~n82835;
  assign n82838 = ~n82836 & n82837;
  assign n82839 = ~n82768 & ~n82838;
  assign n82840 = ~n82832 & ~n82839;
  assign n82841 = P3_DATAO_REG_23_ & n77688;
  assign n82842 = ~n82301 & ~n82359;
  assign n82843 = ~n82300 & ~n82842;
  assign n82844 = ~n82366 & ~n82843;
  assign n82845 = ~n82840 & ~n82841;
  assign n82846 = ~n82844 & n82845;
  assign n82847 = n82840 & n82841;
  assign n82848 = ~n82845 & ~n82847;
  assign n82849 = n82844 & n82848;
  assign n82850 = ~n82846 & ~n82849;
  assign n82851 = n82841 & ~n82844;
  assign n82852 = n82840 & n82851;
  assign n82853 = n82850 & ~n82852;
  assign n82854 = n82764 & ~n82853;
  assign n82855 = ~n82764 & n82853;
  assign n82856 = ~n82854 & ~n82855;
  assign n82857 = n82763 & ~n82856;
  assign n82858 = ~n82764 & n82852;
  assign n82859 = n82764 & ~n82852;
  assign n82860 = n82850 & n82859;
  assign n82861 = ~n82764 & ~n82850;
  assign n82862 = ~n82858 & ~n82860;
  assign n82863 = ~n82861 & n82862;
  assign n82864 = ~n82763 & ~n82863;
  assign n82865 = ~n82857 & ~n82864;
  assign n82866 = P3_DATAO_REG_21_ & n78036;
  assign n82867 = ~n82296 & ~n82391;
  assign n82868 = ~n82390 & ~n82867;
  assign n82869 = ~n82865 & ~n82866;
  assign n82870 = ~n82868 & n82869;
  assign n82871 = n82865 & n82866;
  assign n82872 = ~n82869 & ~n82871;
  assign n82873 = n82868 & n82872;
  assign n82874 = ~n82870 & ~n82873;
  assign n82875 = n82866 & ~n82868;
  assign n82876 = n82865 & n82875;
  assign n82877 = n82874 & ~n82876;
  assign n82878 = n82760 & ~n82877;
  assign n82879 = ~n82760 & n82877;
  assign n82880 = ~n82878 & ~n82879;
  assign n82881 = n82759 & ~n82880;
  assign n82882 = ~n82760 & n82876;
  assign n82883 = ~n82760 & ~n82874;
  assign n82884 = n82760 & ~n82876;
  assign n82885 = n82874 & n82884;
  assign n82886 = ~n82882 & ~n82883;
  assign n82887 = ~n82885 & n82886;
  assign n82888 = ~n82759 & ~n82887;
  assign n82889 = ~n82881 & ~n82888;
  assign n82890 = P3_DATAO_REG_19_ & n77724;
  assign n82891 = ~n82285 & n82404;
  assign n82892 = ~n82284 & ~n82891;
  assign n82893 = ~n82889 & ~n82890;
  assign n82894 = ~n82892 & n82893;
  assign n82895 = n82889 & n82890;
  assign n82896 = ~n82893 & ~n82895;
  assign n82897 = n82892 & n82896;
  assign n82898 = ~n82894 & ~n82897;
  assign n82899 = n82890 & ~n82892;
  assign n82900 = n82889 & n82899;
  assign n82901 = n82898 & ~n82900;
  assign n82902 = n82755 & ~n82901;
  assign n82903 = ~n82755 & n82901;
  assign n82904 = ~n82902 & ~n82903;
  assign n82905 = n82754 & ~n82904;
  assign n82906 = ~n82755 & n82900;
  assign n82907 = ~n82755 & ~n82898;
  assign n82908 = n82755 & ~n82900;
  assign n82909 = n82898 & n82908;
  assign n82910 = ~n82906 & ~n82907;
  assign n82911 = ~n82909 & n82910;
  assign n82912 = ~n82754 & ~n82911;
  assign n82913 = ~n82905 & ~n82912;
  assign n82914 = P3_DATAO_REG_17_ & n77720;
  assign n82915 = ~n82278 & ~n82424;
  assign n82916 = ~n82277 & ~n82915;
  assign n82917 = ~n82431 & ~n82916;
  assign n82918 = ~n82913 & ~n82914;
  assign n82919 = ~n82917 & n82918;
  assign n82920 = n82913 & n82914;
  assign n82921 = ~n82918 & ~n82920;
  assign n82922 = n82917 & n82921;
  assign n82923 = ~n82919 & ~n82922;
  assign n82924 = n82914 & ~n82917;
  assign n82925 = n82913 & n82924;
  assign n82926 = n82923 & ~n82925;
  assign n82927 = n82750 & ~n82926;
  assign n82928 = ~n82750 & n82926;
  assign n82929 = ~n82927 & ~n82928;
  assign n82930 = n82749 & ~n82929;
  assign n82931 = ~n82750 & n82925;
  assign n82932 = n82750 & ~n82925;
  assign n82933 = n82923 & n82932;
  assign n82934 = ~n82750 & ~n82923;
  assign n82935 = ~n82931 & ~n82933;
  assign n82936 = ~n82934 & n82935;
  assign n82937 = ~n82749 & ~n82936;
  assign n82938 = ~n82930 & ~n82937;
  assign n82939 = P3_DATAO_REG_15_ & n77716;
  assign n82940 = ~n82273 & ~n82449;
  assign n82941 = ~n82272 & ~n82940;
  assign n82942 = ~n82456 & ~n82941;
  assign n82943 = ~n82938 & ~n82939;
  assign n82944 = ~n82942 & n82943;
  assign n82945 = n82938 & n82939;
  assign n82946 = ~n82943 & ~n82945;
  assign n82947 = n82942 & n82946;
  assign n82948 = ~n82944 & ~n82947;
  assign n82949 = n82939 & ~n82942;
  assign n82950 = n82938 & n82949;
  assign n82951 = n82948 & ~n82950;
  assign n82952 = n82745 & ~n82951;
  assign n82953 = ~n82745 & n82951;
  assign n82954 = ~n82952 & ~n82953;
  assign n82955 = n82744 & ~n82954;
  assign n82956 = ~n82745 & n82950;
  assign n82957 = n82745 & ~n82950;
  assign n82958 = n82948 & n82957;
  assign n82959 = ~n82745 & ~n82948;
  assign n82960 = ~n82956 & ~n82958;
  assign n82961 = ~n82959 & n82960;
  assign n82962 = ~n82744 & ~n82961;
  assign n82963 = ~n82955 & ~n82962;
  assign n82964 = P3_DATAO_REG_13_ & n77714;
  assign n82965 = ~n82268 & ~n82474;
  assign n82966 = ~n82267 & ~n82965;
  assign n82967 = ~n82481 & ~n82966;
  assign n82968 = ~n82963 & ~n82964;
  assign n82969 = ~n82967 & n82968;
  assign n82970 = n82963 & n82964;
  assign n82971 = ~n82968 & ~n82970;
  assign n82972 = n82967 & n82971;
  assign n82973 = ~n82969 & ~n82972;
  assign n82974 = n82964 & ~n82967;
  assign n82975 = n82963 & n82974;
  assign n82976 = n82973 & ~n82975;
  assign n82977 = n82740 & ~n82976;
  assign n82978 = ~n82740 & n82976;
  assign n82979 = ~n82977 & ~n82978;
  assign n82980 = n82739 & ~n82979;
  assign n82981 = ~n82740 & n82975;
  assign n82982 = n82740 & ~n82975;
  assign n82983 = n82973 & n82982;
  assign n82984 = ~n82740 & ~n82973;
  assign n82985 = ~n82981 & ~n82983;
  assign n82986 = ~n82984 & n82985;
  assign n82987 = ~n82739 & ~n82986;
  assign n82988 = ~n82980 & ~n82987;
  assign n82989 = P3_DATAO_REG_11_ & n77710;
  assign n82990 = ~n82263 & n82499;
  assign n82991 = ~n82262 & ~n82990;
  assign n82992 = ~n82988 & ~n82989;
  assign n82993 = ~n82991 & n82992;
  assign n82994 = n82988 & n82989;
  assign n82995 = ~n82992 & ~n82994;
  assign n82996 = n82991 & n82995;
  assign n82997 = ~n82993 & ~n82996;
  assign n82998 = n82989 & ~n82991;
  assign n82999 = n82988 & n82998;
  assign n83000 = n82997 & ~n82999;
  assign n83001 = n82736 & ~n83000;
  assign n83002 = ~n82736 & n83000;
  assign n83003 = ~n83001 & ~n83002;
  assign n83004 = n82735 & ~n83003;
  assign n83005 = ~n82736 & n82999;
  assign n83006 = n82736 & ~n82999;
  assign n83007 = n82997 & n83006;
  assign n83008 = ~n82736 & ~n82997;
  assign n83009 = ~n83005 & ~n83007;
  assign n83010 = ~n83008 & n83009;
  assign n83011 = ~n82735 & ~n83010;
  assign n83012 = ~n83004 & ~n83011;
  assign n83013 = n82731 & ~n83012;
  assign n83014 = ~n82729 & n82730;
  assign n83015 = n82729 & ~n82730;
  assign n83016 = ~n83014 & ~n83015;
  assign n83017 = n83012 & ~n83016;
  assign n83018 = ~n83013 & ~n83017;
  assign n83019 = ~n82729 & ~n82730;
  assign n83020 = ~n83012 & n83019;
  assign n83021 = n83018 & ~n83020;
  assign n83022 = n82726 & ~n83021;
  assign n83023 = ~n82726 & n83021;
  assign n83024 = ~n83022 & ~n83023;
  assign n83025 = n82718 & ~n83024;
  assign n83026 = n82714 & ~n82717;
  assign n83027 = n83024 & n83026;
  assign n83028 = n82717 & ~n83024;
  assign n83029 = n82714 & n83028;
  assign n83030 = n82717 & n83024;
  assign n83031 = ~n82714 & n83030;
  assign n83032 = ~n83025 & ~n83027;
  assign n83033 = ~n83029 & n83032;
  assign n83034 = ~n83031 & n83033;
  assign n83035 = n82713 & ~n83034;
  assign n83036 = ~n82713 & n83034;
  assign n83037 = ~n83035 & ~n83036;
  assign n83038 = n82704 & ~n83037;
  assign n83039 = n82700 & ~n82703;
  assign n83040 = ~n82573 & ~n82700;
  assign n83041 = ~n82702 & n83040;
  assign n83042 = ~n83039 & ~n83041;
  assign n83043 = n83037 & ~n83042;
  assign n83044 = ~n83038 & ~n83043;
  assign n83045 = n82700 & n82703;
  assign n83046 = ~n83037 & n83045;
  assign n83047 = n83044 & ~n83046;
  assign n83048 = n82699 & ~n83047;
  assign n83049 = ~n82699 & n83047;
  assign n83050 = ~n83048 & ~n83049;
  assign n83051 = n82698 & ~n83050;
  assign n83052 = ~n82699 & ~n83037;
  assign n83053 = n83045 & n83052;
  assign n83054 = ~n82699 & ~n83044;
  assign n83055 = n82699 & ~n83046;
  assign n83056 = n83044 & n83055;
  assign n83057 = ~n83053 & ~n83054;
  assign n83058 = ~n83056 & n83057;
  assign n83059 = ~n82698 & ~n83058;
  assign n83060 = ~n83051 & ~n83059;
  assign n83061 = P3_DATAO_REG_3_ & n80603;
  assign n83062 = ~n82228 & ~n82590;
  assign n83063 = ~n82227 & ~n83062;
  assign n83064 = ~n82597 & ~n83063;
  assign n83065 = ~n83060 & ~n83061;
  assign n83066 = ~n83064 & n83065;
  assign n83067 = n83060 & n83061;
  assign n83068 = ~n83065 & ~n83067;
  assign n83069 = n83064 & n83068;
  assign n83070 = ~n83066 & ~n83069;
  assign n83071 = n83061 & ~n83064;
  assign n83072 = n83060 & n83071;
  assign n83073 = n83070 & ~n83072;
  assign n83074 = n82694 & ~n83073;
  assign n83075 = ~n82694 & n83073;
  assign n83076 = ~n83074 & ~n83075;
  assign n83077 = n82693 & ~n83076;
  assign n83078 = ~n82694 & n83072;
  assign n83079 = n82694 & ~n83072;
  assign n83080 = n83070 & n83079;
  assign n83081 = ~n82694 & ~n83070;
  assign n83082 = ~n83078 & ~n83080;
  assign n83083 = ~n83081 & n83082;
  assign n83084 = ~n82693 & ~n83083;
  assign n83085 = ~n83077 & ~n83084;
  assign n83086 = n80600 & ~n83085;
  assign n83087 = ~n82688 & ~n83085;
  assign n83088 = ~n82689 & ~n83086;
  assign n83089 = ~n83087 & n83088;
  assign n83090 = ~n82694 & ~n83073;
  assign n83091 = ~n82693 & ~n83090;
  assign n83092 = ~n83080 & ~n83091;
  assign n83093 = ~SEL & DIN_30_;
  assign n83094 = P3_DATAO_REG_1_ & n83093;
  assign n83095 = P3_DATAO_REG_2_ & n80599;
  assign n83096 = n83094 & ~n83095;
  assign n83097 = ~n83094 & n83095;
  assign n83098 = ~n83096 & ~n83097;
  assign n83099 = ~n83060 & n83061;
  assign n83100 = ~n83060 & ~n83064;
  assign n83101 = ~n83071 & ~n83099;
  assign n83102 = ~n83100 & n83101;
  assign n83103 = n82700 & ~n83037;
  assign n83104 = ~n82703 & ~n83037;
  assign n83105 = ~n83039 & ~n83103;
  assign n83106 = ~n83104 & n83105;
  assign n83107 = P3_DATAO_REG_4_ & n80603;
  assign n83108 = ~n82712 & n83034;
  assign n83109 = ~n82711 & ~n83108;
  assign n83110 = n82714 & ~n83024;
  assign n83111 = ~n82717 & ~n83024;
  assign n83112 = ~n83026 & ~n83110;
  assign n83113 = ~n83111 & n83112;
  assign n83114 = ~n82725 & n83021;
  assign n83115 = ~n82724 & ~n83114;
  assign n83116 = ~n82736 & ~n83000;
  assign n83117 = ~n82735 & ~n83116;
  assign n83118 = ~n83007 & ~n83117;
  assign n83119 = P3_DATAO_REG_11_ & n77708;
  assign n83120 = ~n82988 & n82989;
  assign n83121 = ~n82988 & ~n82991;
  assign n83122 = ~n82998 & ~n83120;
  assign n83123 = ~n83121 & n83122;
  assign n83124 = ~n82740 & ~n82976;
  assign n83125 = ~n82739 & ~n83124;
  assign n83126 = ~n82983 & ~n83125;
  assign n83127 = ~n82963 & n82964;
  assign n83128 = ~n82963 & ~n82967;
  assign n83129 = ~n82974 & ~n83127;
  assign n83130 = ~n83128 & n83129;
  assign n83131 = ~n82745 & ~n82951;
  assign n83132 = ~n82744 & ~n83131;
  assign n83133 = ~n82958 & ~n83132;
  assign n83134 = ~n82938 & n82939;
  assign n83135 = ~n82938 & ~n82942;
  assign n83136 = ~n82949 & ~n83134;
  assign n83137 = ~n83135 & n83136;
  assign n83138 = ~n82750 & ~n82926;
  assign n83139 = ~n82749 & ~n83138;
  assign n83140 = ~n82933 & ~n83139;
  assign n83141 = P3_DATAO_REG_15_ & n78934;
  assign n83142 = P3_DATAO_REG_16_ & n77716;
  assign n83143 = n83141 & ~n83142;
  assign n83144 = ~n83141 & n83142;
  assign n83145 = ~n83143 & ~n83144;
  assign n83146 = ~n82913 & n82914;
  assign n83147 = ~n82913 & ~n82917;
  assign n83148 = ~n82924 & ~n83146;
  assign n83149 = ~n83147 & n83148;
  assign n83150 = ~n82889 & n82890;
  assign n83151 = ~n82889 & ~n82892;
  assign n83152 = ~n82899 & ~n83150;
  assign n83153 = ~n83151 & n83152;
  assign n83154 = ~n82760 & ~n82877;
  assign n83155 = ~n82759 & ~n83154;
  assign n83156 = ~n82885 & ~n83155;
  assign n83157 = ~n82764 & ~n82853;
  assign n83158 = ~n82763 & ~n83157;
  assign n83159 = ~n82860 & ~n83158;
  assign n83160 = ~n82840 & n82841;
  assign n83161 = ~n82840 & ~n82844;
  assign n83162 = ~n82851 & ~n83160;
  assign n83163 = ~n83161 & n83162;
  assign n83164 = P3_DATAO_REG_22_ & n78036;
  assign n83165 = P3_DATAO_REG_23_ & n77955;
  assign n83166 = n83164 & ~n83165;
  assign n83167 = ~n83164 & n83165;
  assign n83168 = ~n83166 & ~n83167;
  assign n83169 = P3_DATAO_REG_25_ & n77434;
  assign n83170 = P3_DATAO_REG_24_ & n77688;
  assign n83171 = n83169 & ~n83170;
  assign n83172 = ~n83169 & n83170;
  assign n83173 = ~n83171 & ~n83172;
  assign n83174 = P3_DATAO_REG_29_ & n77451;
  assign n83175 = n77440 & n83174;
  assign n83176 = P3_DATAO_REG_29_ & n77440;
  assign n83177 = P3_DATAO_REG_30_ & n77442;
  assign n83178 = ~n77444 & ~n83177;
  assign n83179 = P3_DATAO_REG_31_ & n83178;
  assign n83180 = ~P3_DATAO_REG_31_ & n83177;
  assign n83181 = P3_DATAO_REG_30_ & n77451;
  assign n83182 = ~n83179 & ~n83180;
  assign n83183 = ~n83181 & n83182;
  assign n83184 = n83176 & ~n83183;
  assign n83185 = ~n83176 & n83183;
  assign n83186 = ~n83184 & ~n83185;
  assign n83187 = ~n83174 & n83186;
  assign n83188 = ~n83175 & ~n83187;
  assign n83189 = ~n82782 & n82784;
  assign n83190 = ~n82781 & ~n83189;
  assign n83191 = P3_DATAO_REG_28_ & n77438;
  assign n83192 = n83190 & ~n83191;
  assign n83193 = ~n83190 & n83191;
  assign n83194 = ~n83192 & ~n83193;
  assign n83195 = ~n83188 & n83194;
  assign n83196 = n83188 & ~n83194;
  assign n83197 = ~n83195 & ~n83196;
  assign n83198 = ~n82791 & n82792;
  assign n83199 = ~n82791 & ~n82794;
  assign n83200 = ~n82801 & ~n83198;
  assign n83201 = ~n83199 & n83200;
  assign n83202 = P3_DATAO_REG_26_ & n77436;
  assign n83203 = P3_DATAO_REG_27_ & n77475;
  assign n83204 = n83202 & ~n83203;
  assign n83205 = ~n83202 & n83203;
  assign n83206 = ~n83204 & ~n83205;
  assign n83207 = n83201 & n83206;
  assign n83208 = ~n83201 & ~n83206;
  assign n83209 = ~n83207 & ~n83208;
  assign n83210 = ~n83197 & n83209;
  assign n83211 = n83197 & ~n83209;
  assign n83212 = ~n83210 & ~n83211;
  assign n83213 = ~n82774 & ~n82803;
  assign n83214 = ~n82773 & ~n83213;
  assign n83215 = ~n82811 & ~n83214;
  assign n83216 = ~n83212 & ~n83215;
  assign n83217 = n83212 & n83215;
  assign n83218 = ~n83216 & ~n83217;
  assign n83219 = ~n83173 & n83218;
  assign n83220 = n83173 & ~n83218;
  assign n83221 = ~n83219 & ~n83220;
  assign n83222 = ~n82815 & n82816;
  assign n83223 = ~n82815 & ~n82819;
  assign n83224 = ~n82826 & ~n83222;
  assign n83225 = ~n83223 & n83224;
  assign n83226 = ~n83221 & ~n83225;
  assign n83227 = n83221 & n83225;
  assign n83228 = ~n83226 & ~n83227;
  assign n83229 = ~n82769 & ~n82828;
  assign n83230 = ~n82768 & ~n83229;
  assign n83231 = ~n82835 & ~n83230;
  assign n83232 = ~n83228 & ~n83231;
  assign n83233 = n83228 & n83231;
  assign n83234 = ~n83232 & ~n83233;
  assign n83235 = ~n83168 & n83234;
  assign n83236 = n83168 & ~n83234;
  assign n83237 = ~n83235 & ~n83236;
  assign n83238 = n83163 & n83237;
  assign n83239 = ~n83163 & ~n83237;
  assign n83240 = ~n83238 & ~n83239;
  assign n83241 = n83159 & n83240;
  assign n83242 = ~n83159 & ~n83240;
  assign n83243 = ~n83241 & ~n83242;
  assign n83244 = ~n82865 & n82866;
  assign n83245 = ~n82865 & ~n82868;
  assign n83246 = ~n82875 & ~n83244;
  assign n83247 = ~n83245 & n83246;
  assign n83248 = ~n83243 & ~n83247;
  assign n83249 = n83243 & n83247;
  assign n83250 = ~n83248 & ~n83249;
  assign n83251 = n83156 & n83250;
  assign n83252 = ~n83156 & ~n83250;
  assign n83253 = ~n83251 & ~n83252;
  assign n83254 = P3_DATAO_REG_19_ & n77722;
  assign n83255 = P3_DATAO_REG_21_ & n77726;
  assign n83256 = P3_DATAO_REG_20_ & n77724;
  assign n83257 = n83255 & ~n83256;
  assign n83258 = ~n83255 & n83256;
  assign n83259 = ~n83257 & ~n83258;
  assign n83260 = n83254 & n83259;
  assign n83261 = ~n83254 & ~n83259;
  assign n83262 = ~n83260 & ~n83261;
  assign n83263 = ~n83253 & n83262;
  assign n83264 = n83253 & ~n83262;
  assign n83265 = ~n83263 & ~n83264;
  assign n83266 = P3_DATAO_REG_18_ & n77720;
  assign n83267 = ~n83265 & ~n83266;
  assign n83268 = n83265 & n83266;
  assign n83269 = ~n83267 & ~n83268;
  assign n83270 = n83153 & n83269;
  assign n83271 = ~n83153 & ~n83269;
  assign n83272 = ~n83270 & ~n83271;
  assign n83273 = P3_DATAO_REG_17_ & n77718;
  assign n83274 = ~n83272 & ~n83273;
  assign n83275 = n83272 & n83273;
  assign n83276 = ~n83274 & ~n83275;
  assign n83277 = ~n82755 & ~n82901;
  assign n83278 = ~n82754 & ~n83277;
  assign n83279 = ~n82909 & ~n83278;
  assign n83280 = ~n83276 & ~n83279;
  assign n83281 = n83276 & n83279;
  assign n83282 = ~n83280 & ~n83281;
  assign n83283 = n83149 & n83282;
  assign n83284 = ~n83149 & ~n83282;
  assign n83285 = ~n83283 & ~n83284;
  assign n83286 = ~n83145 & n83285;
  assign n83287 = n83145 & ~n83285;
  assign n83288 = ~n83286 & ~n83287;
  assign n83289 = n83140 & n83288;
  assign n83290 = ~n83140 & ~n83288;
  assign n83291 = ~n83289 & ~n83290;
  assign n83292 = n83137 & n83291;
  assign n83293 = ~n83137 & ~n83291;
  assign n83294 = ~n83292 & ~n83293;
  assign n83295 = P3_DATAO_REG_14_ & n77714;
  assign n83296 = ~n83294 & ~n83295;
  assign n83297 = n83294 & n83295;
  assign n83298 = ~n83296 & ~n83297;
  assign n83299 = n83133 & n83298;
  assign n83300 = ~n83133 & ~n83298;
  assign n83301 = ~n83299 & ~n83300;
  assign n83302 = n83130 & n83301;
  assign n83303 = ~n83130 & ~n83301;
  assign n83304 = ~n83302 & ~n83303;
  assign n83305 = P3_DATAO_REG_13_ & n77712;
  assign n83306 = P3_DATAO_REG_12_ & n77710;
  assign n83307 = n83305 & ~n83306;
  assign n83308 = ~n83305 & n83306;
  assign n83309 = ~n83307 & ~n83308;
  assign n83310 = ~n83304 & n83309;
  assign n83311 = n83304 & ~n83309;
  assign n83312 = ~n83310 & ~n83311;
  assign n83313 = n83126 & n83312;
  assign n83314 = ~n83126 & ~n83312;
  assign n83315 = ~n83313 & ~n83314;
  assign n83316 = n83123 & n83315;
  assign n83317 = ~n83123 & ~n83315;
  assign n83318 = ~n83316 & ~n83317;
  assign n83319 = n83119 & n83318;
  assign n83320 = ~n83119 & ~n83318;
  assign n83321 = ~n83319 & ~n83320;
  assign n83322 = n83118 & n83321;
  assign n83323 = ~n83118 & ~n83321;
  assign n83324 = ~n83322 & ~n83323;
  assign n83325 = P3_DATAO_REG_10_ & n77706;
  assign n83326 = P3_DATAO_REG_9_ & n80109;
  assign n83327 = n83325 & ~n83326;
  assign n83328 = ~n83325 & n83326;
  assign n83329 = ~n83327 & ~n83328;
  assign n83330 = P3_DATAO_REG_8_ & n77704;
  assign n83331 = ~n83329 & ~n83330;
  assign n83332 = n83329 & n83330;
  assign n83333 = ~n83331 & ~n83332;
  assign n83334 = ~n83324 & n83333;
  assign n83335 = n83324 & ~n83333;
  assign n83336 = ~n83334 & ~n83335;
  assign n83337 = n82730 & ~n83012;
  assign n83338 = ~n82729 & ~n83012;
  assign n83339 = ~n83014 & ~n83337;
  assign n83340 = ~n83338 & n83339;
  assign n83341 = ~n83336 & ~n83340;
  assign n83342 = n83336 & n83340;
  assign n83343 = ~n83341 & ~n83342;
  assign n83344 = n83115 & n83343;
  assign n83345 = ~n83115 & ~n83343;
  assign n83346 = ~n83344 & ~n83345;
  assign n83347 = P3_DATAO_REG_7_ & n80609;
  assign n83348 = ~n83346 & ~n83347;
  assign n83349 = n83346 & n83347;
  assign n83350 = ~n83348 & ~n83349;
  assign n83351 = n83113 & n83350;
  assign n83352 = ~n83113 & ~n83350;
  assign n83353 = ~n83351 & ~n83352;
  assign n83354 = n83109 & n83353;
  assign n83355 = ~n83109 & ~n83353;
  assign n83356 = ~n83354 & ~n83355;
  assign n83357 = P3_DATAO_REG_6_ & n80607;
  assign n83358 = P3_DATAO_REG_5_ & n80605;
  assign n83359 = n83357 & ~n83358;
  assign n83360 = ~n83357 & n83358;
  assign n83361 = ~n83359 & ~n83360;
  assign n83362 = ~n83356 & n83361;
  assign n83363 = n83356 & ~n83361;
  assign n83364 = ~n83362 & ~n83363;
  assign n83365 = n83107 & n83364;
  assign n83366 = ~n83107 & ~n83364;
  assign n83367 = ~n83365 & ~n83366;
  assign n83368 = n83106 & n83367;
  assign n83369 = ~n83106 & ~n83367;
  assign n83370 = ~n83368 & ~n83369;
  assign n83371 = P3_DATAO_REG_3_ & n80601;
  assign n83372 = ~n83370 & ~n83371;
  assign n83373 = n83370 & n83371;
  assign n83374 = ~n83372 & ~n83373;
  assign n83375 = ~n82699 & ~n83047;
  assign n83376 = ~n82698 & ~n83375;
  assign n83377 = ~n83056 & ~n83376;
  assign n83378 = ~n83374 & ~n83377;
  assign n83379 = n83374 & n83377;
  assign n83380 = ~n83378 & ~n83379;
  assign n83381 = n83102 & n83380;
  assign n83382 = ~n83102 & ~n83380;
  assign n83383 = ~n83381 & ~n83382;
  assign n83384 = ~n83098 & n83383;
  assign n83385 = n83098 & ~n83383;
  assign n83386 = ~n83384 & ~n83385;
  assign n83387 = n83092 & n83386;
  assign n83388 = ~n83092 & ~n83386;
  assign n83389 = ~n83387 & ~n83388;
  assign n83390 = n83089 & n83389;
  assign n83391 = ~n83089 & ~n83389;
  assign n83392 = ~n83390 & ~n83391;
  assign n83393 = ~SEL & DIN_31_;
  assign n83394 = ~P3_DATAO_REG_0_ & n83393;
  assign n83395 = P3_DATAO_REG_0_ & n83093;
  assign n83396 = n80602 & ~n82612;
  assign n83397 = ~n80602 & n82612;
  assign n83398 = ~n83396 & ~n83397;
  assign n83399 = n82686 & ~n83398;
  assign n83400 = ~n80602 & n82603;
  assign n83401 = ~n80602 & ~n82610;
  assign n83402 = ~n82611 & ~n83400;
  assign n83403 = ~n83401 & n83402;
  assign n83404 = ~n82686 & ~n83403;
  assign n83405 = ~n83399 & ~n83404;
  assign n83406 = P3_DATAO_REG_0_ & n80599;
  assign n83407 = n83405 & ~n83406;
  assign n83408 = ~n82614 & ~n82664;
  assign n83409 = ~n82683 & n83408;
  assign n83410 = ~n82685 & ~n83409;
  assign n83411 = n82678 & ~n83410;
  assign n83412 = ~n82614 & n82684;
  assign n83413 = ~n82685 & ~n83412;
  assign n83414 = ~n82678 & n83413;
  assign n83415 = ~n83411 & ~n83414;
  assign n83416 = P3_DATAO_REG_0_ & n80603;
  assign n83417 = P3_DATAO_REG_0_ & n80605;
  assign n83418 = P3_DATAO_REG_0_ & n80607;
  assign n83419 = ~n82633 & ~n82639;
  assign n83420 = n82638 & ~n83419;
  assign n83421 = ~n82638 & n83419;
  assign n83422 = ~n83420 & ~n83421;
  assign n83423 = n83418 & ~n83422;
  assign n83424 = ~n83418 & n83422;
  assign n83425 = P3_DATAO_REG_0_ & n80609;
  assign n83426 = n77705 & ~n80585;
  assign n83427 = ~n80410 & ~n80585;
  assign n83428 = ~n80411 & ~n83426;
  assign n83429 = ~n83427 & n83428;
  assign n83430 = n83425 & ~n83429;
  assign n83431 = ~n82620 & ~n82623;
  assign n83432 = n82620 & n82623;
  assign n83433 = ~n83431 & ~n83432;
  assign n83434 = n82630 & n83433;
  assign n83435 = ~n82630 & n83431;
  assign n83436 = n82620 & n82631;
  assign n83437 = ~n83434 & ~n83435;
  assign n83438 = ~n83436 & n83437;
  assign n83439 = ~n83429 & n83438;
  assign n83440 = n83425 & n83438;
  assign n83441 = ~n83430 & ~n83439;
  assign n83442 = ~n83440 & n83441;
  assign n83443 = ~n83424 & ~n83442;
  assign n83444 = ~n83423 & ~n83443;
  assign n83445 = n83417 & ~n83444;
  assign n83446 = ~n82615 & n82646;
  assign n83447 = ~n82647 & ~n83446;
  assign n83448 = n82641 & ~n83447;
  assign n83449 = ~n82615 & ~n82646;
  assign n83450 = ~n82641 & n83449;
  assign n83451 = n82642 & n82646;
  assign n83452 = ~n83448 & ~n83450;
  assign n83453 = ~n83451 & n83452;
  assign n83454 = ~n83417 & ~n83423;
  assign n83455 = ~n83443 & n83454;
  assign n83456 = n83453 & ~n83455;
  assign n83457 = ~n83445 & ~n83456;
  assign n83458 = n83416 & ~n83457;
  assign n83459 = n82662 & ~n82663;
  assign n83460 = n82650 & n83459;
  assign n83461 = ~n82650 & n82664;
  assign n83462 = ~n83460 & ~n83461;
  assign n83463 = n82650 & ~n82663;
  assign n83464 = ~n82650 & n82663;
  assign n83465 = ~n83463 & ~n83464;
  assign n83466 = ~n82662 & n83465;
  assign n83467 = n83462 & ~n83466;
  assign n83468 = n83416 & ~n83467;
  assign n83469 = ~n83457 & ~n83467;
  assign n83470 = ~n83458 & ~n83468;
  assign n83471 = ~n83469 & n83470;
  assign n83472 = n83415 & ~n83471;
  assign n83473 = P3_DATAO_REG_0_ & n80601;
  assign n83474 = n83415 & n83473;
  assign n83475 = ~n83471 & n83473;
  assign n83476 = ~n83472 & ~n83474;
  assign n83477 = ~n83475 & n83476;
  assign n83478 = ~n83407 & ~n83477;
  assign n83479 = ~n83405 & n83406;
  assign n83480 = ~n83478 & ~n83479;
  assign n83481 = n83395 & ~n83480;
  assign n83482 = ~n83395 & ~n83406;
  assign n83483 = n83405 & n83482;
  assign n83484 = n82689 & n83085;
  assign n83485 = ~n83472 & ~n83475;
  assign n83486 = ~n83395 & n83485;
  assign n83487 = ~n83474 & n83486;
  assign n83488 = ~n83479 & n83487;
  assign n83489 = ~n83483 & ~n83484;
  assign n83490 = ~n83488 & n83489;
  assign n83491 = ~n80600 & ~n83085;
  assign n83492 = ~n82688 & n83491;
  assign n83493 = n80600 & n83085;
  assign n83494 = ~n83491 & ~n83493;
  assign n83495 = n82688 & n83494;
  assign n83496 = ~n83492 & ~n83495;
  assign n83497 = n83490 & n83496;
  assign n83498 = ~n83394 & ~n83481;
  assign n83499 = ~n83497 & n83498;
  assign n83500 = ~n83392 & ~n83499;
  assign n83501 = n83392 & n83499;
  assign n83502 = P3_DATAO_REG_31_ & ~n83393;
  assign n83503 = ~P3_DATAO_REG_31_ & n83393;
  assign n83504 = ~n83502 & ~n83503;
  assign n83505 = ~n83500 & ~n83501;
  assign n83506 = n83504 & n83505;
  assign n83507 = ~n83395 & ~n83479;
  assign n83508 = ~n83478 & n83507;
  assign n83509 = ~n83484 & n83496;
  assign n83510 = ~n83508 & n83509;
  assign n83511 = n83498 & ~n83510;
  assign n83512 = ~n83392 & ~n83511;
  assign n83513 = n83392 & n83511;
  assign n83514 = ~n83512 & ~n83513;
  assign n83515 = ~n83504 & ~n83514;
  assign n83516 = ~n83506 & ~n83515;
  assign n83517 = ~n12802 & ~n83516;
  assign n83518 = ~n80598 & ~n83517;
  assign n83519 = n80592 & ~n83518;
  assign n83520 = n80597 & ~n83519;
  assign n83521 = ~n77418 & n80597;
  assign n14841 = ~n83520 & ~n83521;
  assign n83523 = P2_P1_INSTQUEUE_REG_15__6_ & ~n77424;
  assign n83524 = P2_BUF1_REG_6_ & n12802;
  assign n83525 = n77435 & ~n77612;
  assign n83526 = ~n77435 & n77612;
  assign n83527 = ~n83525 & ~n83526;
  assign n83528 = n77553 & ~n83527;
  assign n83529 = ~n77435 & ~n77612;
  assign n83530 = ~n77553 & n83529;
  assign n83531 = n77554 & n77612;
  assign n83532 = ~n83528 & ~n83530;
  assign n83533 = ~n83531 & n83532;
  assign n83534 = ~n12802 & ~n83533;
  assign n83535 = ~n83524 & ~n83534;
  assign n83536 = n77374 & ~n83535;
  assign n83537 = n77432 & n83536;
  assign n83538 = ~n76765 & n77426;
  assign n83539 = n77369 & n83538;
  assign n83540 = P2_BUF1_REG_22_ & n12802;
  assign n83541 = n80413 & ~n80582;
  assign n83542 = ~n80413 & n80582;
  assign n83543 = ~n83541 & ~n83542;
  assign n83544 = n80573 & ~n83543;
  assign n83545 = ~n80413 & ~n80582;
  assign n83546 = ~n80573 & n83545;
  assign n83547 = n80574 & n80582;
  assign n83548 = ~n83544 & ~n83546;
  assign n83549 = ~n83547 & n83548;
  assign n83550 = ~n12802 & ~n83549;
  assign n83551 = ~n83540 & ~n83550;
  assign n83552 = n80592 & ~n83551;
  assign n83553 = n77420 & n83552;
  assign n83554 = P2_BUF1_REG_30_ & n12802;
  assign n83555 = n83395 & ~n83509;
  assign n83556 = ~n83395 & n83509;
  assign n83557 = ~n83555 & ~n83556;
  assign n83558 = n83480 & ~n83557;
  assign n83559 = ~n83395 & ~n83509;
  assign n83560 = ~n83480 & n83559;
  assign n83561 = n83481 & n83509;
  assign n83562 = ~n83558 & ~n83560;
  assign n83563 = ~n83561 & n83562;
  assign n83564 = ~n12802 & ~n83563;
  assign n83565 = ~n83554 & ~n83564;
  assign n83566 = n80592 & ~n83565;
  assign n83567 = n77418 & n83566;
  assign n83568 = ~n83523 & ~n83537;
  assign n83569 = ~n83539 & n83568;
  assign n83570 = ~n83553 & n83569;
  assign n14846 = n83567 | ~n83570;
  assign n83572 = P2_P1_INSTQUEUE_REG_15__5_ & ~n77424;
  assign n83573 = P2_BUF1_REG_5_ & n12802;
  assign n83574 = ~n77437 & ~n77515;
  assign n83575 = n77437 & n77515;
  assign n83576 = ~n83574 & ~n83575;
  assign n83577 = n77551 & ~n83576;
  assign n83578 = ~n77516 & ~n77517;
  assign n83579 = ~n77551 & ~n83578;
  assign n83580 = ~n83577 & ~n83579;
  assign n83581 = ~n12802 & ~n83580;
  assign n83582 = ~n83573 & ~n83581;
  assign n83583 = n77374 & ~n83582;
  assign n83584 = n77432 & n83583;
  assign n83585 = ~n76734 & n77426;
  assign n83586 = n77369 & n83585;
  assign n83587 = P2_BUF1_REG_21_ & n12802;
  assign n83588 = ~n80414 & ~n80418;
  assign n83589 = n80414 & n80418;
  assign n83590 = ~n83588 & ~n83589;
  assign n83591 = n80571 & ~n83590;
  assign n83592 = ~n80571 & n83590;
  assign n83593 = ~n83591 & ~n83592;
  assign n83594 = ~n12802 & ~n83593;
  assign n83595 = ~n83587 & ~n83594;
  assign n83596 = n80592 & ~n83595;
  assign n83597 = n77420 & n83596;
  assign n83598 = P2_BUF1_REG_29_ & n12802;
  assign n83599 = ~n83405 & ~n83406;
  assign n83600 = n83405 & n83406;
  assign n83601 = ~n83599 & ~n83600;
  assign n83602 = n83477 & ~n83601;
  assign n83603 = ~n83407 & ~n83479;
  assign n83604 = ~n83477 & ~n83603;
  assign n83605 = ~n83602 & ~n83604;
  assign n83606 = ~n12802 & ~n83605;
  assign n83607 = ~n83598 & ~n83606;
  assign n83608 = n80592 & ~n83607;
  assign n83609 = n77418 & n83608;
  assign n83610 = ~n83572 & ~n83584;
  assign n83611 = ~n83586 & n83610;
  assign n83612 = ~n83597 & n83611;
  assign n14851 = n83609 | ~n83612;
  assign n83614 = P2_P1_INSTQUEUE_REG_15__4_ & ~n77424;
  assign n83615 = P2_BUF1_REG_4_ & n12802;
  assign n83616 = n77518 & ~n77548;
  assign n83617 = ~n77518 & n77548;
  assign n83618 = ~n83616 & ~n83617;
  assign n83619 = n77539 & ~n83618;
  assign n83620 = ~n77518 & ~n77548;
  assign n83621 = ~n77539 & n83620;
  assign n83622 = n77540 & n77548;
  assign n83623 = ~n83619 & ~n83621;
  assign n83624 = ~n83622 & n83623;
  assign n83625 = ~n12802 & ~n83624;
  assign n83626 = ~n83615 & ~n83625;
  assign n83627 = n77374 & ~n83626;
  assign n83628 = n77432 & n83627;
  assign n83629 = ~n76797 & n77426;
  assign n83630 = n77369 & n83629;
  assign n83631 = P2_BUF1_REG_20_ & n12802;
  assign n83632 = ~n80421 & ~n80568;
  assign n83633 = n80421 & n80568;
  assign n83634 = ~n83632 & ~n83633;
  assign n83635 = n80561 & n83634;
  assign n83636 = ~n80561 & n83632;
  assign n83637 = n80562 & n80568;
  assign n83638 = ~n83635 & ~n83636;
  assign n83639 = ~n83637 & n83638;
  assign n83640 = ~n12802 & ~n83639;
  assign n83641 = ~n83631 & ~n83640;
  assign n83642 = n80592 & ~n83641;
  assign n83643 = n77420 & n83642;
  assign n83644 = P2_BUF1_REG_28_ & n12802;
  assign n83645 = n83471 & ~n83473;
  assign n83646 = ~n83475 & ~n83645;
  assign n83647 = ~n83415 & n83646;
  assign n83648 = n83415 & n83645;
  assign n83649 = ~n83471 & n83474;
  assign n83650 = ~n83647 & ~n83648;
  assign n83651 = ~n83649 & n83650;
  assign n83652 = ~n12802 & ~n83651;
  assign n83653 = ~n83644 & ~n83652;
  assign n83654 = n80592 & ~n83653;
  assign n83655 = n77418 & n83654;
  assign n83656 = ~n83614 & ~n83628;
  assign n83657 = ~n83630 & n83656;
  assign n83658 = ~n83643 & n83657;
  assign n14856 = n83655 | ~n83658;
  assign n83660 = P2_P1_INSTQUEUE_REG_15__3_ & ~n77424;
  assign n83661 = P2_BUF1_REG_3_ & n12802;
  assign n83662 = ~n77519 & ~n77523;
  assign n83663 = n77519 & n77523;
  assign n83664 = ~n83662 & ~n83663;
  assign n83665 = n77537 & ~n83664;
  assign n83666 = ~n77524 & ~n77525;
  assign n83667 = ~n77537 & ~n83666;
  assign n83668 = ~n83665 & ~n83667;
  assign n83669 = ~n12802 & ~n83668;
  assign n83670 = ~n83661 & ~n83669;
  assign n83671 = n77374 & ~n83670;
  assign n83672 = n77432 & n83671;
  assign n83673 = ~n76859 & n77426;
  assign n83674 = n77369 & n83673;
  assign n83675 = P2_BUF1_REG_19_ & n12802;
  assign n83676 = ~n80422 & ~n80426;
  assign n83677 = n80422 & n80426;
  assign n83678 = ~n83676 & ~n83677;
  assign n83679 = n80559 & ~n83678;
  assign n83680 = ~n80427 & ~n80428;
  assign n83681 = ~n80559 & ~n83680;
  assign n83682 = ~n83679 & ~n83681;
  assign n83683 = ~n12802 & ~n83682;
  assign n83684 = ~n83675 & ~n83683;
  assign n83685 = n80592 & ~n83684;
  assign n83686 = n77420 & n83685;
  assign n83687 = P2_BUF1_REG_27_ & n12802;
  assign n83688 = ~n83416 & n83467;
  assign n83689 = ~n83468 & ~n83688;
  assign n83690 = n83457 & n83689;
  assign n83691 = ~n83457 & ~n83689;
  assign n83692 = ~n83690 & ~n83691;
  assign n83693 = ~n12802 & ~n83692;
  assign n83694 = ~n83687 & ~n83693;
  assign n83695 = n80592 & ~n83694;
  assign n83696 = n77418 & n83695;
  assign n83697 = ~n83660 & ~n83672;
  assign n83698 = ~n83674 & n83697;
  assign n83699 = ~n83686 & n83698;
  assign n14861 = n83696 | ~n83699;
  assign n83701 = P2_P1_INSTQUEUE_REG_15__2_ & ~n77424;
  assign n83702 = P2_BUF1_REG_2_ & n12802;
  assign n83703 = n77529 & ~n77535;
  assign n83704 = ~n77529 & n77535;
  assign n83705 = ~n83703 & ~n83704;
  assign n83706 = ~n77528 & n83705;
  assign n83707 = n77528 & n83704;
  assign n83708 = n77530 & ~n77535;
  assign n83709 = ~n83706 & ~n83707;
  assign n83710 = ~n83708 & n83709;
  assign n83711 = ~n12802 & ~n83710;
  assign n83712 = ~n83702 & ~n83711;
  assign n83713 = n77374 & ~n83712;
  assign n83714 = n77432 & n83713;
  assign n83715 = ~n76890 & n77426;
  assign n83716 = n77369 & n83715;
  assign n83717 = P2_BUF1_REG_18_ & n12802;
  assign n83718 = n80429 & ~n80556;
  assign n83719 = ~n80429 & n80556;
  assign n83720 = ~n83718 & ~n83719;
  assign n83721 = n80547 & ~n83720;
  assign n83722 = ~n80429 & ~n80556;
  assign n83723 = ~n80547 & n83722;
  assign n83724 = n80548 & n80556;
  assign n83725 = ~n83721 & ~n83723;
  assign n83726 = ~n83724 & n83725;
  assign n83727 = ~n12802 & ~n83726;
  assign n83728 = ~n83717 & ~n83727;
  assign n83729 = n80592 & ~n83728;
  assign n83730 = n77420 & n83729;
  assign n83731 = P2_BUF1_REG_26_ & n12802;
  assign n83732 = n83417 & ~n83453;
  assign n83733 = ~n83417 & n83453;
  assign n83734 = ~n83732 & ~n83733;
  assign n83735 = n83444 & ~n83734;
  assign n83736 = ~n83417 & ~n83453;
  assign n83737 = ~n83444 & n83736;
  assign n83738 = n83445 & n83453;
  assign n83739 = ~n83735 & ~n83737;
  assign n83740 = ~n83738 & n83739;
  assign n83741 = ~n12802 & ~n83740;
  assign n83742 = ~n83731 & ~n83741;
  assign n83743 = n80592 & ~n83742;
  assign n83744 = n77418 & n83743;
  assign n83745 = ~n83701 & ~n83714;
  assign n83746 = ~n83716 & n83745;
  assign n83747 = ~n83730 & n83746;
  assign n14866 = n83744 | ~n83747;
  assign n83749 = P2_P1_INSTQUEUE_REG_15__1_ & ~n77424;
  assign n83750 = P2_BUF1_REG_1_ & n12802;
  assign n83751 = P3_DATAO_REG_1_ & n77444;
  assign n83752 = P3_DATAO_REG_0_ & n77442;
  assign n83753 = n83751 & ~n83752;
  assign n83754 = ~n83751 & n83752;
  assign n83755 = ~n83753 & ~n83754;
  assign n83756 = ~n12802 & ~n83755;
  assign n83757 = ~n83750 & ~n83756;
  assign n83758 = n77374 & ~n83757;
  assign n83759 = n77432 & n83758;
  assign n83760 = ~n76925 & n77426;
  assign n83761 = n77369 & n83760;
  assign n83762 = P2_BUF1_REG_17_ & n12802;
  assign n83763 = ~n80537 & ~n80545;
  assign n83764 = n80544 & n83763;
  assign n83765 = ~n80544 & ~n83763;
  assign n83766 = ~n83764 & ~n83765;
  assign n83767 = ~n12802 & ~n83766;
  assign n83768 = ~n83762 & ~n83767;
  assign n83769 = n80592 & ~n83768;
  assign n83770 = n77420 & n83769;
  assign n83771 = P2_BUF1_REG_25_ & n12802;
  assign n83772 = ~n83418 & ~n83422;
  assign n83773 = n83418 & n83422;
  assign n83774 = ~n83772 & ~n83773;
  assign n83775 = n83442 & ~n83774;
  assign n83776 = ~n83423 & ~n83424;
  assign n83777 = ~n83442 & ~n83776;
  assign n83778 = ~n83775 & ~n83777;
  assign n83779 = ~n12802 & ~n83778;
  assign n83780 = ~n83771 & ~n83779;
  assign n83781 = n80592 & ~n83780;
  assign n83782 = n77418 & n83781;
  assign n83783 = ~n83749 & ~n83759;
  assign n83784 = ~n83761 & n83783;
  assign n83785 = ~n83770 & n83784;
  assign n14871 = n83782 | ~n83785;
  assign n83787 = P2_P1_INSTQUEUE_REG_15__0_ & ~n77424;
  assign n83788 = P2_BUF1_REG_0_ & n12802;
  assign n83789 = ~n12802 & n77527;
  assign n83790 = ~n83788 & ~n83789;
  assign n83791 = n77374 & ~n83790;
  assign n83792 = n77432 & n83791;
  assign n83793 = ~n76956 & n77426;
  assign n83794 = n77369 & n83793;
  assign n83795 = P2_BUF1_REG_16_ & n12802;
  assign n83796 = n80439 & ~n80534;
  assign n83797 = ~n80439 & n80534;
  assign n83798 = ~n83796 & ~n83797;
  assign n83799 = ~n80438 & n83798;
  assign n83800 = n80438 & n83797;
  assign n83801 = n80440 & ~n80534;
  assign n83802 = ~n83799 & ~n83800;
  assign n83803 = ~n83801 & n83802;
  assign n83804 = ~n12802 & ~n83803;
  assign n83805 = ~n83795 & ~n83804;
  assign n83806 = n80592 & ~n83805;
  assign n83807 = n77420 & n83806;
  assign n83808 = P2_BUF1_REG_24_ & n12802;
  assign n83809 = n83425 & ~n83438;
  assign n83810 = ~n83425 & n83438;
  assign n83811 = ~n83809 & ~n83810;
  assign n83812 = n83429 & ~n83811;
  assign n83813 = ~n83425 & ~n83438;
  assign n83814 = ~n83429 & n83813;
  assign n83815 = n83430 & n83438;
  assign n83816 = ~n83812 & ~n83814;
  assign n83817 = ~n83815 & n83816;
  assign n83818 = ~n12802 & ~n83817;
  assign n83819 = ~n83808 & ~n83818;
  assign n83820 = n80592 & ~n83819;
  assign n83821 = n77418 & n83820;
  assign n83822 = ~n83787 & ~n83792;
  assign n83823 = ~n83794 & n83822;
  assign n83824 = ~n83807 & n83823;
  assign n14876 = n83821 | ~n83824;
  assign n83826 = P2_P1_INSTQUEUEWR_ADDR_REG_3_ & P2_P1_INSTQUEUEWR_ADDR_REG_1_;
  assign n83827 = P2_P1_INSTQUEUEWR_ADDR_REG_2_ & ~P2_P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n83828 = n83826 & n83827;
  assign n83829 = P2_P1_STATE2_REG_3_ & ~n83828;
  assign n83830 = n77374 & ~n83829;
  assign n83831 = n77382 & n77392;
  assign n83832 = ~n83828 & ~n83831;
  assign n83833 = P2_P1_INSTQUEUEWR_ADDR_REG_0_ & ~n77397;
  assign n83834 = n77417 & n83833;
  assign n83835 = n77395 & n77419;
  assign n83836 = ~n83834 & ~n83835;
  assign n83837 = n77391 & ~n83836;
  assign n83838 = n83832 & ~n83837;
  assign n83839 = n83830 & ~n83838;
  assign n83840 = P2_P1_INSTQUEUE_REG_14__7_ & ~n83839;
  assign n83841 = n77427 & n83828;
  assign n83842 = n77429 & n83836;
  assign n83843 = n77391 & ~n83842;
  assign n83844 = ~n83832 & ~n83843;
  assign n83845 = n77701 & n83844;
  assign n83846 = n80593 & n83835;
  assign n83847 = ~n83840 & ~n83841;
  assign n83848 = ~n83845 & n83847;
  assign n83849 = ~n83846 & n83848;
  assign n83850 = ~n83519 & n83849;
  assign n83851 = ~n83834 & n83849;
  assign n14881 = ~n83850 & ~n83851;
  assign n83853 = P2_P1_INSTQUEUE_REG_14__6_ & ~n83839;
  assign n83854 = n83536 & n83844;
  assign n83855 = n83538 & n83828;
  assign n83856 = n83552 & n83835;
  assign n83857 = n83566 & n83834;
  assign n83858 = ~n83853 & ~n83854;
  assign n83859 = ~n83855 & n83858;
  assign n83860 = ~n83856 & n83859;
  assign n14886 = n83857 | ~n83860;
  assign n83862 = P2_P1_INSTQUEUE_REG_14__5_ & ~n83839;
  assign n83863 = n83583 & n83844;
  assign n83864 = n83585 & n83828;
  assign n83865 = n83596 & n83835;
  assign n83866 = n83608 & n83834;
  assign n83867 = ~n83862 & ~n83863;
  assign n83868 = ~n83864 & n83867;
  assign n83869 = ~n83865 & n83868;
  assign n14891 = n83866 | ~n83869;
  assign n83871 = P2_P1_INSTQUEUE_REG_14__4_ & ~n83839;
  assign n83872 = n83627 & n83844;
  assign n83873 = n83629 & n83828;
  assign n83874 = n83642 & n83835;
  assign n83875 = n83654 & n83834;
  assign n83876 = ~n83871 & ~n83872;
  assign n83877 = ~n83873 & n83876;
  assign n83878 = ~n83874 & n83877;
  assign n14896 = n83875 | ~n83878;
  assign n83880 = P2_P1_INSTQUEUE_REG_14__3_ & ~n83839;
  assign n83881 = n83671 & n83844;
  assign n83882 = n83673 & n83828;
  assign n83883 = n83685 & n83835;
  assign n83884 = n83695 & n83834;
  assign n83885 = ~n83880 & ~n83881;
  assign n83886 = ~n83882 & n83885;
  assign n83887 = ~n83883 & n83886;
  assign n14901 = n83884 | ~n83887;
  assign n83889 = P2_P1_INSTQUEUE_REG_14__2_ & ~n83839;
  assign n83890 = n83713 & n83844;
  assign n83891 = n83715 & n83828;
  assign n83892 = n83729 & n83835;
  assign n83893 = n83743 & n83834;
  assign n83894 = ~n83889 & ~n83890;
  assign n83895 = ~n83891 & n83894;
  assign n83896 = ~n83892 & n83895;
  assign n14906 = n83893 | ~n83896;
  assign n83898 = P2_P1_INSTQUEUE_REG_14__1_ & ~n83839;
  assign n83899 = n83758 & n83844;
  assign n83900 = n83760 & n83828;
  assign n83901 = n83769 & n83835;
  assign n83902 = n83781 & n83834;
  assign n83903 = ~n83898 & ~n83899;
  assign n83904 = ~n83900 & n83903;
  assign n83905 = ~n83901 & n83904;
  assign n14911 = n83902 | ~n83905;
  assign n83907 = P2_P1_INSTQUEUE_REG_14__0_ & ~n83839;
  assign n83908 = n83791 & n83844;
  assign n83909 = n83793 & n83828;
  assign n83910 = n83806 & n83835;
  assign n83911 = n83820 & n83834;
  assign n83912 = ~n83907 & ~n83908;
  assign n83913 = ~n83909 & n83912;
  assign n83914 = ~n83910 & n83913;
  assign n14916 = n83911 | ~n83914;
  assign n83916 = P2_P1_INSTQUEUEWR_ADDR_REG_3_ & P2_P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n83917 = n77383 & n83916;
  assign n83918 = P2_P1_STATE2_REG_3_ & ~n83917;
  assign n83919 = n77374 & ~n83918;
  assign n83920 = n77382 & n77393;
  assign n83921 = ~n83917 & ~n83920;
  assign n83922 = ~P2_P1_INSTQUEUEWR_ADDR_REG_0_ & n77397;
  assign n83923 = n77417 & n83922;
  assign n83924 = n77396 & n77419;
  assign n83925 = ~n83923 & ~n83924;
  assign n83926 = n77391 & ~n83925;
  assign n83927 = n83921 & ~n83926;
  assign n83928 = n83919 & ~n83927;
  assign n83929 = P2_P1_INSTQUEUE_REG_13__7_ & ~n83928;
  assign n83930 = n77427 & n83917;
  assign n83931 = n77429 & n83925;
  assign n83932 = n77391 & ~n83931;
  assign n83933 = ~n83921 & ~n83932;
  assign n83934 = n77701 & n83933;
  assign n83935 = n80593 & n83924;
  assign n83936 = ~n83929 & ~n83930;
  assign n83937 = ~n83934 & n83936;
  assign n83938 = ~n83935 & n83937;
  assign n83939 = ~n83519 & n83938;
  assign n83940 = ~n83923 & n83938;
  assign n14921 = ~n83939 & ~n83940;
  assign n83942 = P2_P1_INSTQUEUE_REG_13__6_ & ~n83928;
  assign n83943 = n83536 & n83933;
  assign n83944 = n83538 & n83917;
  assign n83945 = n83552 & n83924;
  assign n83946 = n83566 & n83923;
  assign n83947 = ~n83942 & ~n83943;
  assign n83948 = ~n83944 & n83947;
  assign n83949 = ~n83945 & n83948;
  assign n14926 = n83946 | ~n83949;
  assign n83951 = P2_P1_INSTQUEUE_REG_13__5_ & ~n83928;
  assign n83952 = n83583 & n83933;
  assign n83953 = n83585 & n83917;
  assign n83954 = n83596 & n83924;
  assign n83955 = n83608 & n83923;
  assign n83956 = ~n83951 & ~n83952;
  assign n83957 = ~n83953 & n83956;
  assign n83958 = ~n83954 & n83957;
  assign n14931 = n83955 | ~n83958;
  assign n83960 = P2_P1_INSTQUEUE_REG_13__4_ & ~n83928;
  assign n83961 = n83627 & n83933;
  assign n83962 = n83629 & n83917;
  assign n83963 = n83642 & n83924;
  assign n83964 = n83654 & n83923;
  assign n83965 = ~n83960 & ~n83961;
  assign n83966 = ~n83962 & n83965;
  assign n83967 = ~n83963 & n83966;
  assign n14936 = n83964 | ~n83967;
  assign n83969 = P2_P1_INSTQUEUE_REG_13__3_ & ~n83928;
  assign n83970 = n83671 & n83933;
  assign n83971 = n83673 & n83917;
  assign n83972 = n83685 & n83924;
  assign n83973 = n83695 & n83923;
  assign n83974 = ~n83969 & ~n83970;
  assign n83975 = ~n83971 & n83974;
  assign n83976 = ~n83972 & n83975;
  assign n14941 = n83973 | ~n83976;
  assign n83978 = P2_P1_INSTQUEUE_REG_13__2_ & ~n83928;
  assign n83979 = n83713 & n83933;
  assign n83980 = n83715 & n83917;
  assign n83981 = n83729 & n83924;
  assign n83982 = n83743 & n83923;
  assign n83983 = ~n83978 & ~n83979;
  assign n83984 = ~n83980 & n83983;
  assign n83985 = ~n83981 & n83984;
  assign n14946 = n83982 | ~n83985;
  assign n83987 = P2_P1_INSTQUEUE_REG_13__1_ & ~n83928;
  assign n83988 = n83758 & n83933;
  assign n83989 = n83760 & n83917;
  assign n83990 = n83769 & n83924;
  assign n83991 = n83781 & n83923;
  assign n83992 = ~n83987 & ~n83988;
  assign n83993 = ~n83989 & n83992;
  assign n83994 = ~n83990 & n83993;
  assign n14951 = n83991 | ~n83994;
  assign n83996 = P2_P1_INSTQUEUE_REG_13__0_ & ~n83928;
  assign n83997 = n83791 & n83933;
  assign n83998 = n83793 & n83917;
  assign n83999 = n83806 & n83924;
  assign n84000 = n83820 & n83923;
  assign n84001 = ~n83996 & ~n83997;
  assign n84002 = ~n83998 & n84001;
  assign n84003 = ~n83999 & n84002;
  assign n14956 = n84000 | ~n84003;
  assign n84005 = P2_P1_INSTQUEUEWR_ADDR_REG_3_ & ~P2_P1_INSTQUEUEWR_ADDR_REG_1_;
  assign n84006 = n83827 & n84005;
  assign n84007 = P2_P1_STATE2_REG_3_ & ~n84006;
  assign n84008 = n77374 & ~n84007;
  assign n84009 = P2_P1_INSTQUEUEWR_ADDR_REG_0_ & n77397;
  assign n84010 = n77417 & n84009;
  assign n84011 = ~P2_P1_INSTQUEUEWR_ADDR_REG_0_ & n77394;
  assign n84012 = n77419 & n84011;
  assign n84013 = ~n84010 & ~n84012;
  assign n84014 = n77391 & ~n84013;
  assign n84015 = n77382 & n77385;
  assign n84016 = ~n84014 & ~n84015;
  assign n84017 = n84008 & ~n84016;
  assign n84018 = P2_P1_INSTQUEUE_REG_12__7_ & ~n84017;
  assign n84019 = n77427 & n84006;
  assign n84020 = n77429 & n84013;
  assign n84021 = n77391 & ~n84020;
  assign n84022 = n84015 & ~n84021;
  assign n84023 = n77701 & n84022;
  assign n84024 = n80593 & n84012;
  assign n84025 = ~n84018 & ~n84019;
  assign n84026 = ~n84023 & n84025;
  assign n84027 = ~n84024 & n84026;
  assign n84028 = ~n83519 & n84027;
  assign n84029 = ~n84010 & n84027;
  assign n14961 = ~n84028 & ~n84029;
  assign n84031 = P2_P1_INSTQUEUE_REG_12__6_ & ~n84017;
  assign n84032 = n83536 & n84022;
  assign n84033 = n83538 & n84006;
  assign n84034 = n83552 & n84012;
  assign n84035 = n83566 & n84010;
  assign n84036 = ~n84031 & ~n84032;
  assign n84037 = ~n84033 & n84036;
  assign n84038 = ~n84034 & n84037;
  assign n14966 = n84035 | ~n84038;
  assign n84040 = P2_P1_INSTQUEUE_REG_12__5_ & ~n84017;
  assign n84041 = n83583 & n84022;
  assign n84042 = n83585 & n84006;
  assign n84043 = n83596 & n84012;
  assign n84044 = n83608 & n84010;
  assign n84045 = ~n84040 & ~n84041;
  assign n84046 = ~n84042 & n84045;
  assign n84047 = ~n84043 & n84046;
  assign n14971 = n84044 | ~n84047;
  assign n84049 = P2_P1_INSTQUEUE_REG_12__4_ & ~n84017;
  assign n84050 = n83627 & n84022;
  assign n84051 = n83629 & n84006;
  assign n84052 = n83642 & n84012;
  assign n84053 = n83654 & n84010;
  assign n84054 = ~n84049 & ~n84050;
  assign n84055 = ~n84051 & n84054;
  assign n84056 = ~n84052 & n84055;
  assign n14976 = n84053 | ~n84056;
  assign n84058 = P2_P1_INSTQUEUE_REG_12__3_ & ~n84017;
  assign n84059 = n83671 & n84022;
  assign n84060 = n83673 & n84006;
  assign n84061 = n83685 & n84012;
  assign n84062 = n83695 & n84010;
  assign n84063 = ~n84058 & ~n84059;
  assign n84064 = ~n84060 & n84063;
  assign n84065 = ~n84061 & n84064;
  assign n14981 = n84062 | ~n84065;
  assign n84067 = P2_P1_INSTQUEUE_REG_12__2_ & ~n84017;
  assign n84068 = n83713 & n84022;
  assign n84069 = n83715 & n84006;
  assign n84070 = n83729 & n84012;
  assign n84071 = n83743 & n84010;
  assign n84072 = ~n84067 & ~n84068;
  assign n84073 = ~n84069 & n84072;
  assign n84074 = ~n84070 & n84073;
  assign n14986 = n84071 | ~n84074;
  assign n84076 = P2_P1_INSTQUEUE_REG_12__1_ & ~n84017;
  assign n84077 = n83758 & n84022;
  assign n84078 = n83760 & n84006;
  assign n84079 = n83769 & n84012;
  assign n84080 = n83781 & n84010;
  assign n84081 = ~n84076 & ~n84077;
  assign n84082 = ~n84078 & n84081;
  assign n84083 = ~n84079 & n84082;
  assign n14991 = n84080 | ~n84083;
  assign n84085 = P2_P1_INSTQUEUE_REG_12__0_ & ~n84017;
  assign n84086 = n83791 & n84022;
  assign n84087 = n83793 & n84006;
  assign n84088 = n83806 & n84012;
  assign n84089 = n83820 & n84010;
  assign n84090 = ~n84085 & ~n84086;
  assign n84091 = ~n84087 & n84090;
  assign n84092 = ~n84088 & n84091;
  assign n14996 = n84089 | ~n84092;
  assign n84094 = P2_P1_INSTQUEUEWR_ADDR_REG_3_ & ~P2_P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n84095 = n77367 & n84094;
  assign n84096 = P2_P1_STATE2_REG_3_ & ~n84095;
  assign n84097 = n77374 & ~n84096;
  assign n84098 = n77378 & ~n77381;
  assign n84099 = n77386 & n84098;
  assign n84100 = ~n84095 & ~n84099;
  assign n84101 = n77405 & ~n77416;
  assign n84102 = n77398 & n84101;
  assign n84103 = n77402 & n77411;
  assign n84104 = ~n84102 & ~n84103;
  assign n84105 = n77391 & ~n84104;
  assign n84106 = n84100 & ~n84105;
  assign n84107 = n84097 & ~n84106;
  assign n84108 = P2_P1_INSTQUEUE_REG_11__7_ & ~n84107;
  assign n84109 = n77427 & n84095;
  assign n84110 = n77429 & n84104;
  assign n84111 = n77391 & ~n84110;
  assign n84112 = ~n84100 & ~n84111;
  assign n84113 = n77701 & n84112;
  assign n84114 = n80593 & n84103;
  assign n84115 = ~n84108 & ~n84109;
  assign n84116 = ~n84113 & n84115;
  assign n84117 = ~n84114 & n84116;
  assign n84118 = ~n83519 & n84117;
  assign n84119 = ~n84102 & n84117;
  assign n15001 = ~n84118 & ~n84119;
  assign n84121 = P2_P1_INSTQUEUE_REG_11__6_ & ~n84107;
  assign n84122 = n83536 & n84112;
  assign n84123 = n83538 & n84095;
  assign n84124 = n83552 & n84103;
  assign n84125 = n83566 & n84102;
  assign n84126 = ~n84121 & ~n84122;
  assign n84127 = ~n84123 & n84126;
  assign n84128 = ~n84124 & n84127;
  assign n15006 = n84125 | ~n84128;
  assign n84130 = P2_P1_INSTQUEUE_REG_11__5_ & ~n84107;
  assign n84131 = n83583 & n84112;
  assign n84132 = n83585 & n84095;
  assign n84133 = n83596 & n84103;
  assign n84134 = n83608 & n84102;
  assign n84135 = ~n84130 & ~n84131;
  assign n84136 = ~n84132 & n84135;
  assign n84137 = ~n84133 & n84136;
  assign n15011 = n84134 | ~n84137;
  assign n84139 = P2_P1_INSTQUEUE_REG_11__4_ & ~n84107;
  assign n84140 = n83627 & n84112;
  assign n84141 = n83629 & n84095;
  assign n84142 = n83642 & n84103;
  assign n84143 = n83654 & n84102;
  assign n84144 = ~n84139 & ~n84140;
  assign n84145 = ~n84141 & n84144;
  assign n84146 = ~n84142 & n84145;
  assign n15016 = n84143 | ~n84146;
  assign n84148 = P2_P1_INSTQUEUE_REG_11__3_ & ~n84107;
  assign n84149 = n83671 & n84112;
  assign n84150 = n83673 & n84095;
  assign n84151 = n83685 & n84103;
  assign n84152 = n83695 & n84102;
  assign n84153 = ~n84148 & ~n84149;
  assign n84154 = ~n84150 & n84153;
  assign n84155 = ~n84151 & n84154;
  assign n15021 = n84152 | ~n84155;
  assign n84157 = P2_P1_INSTQUEUE_REG_11__2_ & ~n84107;
  assign n84158 = n83713 & n84112;
  assign n84159 = n83715 & n84095;
  assign n84160 = n83729 & n84103;
  assign n84161 = n83743 & n84102;
  assign n84162 = ~n84157 & ~n84158;
  assign n84163 = ~n84159 & n84162;
  assign n84164 = ~n84160 & n84163;
  assign n15026 = n84161 | ~n84164;
  assign n84166 = P2_P1_INSTQUEUE_REG_11__1_ & ~n84107;
  assign n84167 = n83758 & n84112;
  assign n84168 = n83760 & n84095;
  assign n84169 = n83769 & n84103;
  assign n84170 = n83781 & n84102;
  assign n84171 = ~n84166 & ~n84167;
  assign n84172 = ~n84168 & n84171;
  assign n84173 = ~n84169 & n84172;
  assign n15031 = n84170 | ~n84173;
  assign n84175 = P2_P1_INSTQUEUE_REG_11__0_ & ~n84107;
  assign n84176 = n83791 & n84112;
  assign n84177 = n83793 & n84095;
  assign n84178 = n83806 & n84103;
  assign n84179 = n83820 & n84102;
  assign n84180 = ~n84175 & ~n84176;
  assign n84181 = ~n84177 & n84180;
  assign n84182 = ~n84178 & n84181;
  assign n15036 = n84179 | ~n84182;
  assign n84184 = ~P2_P1_INSTQUEUEWR_ADDR_REG_2_ & ~P2_P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n84185 = n83826 & n84184;
  assign n84186 = P2_P1_STATE2_REG_3_ & ~n84185;
  assign n84187 = n77374 & ~n84186;
  assign n84188 = n77392 & n84098;
  assign n84189 = ~n84185 & ~n84188;
  assign n84190 = n83833 & n84101;
  assign n84191 = n77395 & n77411;
  assign n84192 = ~n84190 & ~n84191;
  assign n84193 = n77391 & ~n84192;
  assign n84194 = n84189 & ~n84193;
  assign n84195 = n84187 & ~n84194;
  assign n84196 = P2_P1_INSTQUEUE_REG_10__7_ & ~n84195;
  assign n84197 = n77427 & n84185;
  assign n84198 = n77429 & n84192;
  assign n84199 = n77391 & ~n84198;
  assign n84200 = ~n84189 & ~n84199;
  assign n84201 = n77701 & n84200;
  assign n84202 = n80593 & n84191;
  assign n84203 = ~n84196 & ~n84197;
  assign n84204 = ~n84201 & n84203;
  assign n84205 = ~n84202 & n84204;
  assign n84206 = ~n83519 & n84205;
  assign n84207 = ~n84190 & n84205;
  assign n15041 = ~n84206 & ~n84207;
  assign n84209 = P2_P1_INSTQUEUE_REG_10__6_ & ~n84195;
  assign n84210 = n83536 & n84200;
  assign n84211 = n83538 & n84185;
  assign n84212 = n83552 & n84191;
  assign n84213 = n83566 & n84190;
  assign n84214 = ~n84209 & ~n84210;
  assign n84215 = ~n84211 & n84214;
  assign n84216 = ~n84212 & n84215;
  assign n15046 = n84213 | ~n84216;
  assign n84218 = P2_P1_INSTQUEUE_REG_10__5_ & ~n84195;
  assign n84219 = n83583 & n84200;
  assign n84220 = n83585 & n84185;
  assign n84221 = n83596 & n84191;
  assign n84222 = n83608 & n84190;
  assign n84223 = ~n84218 & ~n84219;
  assign n84224 = ~n84220 & n84223;
  assign n84225 = ~n84221 & n84224;
  assign n15051 = n84222 | ~n84225;
  assign n84227 = P2_P1_INSTQUEUE_REG_10__4_ & ~n84195;
  assign n84228 = n83627 & n84200;
  assign n84229 = n83629 & n84185;
  assign n84230 = n83642 & n84191;
  assign n84231 = n83654 & n84190;
  assign n84232 = ~n84227 & ~n84228;
  assign n84233 = ~n84229 & n84232;
  assign n84234 = ~n84230 & n84233;
  assign n15056 = n84231 | ~n84234;
  assign n84236 = P2_P1_INSTQUEUE_REG_10__3_ & ~n84195;
  assign n84237 = n83671 & n84200;
  assign n84238 = n83673 & n84185;
  assign n84239 = n83685 & n84191;
  assign n84240 = n83695 & n84190;
  assign n84241 = ~n84236 & ~n84237;
  assign n84242 = ~n84238 & n84241;
  assign n84243 = ~n84239 & n84242;
  assign n15061 = n84240 | ~n84243;
  assign n84245 = P2_P1_INSTQUEUE_REG_10__2_ & ~n84195;
  assign n84246 = n83713 & n84200;
  assign n84247 = n83715 & n84185;
  assign n84248 = n83729 & n84191;
  assign n84249 = n83743 & n84190;
  assign n84250 = ~n84245 & ~n84246;
  assign n84251 = ~n84247 & n84250;
  assign n84252 = ~n84248 & n84251;
  assign n15066 = n84249 | ~n84252;
  assign n84254 = P2_P1_INSTQUEUE_REG_10__1_ & ~n84195;
  assign n84255 = n83758 & n84200;
  assign n84256 = n83760 & n84185;
  assign n84257 = n83769 & n84191;
  assign n84258 = n83781 & n84190;
  assign n84259 = ~n84254 & ~n84255;
  assign n84260 = ~n84256 & n84259;
  assign n84261 = ~n84257 & n84260;
  assign n15071 = n84258 | ~n84261;
  assign n84263 = P2_P1_INSTQUEUE_REG_10__0_ & ~n84195;
  assign n84264 = n83791 & n84200;
  assign n84265 = n83793 & n84185;
  assign n84266 = n83806 & n84191;
  assign n84267 = n83820 & n84190;
  assign n84268 = ~n84263 & ~n84264;
  assign n84269 = ~n84265 & n84268;
  assign n84270 = ~n84266 & n84269;
  assign n15076 = n84267 | ~n84270;
  assign n84272 = n77383 & n84094;
  assign n84273 = P2_P1_STATE2_REG_3_ & ~n84272;
  assign n84274 = n77374 & ~n84273;
  assign n84275 = n77393 & n84098;
  assign n84276 = ~n84272 & ~n84275;
  assign n84277 = n83922 & n84101;
  assign n84278 = n77396 & n77411;
  assign n84279 = ~n84277 & ~n84278;
  assign n84280 = n77391 & ~n84279;
  assign n84281 = n84276 & ~n84280;
  assign n84282 = n84274 & ~n84281;
  assign n84283 = P2_P1_INSTQUEUE_REG_9__7_ & ~n84282;
  assign n84284 = n77427 & n84272;
  assign n84285 = n77429 & n84279;
  assign n84286 = n77391 & ~n84285;
  assign n84287 = ~n84276 & ~n84286;
  assign n84288 = n77701 & n84287;
  assign n84289 = n80593 & n84278;
  assign n84290 = ~n84283 & ~n84284;
  assign n84291 = ~n84288 & n84290;
  assign n84292 = ~n84289 & n84291;
  assign n84293 = ~n83519 & n84292;
  assign n84294 = ~n84277 & n84292;
  assign n15081 = ~n84293 & ~n84294;
  assign n84296 = P2_P1_INSTQUEUE_REG_9__6_ & ~n84282;
  assign n84297 = n83536 & n84287;
  assign n84298 = n83538 & n84272;
  assign n84299 = n83552 & n84278;
  assign n84300 = n83566 & n84277;
  assign n84301 = ~n84296 & ~n84297;
  assign n84302 = ~n84298 & n84301;
  assign n84303 = ~n84299 & n84302;
  assign n15086 = n84300 | ~n84303;
  assign n84305 = P2_P1_INSTQUEUE_REG_9__5_ & ~n84282;
  assign n84306 = n83583 & n84287;
  assign n84307 = n83585 & n84272;
  assign n84308 = n83596 & n84278;
  assign n84309 = n83608 & n84277;
  assign n84310 = ~n84305 & ~n84306;
  assign n84311 = ~n84307 & n84310;
  assign n84312 = ~n84308 & n84311;
  assign n15091 = n84309 | ~n84312;
  assign n84314 = P2_P1_INSTQUEUE_REG_9__4_ & ~n84282;
  assign n84315 = n83627 & n84287;
  assign n84316 = n83629 & n84272;
  assign n84317 = n83642 & n84278;
  assign n84318 = n83654 & n84277;
  assign n84319 = ~n84314 & ~n84315;
  assign n84320 = ~n84316 & n84319;
  assign n84321 = ~n84317 & n84320;
  assign n15096 = n84318 | ~n84321;
  assign n84323 = P2_P1_INSTQUEUE_REG_9__3_ & ~n84282;
  assign n84324 = n83671 & n84287;
  assign n84325 = n83673 & n84272;
  assign n84326 = n83685 & n84278;
  assign n84327 = n83695 & n84277;
  assign n84328 = ~n84323 & ~n84324;
  assign n84329 = ~n84325 & n84328;
  assign n84330 = ~n84326 & n84329;
  assign n15101 = n84327 | ~n84330;
  assign n84332 = P2_P1_INSTQUEUE_REG_9__2_ & ~n84282;
  assign n84333 = n83713 & n84287;
  assign n84334 = n83715 & n84272;
  assign n84335 = n83729 & n84278;
  assign n84336 = n83743 & n84277;
  assign n84337 = ~n84332 & ~n84333;
  assign n84338 = ~n84334 & n84337;
  assign n84339 = ~n84335 & n84338;
  assign n15106 = n84336 | ~n84339;
  assign n84341 = P2_P1_INSTQUEUE_REG_9__1_ & ~n84282;
  assign n84342 = n83758 & n84287;
  assign n84343 = n83760 & n84272;
  assign n84344 = n83769 & n84278;
  assign n84345 = n83781 & n84277;
  assign n84346 = ~n84341 & ~n84342;
  assign n84347 = ~n84343 & n84346;
  assign n84348 = ~n84344 & n84347;
  assign n15111 = n84345 | ~n84348;
  assign n84350 = P2_P1_INSTQUEUE_REG_9__0_ & ~n84282;
  assign n84351 = n83791 & n84287;
  assign n84352 = n83793 & n84272;
  assign n84353 = n83806 & n84278;
  assign n84354 = n83820 & n84277;
  assign n84355 = ~n84350 & ~n84351;
  assign n84356 = ~n84352 & n84355;
  assign n84357 = ~n84353 & n84356;
  assign n15116 = n84354 | ~n84357;
  assign n84359 = n84005 & n84184;
  assign n84360 = P2_P1_STATE2_REG_3_ & ~n84359;
  assign n84361 = n77374 & ~n84360;
  assign n84362 = n84009 & n84101;
  assign n84363 = n77411 & n84011;
  assign n84364 = ~n84362 & ~n84363;
  assign n84365 = n77391 & ~n84364;
  assign n84366 = n77385 & n84098;
  assign n84367 = ~n84365 & ~n84366;
  assign n84368 = n84361 & ~n84367;
  assign n84369 = P2_P1_INSTQUEUE_REG_8__7_ & ~n84368;
  assign n84370 = n77427 & n84359;
  assign n84371 = n77429 & n84364;
  assign n84372 = n77391 & ~n84371;
  assign n84373 = n84366 & ~n84372;
  assign n84374 = n77701 & n84373;
  assign n84375 = n80593 & n84363;
  assign n84376 = ~n84369 & ~n84370;
  assign n84377 = ~n84374 & n84376;
  assign n84378 = ~n84375 & n84377;
  assign n84379 = ~n83519 & n84378;
  assign n84380 = ~n84362 & n84378;
  assign n15121 = ~n84379 & ~n84380;
  assign n84382 = P2_P1_INSTQUEUE_REG_8__6_ & ~n84368;
  assign n84383 = n83536 & n84373;
  assign n84384 = n83538 & n84359;
  assign n84385 = n83552 & n84363;
  assign n84386 = n83566 & n84362;
  assign n84387 = ~n84382 & ~n84383;
  assign n84388 = ~n84384 & n84387;
  assign n84389 = ~n84385 & n84388;
  assign n15126 = n84386 | ~n84389;
  assign n84391 = P2_P1_INSTQUEUE_REG_8__5_ & ~n84368;
  assign n84392 = n83583 & n84373;
  assign n84393 = n83585 & n84359;
  assign n84394 = n83596 & n84363;
  assign n84395 = n83608 & n84362;
  assign n84396 = ~n84391 & ~n84392;
  assign n84397 = ~n84393 & n84396;
  assign n84398 = ~n84394 & n84397;
  assign n15131 = n84395 | ~n84398;
  assign n84400 = P2_P1_INSTQUEUE_REG_8__4_ & ~n84368;
  assign n84401 = n83627 & n84373;
  assign n84402 = n83629 & n84359;
  assign n84403 = n83642 & n84363;
  assign n84404 = n83654 & n84362;
  assign n84405 = ~n84400 & ~n84401;
  assign n84406 = ~n84402 & n84405;
  assign n84407 = ~n84403 & n84406;
  assign n15136 = n84404 | ~n84407;
  assign n84409 = P2_P1_INSTQUEUE_REG_8__3_ & ~n84368;
  assign n84410 = n83671 & n84373;
  assign n84411 = n83673 & n84359;
  assign n84412 = n83685 & n84363;
  assign n84413 = n83695 & n84362;
  assign n84414 = ~n84409 & ~n84410;
  assign n84415 = ~n84411 & n84414;
  assign n84416 = ~n84412 & n84415;
  assign n15141 = n84413 | ~n84416;
  assign n84418 = P2_P1_INSTQUEUE_REG_8__2_ & ~n84368;
  assign n84419 = n83713 & n84373;
  assign n84420 = n83715 & n84359;
  assign n84421 = n83729 & n84363;
  assign n84422 = n83743 & n84362;
  assign n84423 = ~n84418 & ~n84419;
  assign n84424 = ~n84420 & n84423;
  assign n84425 = ~n84421 & n84424;
  assign n15146 = n84422 | ~n84425;
  assign n84427 = P2_P1_INSTQUEUE_REG_8__1_ & ~n84368;
  assign n84428 = n83758 & n84373;
  assign n84429 = n83760 & n84359;
  assign n84430 = n83769 & n84363;
  assign n84431 = n83781 & n84362;
  assign n84432 = ~n84427 & ~n84428;
  assign n84433 = ~n84429 & n84432;
  assign n84434 = ~n84430 & n84433;
  assign n15151 = n84431 | ~n84434;
  assign n84436 = P2_P1_INSTQUEUE_REG_8__0_ & ~n84368;
  assign n84437 = n83791 & n84373;
  assign n84438 = n83793 & n84359;
  assign n84439 = n83806 & n84363;
  assign n84440 = n83820 & n84362;
  assign n84441 = ~n84436 & ~n84437;
  assign n84442 = ~n84438 & n84441;
  assign n84443 = ~n84439 & n84442;
  assign n15156 = n84440 | ~n84443;
  assign n84445 = P2_P1_STATE2_REG_3_ & ~n77379;
  assign n84446 = n77374 & ~n84445;
  assign n84447 = ~n77379 & ~n77407;
  assign n84448 = ~n77405 & n77416;
  assign n84449 = n77398 & n84448;
  assign n84450 = ~n77415 & ~n84449;
  assign n84451 = n77391 & ~n84450;
  assign n84452 = n84447 & ~n84451;
  assign n84453 = n84446 & ~n84452;
  assign n84454 = P2_P1_INSTQUEUE_REG_7__7_ & ~n84453;
  assign n84455 = n77379 & n77427;
  assign n84456 = n77429 & n84450;
  assign n84457 = n77391 & ~n84456;
  assign n84458 = ~n84447 & ~n84457;
  assign n84459 = n77701 & n84458;
  assign n84460 = n77415 & n80593;
  assign n84461 = ~n84454 & ~n84455;
  assign n84462 = ~n84459 & n84461;
  assign n84463 = ~n84460 & n84462;
  assign n84464 = ~n83519 & n84463;
  assign n84465 = ~n84449 & n84463;
  assign n15161 = ~n84464 & ~n84465;
  assign n84467 = P2_P1_INSTQUEUE_REG_7__6_ & ~n84453;
  assign n84468 = n83536 & n84458;
  assign n84469 = n77379 & n83538;
  assign n84470 = n77415 & n83552;
  assign n84471 = n83566 & n84449;
  assign n84472 = ~n84467 & ~n84468;
  assign n84473 = ~n84469 & n84472;
  assign n84474 = ~n84470 & n84473;
  assign n15166 = n84471 | ~n84474;
  assign n84476 = P2_P1_INSTQUEUE_REG_7__5_ & ~n84453;
  assign n84477 = n83583 & n84458;
  assign n84478 = n77379 & n83585;
  assign n84479 = n77415 & n83596;
  assign n84480 = n83608 & n84449;
  assign n84481 = ~n84476 & ~n84477;
  assign n84482 = ~n84478 & n84481;
  assign n84483 = ~n84479 & n84482;
  assign n15171 = n84480 | ~n84483;
  assign n84485 = P2_P1_INSTQUEUE_REG_7__4_ & ~n84453;
  assign n84486 = n83627 & n84458;
  assign n84487 = n77379 & n83629;
  assign n84488 = n77415 & n83642;
  assign n84489 = n83654 & n84449;
  assign n84490 = ~n84485 & ~n84486;
  assign n84491 = ~n84487 & n84490;
  assign n84492 = ~n84488 & n84491;
  assign n15176 = n84489 | ~n84492;
  assign n84494 = P2_P1_INSTQUEUE_REG_7__3_ & ~n84453;
  assign n84495 = n83671 & n84458;
  assign n84496 = n77379 & n83673;
  assign n84497 = n77415 & n83685;
  assign n84498 = n83695 & n84449;
  assign n84499 = ~n84494 & ~n84495;
  assign n84500 = ~n84496 & n84499;
  assign n84501 = ~n84497 & n84500;
  assign n15181 = n84498 | ~n84501;
  assign n84503 = P2_P1_INSTQUEUE_REG_7__2_ & ~n84453;
  assign n84504 = n83713 & n84458;
  assign n84505 = n77379 & n83715;
  assign n84506 = n77415 & n83729;
  assign n84507 = n83743 & n84449;
  assign n84508 = ~n84503 & ~n84504;
  assign n84509 = ~n84505 & n84508;
  assign n84510 = ~n84506 & n84509;
  assign n15186 = n84507 | ~n84510;
  assign n84512 = P2_P1_INSTQUEUE_REG_7__1_ & ~n84453;
  assign n84513 = n83758 & n84458;
  assign n84514 = n77379 & n83760;
  assign n84515 = n77415 & n83769;
  assign n84516 = n83781 & n84449;
  assign n84517 = ~n84512 & ~n84513;
  assign n84518 = ~n84514 & n84517;
  assign n84519 = ~n84515 & n84518;
  assign n15191 = n84516 | ~n84519;
  assign n84521 = P2_P1_INSTQUEUE_REG_7__0_ & ~n84453;
  assign n84522 = n83791 & n84458;
  assign n84523 = n77379 & n83793;
  assign n84524 = n77415 & n83806;
  assign n84525 = n83820 & n84449;
  assign n84526 = ~n84521 & ~n84522;
  assign n84527 = ~n84523 & n84526;
  assign n84528 = ~n84524 & n84527;
  assign n15196 = n84525 | ~n84528;
  assign n84530 = ~P2_P1_INSTQUEUEWR_ADDR_REG_3_ & P2_P1_INSTQUEUEWR_ADDR_REG_1_;
  assign n84531 = n83827 & n84530;
  assign n84532 = P2_P1_STATE2_REG_3_ & ~n84531;
  assign n84533 = n77374 & ~n84532;
  assign n84534 = n77392 & n77406;
  assign n84535 = ~n84531 & ~n84534;
  assign n84536 = n83833 & n84448;
  assign n84537 = n77395 & n77414;
  assign n84538 = ~n84536 & ~n84537;
  assign n84539 = n77391 & ~n84538;
  assign n84540 = n84535 & ~n84539;
  assign n84541 = n84533 & ~n84540;
  assign n84542 = P2_P1_INSTQUEUE_REG_6__7_ & ~n84541;
  assign n84543 = n77427 & n84531;
  assign n84544 = n77429 & n84538;
  assign n84545 = n77391 & ~n84544;
  assign n84546 = ~n84535 & ~n84545;
  assign n84547 = n77701 & n84546;
  assign n84548 = n80593 & n84537;
  assign n84549 = ~n84542 & ~n84543;
  assign n84550 = ~n84547 & n84549;
  assign n84551 = ~n84548 & n84550;
  assign n84552 = ~n83519 & n84551;
  assign n84553 = ~n84536 & n84551;
  assign n15201 = ~n84552 & ~n84553;
  assign n84555 = P2_P1_INSTQUEUE_REG_6__6_ & ~n84541;
  assign n84556 = n83536 & n84546;
  assign n84557 = n83538 & n84531;
  assign n84558 = n83552 & n84537;
  assign n84559 = n83566 & n84536;
  assign n84560 = ~n84555 & ~n84556;
  assign n84561 = ~n84557 & n84560;
  assign n84562 = ~n84558 & n84561;
  assign n15206 = n84559 | ~n84562;
  assign n84564 = P2_P1_INSTQUEUE_REG_6__5_ & ~n84541;
  assign n84565 = n83583 & n84546;
  assign n84566 = n83585 & n84531;
  assign n84567 = n83596 & n84537;
  assign n84568 = n83608 & n84536;
  assign n84569 = ~n84564 & ~n84565;
  assign n84570 = ~n84566 & n84569;
  assign n84571 = ~n84567 & n84570;
  assign n15211 = n84568 | ~n84571;
  assign n84573 = P2_P1_INSTQUEUE_REG_6__4_ & ~n84541;
  assign n84574 = n83627 & n84546;
  assign n84575 = n83629 & n84531;
  assign n84576 = n83642 & n84537;
  assign n84577 = n83654 & n84536;
  assign n84578 = ~n84573 & ~n84574;
  assign n84579 = ~n84575 & n84578;
  assign n84580 = ~n84576 & n84579;
  assign n15216 = n84577 | ~n84580;
  assign n84582 = P2_P1_INSTQUEUE_REG_6__3_ & ~n84541;
  assign n84583 = n83671 & n84546;
  assign n84584 = n83673 & n84531;
  assign n84585 = n83685 & n84537;
  assign n84586 = n83695 & n84536;
  assign n84587 = ~n84582 & ~n84583;
  assign n84588 = ~n84584 & n84587;
  assign n84589 = ~n84585 & n84588;
  assign n15221 = n84586 | ~n84589;
  assign n84591 = P2_P1_INSTQUEUE_REG_6__2_ & ~n84541;
  assign n84592 = n83713 & n84546;
  assign n84593 = n83715 & n84531;
  assign n84594 = n83729 & n84537;
  assign n84595 = n83743 & n84536;
  assign n84596 = ~n84591 & ~n84592;
  assign n84597 = ~n84593 & n84596;
  assign n84598 = ~n84594 & n84597;
  assign n15226 = n84595 | ~n84598;
  assign n84600 = P2_P1_INSTQUEUE_REG_6__1_ & ~n84541;
  assign n84601 = n83758 & n84546;
  assign n84602 = n83760 & n84531;
  assign n84603 = n83769 & n84537;
  assign n84604 = n83781 & n84536;
  assign n84605 = ~n84600 & ~n84601;
  assign n84606 = ~n84602 & n84605;
  assign n84607 = ~n84603 & n84606;
  assign n15231 = n84604 | ~n84607;
  assign n84609 = P2_P1_INSTQUEUE_REG_6__0_ & ~n84541;
  assign n84610 = n83791 & n84546;
  assign n84611 = n83793 & n84531;
  assign n84612 = n83806 & n84537;
  assign n84613 = n83820 & n84536;
  assign n84614 = ~n84609 & ~n84610;
  assign n84615 = ~n84611 & n84614;
  assign n84616 = ~n84612 & n84615;
  assign n15236 = n84613 | ~n84616;
  assign n84618 = ~P2_P1_INSTQUEUEWR_ADDR_REG_3_ & P2_P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n84619 = n77383 & n84618;
  assign n84620 = P2_P1_STATE2_REG_3_ & ~n84619;
  assign n84621 = n77374 & ~n84620;
  assign n84622 = n77393 & n77406;
  assign n84623 = ~n84619 & ~n84622;
  assign n84624 = n83922 & n84448;
  assign n84625 = n77396 & n77414;
  assign n84626 = ~n84624 & ~n84625;
  assign n84627 = n77391 & ~n84626;
  assign n84628 = n84623 & ~n84627;
  assign n84629 = n84621 & ~n84628;
  assign n84630 = P2_P1_INSTQUEUE_REG_5__7_ & ~n84629;
  assign n84631 = n77427 & n84619;
  assign n84632 = n77429 & n84626;
  assign n84633 = n77391 & ~n84632;
  assign n84634 = ~n84623 & ~n84633;
  assign n84635 = n77701 & n84634;
  assign n84636 = n80593 & n84625;
  assign n84637 = ~n84630 & ~n84631;
  assign n84638 = ~n84635 & n84637;
  assign n84639 = ~n84636 & n84638;
  assign n84640 = ~n83519 & n84639;
  assign n84641 = ~n84624 & n84639;
  assign n15241 = ~n84640 & ~n84641;
  assign n84643 = P2_P1_INSTQUEUE_REG_5__6_ & ~n84629;
  assign n84644 = n83536 & n84634;
  assign n84645 = n83538 & n84619;
  assign n84646 = n83552 & n84625;
  assign n84647 = n83566 & n84624;
  assign n84648 = ~n84643 & ~n84644;
  assign n84649 = ~n84645 & n84648;
  assign n84650 = ~n84646 & n84649;
  assign n15246 = n84647 | ~n84650;
  assign n84652 = P2_P1_INSTQUEUE_REG_5__5_ & ~n84629;
  assign n84653 = n83583 & n84634;
  assign n84654 = n83585 & n84619;
  assign n84655 = n83596 & n84625;
  assign n84656 = n83608 & n84624;
  assign n84657 = ~n84652 & ~n84653;
  assign n84658 = ~n84654 & n84657;
  assign n84659 = ~n84655 & n84658;
  assign n15251 = n84656 | ~n84659;
  assign n84661 = P2_P1_INSTQUEUE_REG_5__4_ & ~n84629;
  assign n84662 = n83627 & n84634;
  assign n84663 = n83629 & n84619;
  assign n84664 = n83642 & n84625;
  assign n84665 = n83654 & n84624;
  assign n84666 = ~n84661 & ~n84662;
  assign n84667 = ~n84663 & n84666;
  assign n84668 = ~n84664 & n84667;
  assign n15256 = n84665 | ~n84668;
  assign n84670 = P2_P1_INSTQUEUE_REG_5__3_ & ~n84629;
  assign n84671 = n83671 & n84634;
  assign n84672 = n83673 & n84619;
  assign n84673 = n83685 & n84625;
  assign n84674 = n83695 & n84624;
  assign n84675 = ~n84670 & ~n84671;
  assign n84676 = ~n84672 & n84675;
  assign n84677 = ~n84673 & n84676;
  assign n15261 = n84674 | ~n84677;
  assign n84679 = P2_P1_INSTQUEUE_REG_5__2_ & ~n84629;
  assign n84680 = n83713 & n84634;
  assign n84681 = n83715 & n84619;
  assign n84682 = n83729 & n84625;
  assign n84683 = n83743 & n84624;
  assign n84684 = ~n84679 & ~n84680;
  assign n84685 = ~n84681 & n84684;
  assign n84686 = ~n84682 & n84685;
  assign n15266 = n84683 | ~n84686;
  assign n84688 = P2_P1_INSTQUEUE_REG_5__1_ & ~n84629;
  assign n84689 = n83758 & n84634;
  assign n84690 = n83760 & n84619;
  assign n84691 = n83769 & n84625;
  assign n84692 = n83781 & n84624;
  assign n84693 = ~n84688 & ~n84689;
  assign n84694 = ~n84690 & n84693;
  assign n84695 = ~n84691 & n84694;
  assign n15271 = n84692 | ~n84695;
  assign n84697 = P2_P1_INSTQUEUE_REG_5__0_ & ~n84629;
  assign n84698 = n83791 & n84634;
  assign n84699 = n83793 & n84619;
  assign n84700 = n83806 & n84625;
  assign n84701 = n83820 & n84624;
  assign n84702 = ~n84697 & ~n84698;
  assign n84703 = ~n84699 & n84702;
  assign n84704 = ~n84700 & n84703;
  assign n15276 = n84701 | ~n84704;
  assign n84706 = ~P2_P1_INSTQUEUEWR_ADDR_REG_3_ & ~P2_P1_INSTQUEUEWR_ADDR_REG_1_;
  assign n84707 = n83827 & n84706;
  assign n84708 = P2_P1_STATE2_REG_3_ & ~n84707;
  assign n84709 = n77374 & ~n84708;
  assign n84710 = n84009 & n84448;
  assign n84711 = n77414 & n84011;
  assign n84712 = ~n84710 & ~n84711;
  assign n84713 = n77391 & ~n84712;
  assign n84714 = n77385 & n77406;
  assign n84715 = ~n84713 & ~n84714;
  assign n84716 = n84709 & ~n84715;
  assign n84717 = P2_P1_INSTQUEUE_REG_4__7_ & ~n84716;
  assign n84718 = n77427 & n84707;
  assign n84719 = n77391 & ~n77429;
  assign n84720 = n84714 & ~n84719;
  assign n84721 = n77701 & n84720;
  assign n84722 = n80593 & n84711;
  assign n84723 = ~n84717 & ~n84718;
  assign n84724 = ~n84721 & n84723;
  assign n84725 = ~n84722 & n84724;
  assign n84726 = ~n83519 & n84725;
  assign n84727 = ~n84710 & n84725;
  assign n15281 = ~n84726 & ~n84727;
  assign n84729 = P2_P1_INSTQUEUE_REG_4__6_ & ~n84716;
  assign n84730 = n83536 & n84720;
  assign n84731 = n83538 & n84707;
  assign n84732 = n83552 & n84711;
  assign n84733 = n83566 & n84710;
  assign n84734 = ~n84729 & ~n84730;
  assign n84735 = ~n84731 & n84734;
  assign n84736 = ~n84732 & n84735;
  assign n15286 = n84733 | ~n84736;
  assign n84738 = P2_P1_INSTQUEUE_REG_4__5_ & ~n84716;
  assign n84739 = n83583 & n84720;
  assign n84740 = n83585 & n84707;
  assign n84741 = n83596 & n84711;
  assign n84742 = n83608 & n84710;
  assign n84743 = ~n84738 & ~n84739;
  assign n84744 = ~n84740 & n84743;
  assign n84745 = ~n84741 & n84744;
  assign n15291 = n84742 | ~n84745;
  assign n84747 = P2_P1_INSTQUEUE_REG_4__4_ & ~n84716;
  assign n84748 = n83627 & n84720;
  assign n84749 = n83629 & n84707;
  assign n84750 = n83642 & n84711;
  assign n84751 = n83654 & n84710;
  assign n84752 = ~n84747 & ~n84748;
  assign n84753 = ~n84749 & n84752;
  assign n84754 = ~n84750 & n84753;
  assign n15296 = n84751 | ~n84754;
  assign n84756 = P2_P1_INSTQUEUE_REG_4__3_ & ~n84716;
  assign n84757 = n83671 & n84720;
  assign n84758 = n83673 & n84707;
  assign n84759 = n83685 & n84711;
  assign n84760 = n83695 & n84710;
  assign n84761 = ~n84756 & ~n84757;
  assign n84762 = ~n84758 & n84761;
  assign n84763 = ~n84759 & n84762;
  assign n15301 = n84760 | ~n84763;
  assign n84765 = P2_P1_INSTQUEUE_REG_4__2_ & ~n84716;
  assign n84766 = n83713 & n84720;
  assign n84767 = n83715 & n84707;
  assign n84768 = n83729 & n84711;
  assign n84769 = n83743 & n84710;
  assign n84770 = ~n84765 & ~n84766;
  assign n84771 = ~n84767 & n84770;
  assign n84772 = ~n84768 & n84771;
  assign n15306 = n84769 | ~n84772;
  assign n84774 = P2_P1_INSTQUEUE_REG_4__1_ & ~n84716;
  assign n84775 = n83758 & n84720;
  assign n84776 = n83760 & n84707;
  assign n84777 = n83769 & n84711;
  assign n84778 = n83781 & n84710;
  assign n84779 = ~n84774 & ~n84775;
  assign n84780 = ~n84776 & n84779;
  assign n84781 = ~n84777 & n84780;
  assign n15311 = n84778 | ~n84781;
  assign n84783 = P2_P1_INSTQUEUE_REG_4__0_ & ~n84716;
  assign n84784 = n83791 & n84720;
  assign n84785 = n83793 & n84707;
  assign n84786 = n83806 & n84711;
  assign n84787 = n83820 & n84710;
  assign n84788 = ~n84783 & ~n84784;
  assign n84789 = ~n84785 & n84788;
  assign n84790 = ~n84786 & n84789;
  assign n15316 = n84787 | ~n84790;
  assign n84792 = ~P2_P1_INSTQUEUEWR_ADDR_REG_3_ & ~P2_P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n84793 = n77367 & n84792;
  assign n84794 = P2_P1_STATE2_REG_3_ & ~n84793;
  assign n84795 = n77374 & ~n84794;
  assign n84796 = n77378 & n77381;
  assign n84797 = n77386 & n84796;
  assign n84798 = ~n84793 & ~n84797;
  assign n84799 = n77405 & n77416;
  assign n84800 = n77398 & n84799;
  assign n84801 = n77401 & n77410;
  assign n84802 = n77402 & n84801;
  assign n84803 = ~n84800 & ~n84802;
  assign n84804 = n77391 & ~n84803;
  assign n84805 = n84798 & ~n84804;
  assign n84806 = n84795 & ~n84805;
  assign n84807 = P2_P1_INSTQUEUE_REG_3__7_ & ~n84806;
  assign n84808 = n77427 & n84793;
  assign n84809 = ~n84719 & ~n84798;
  assign n84810 = n77701 & n84809;
  assign n84811 = n80593 & n84802;
  assign n84812 = ~n84807 & ~n84808;
  assign n84813 = ~n84810 & n84812;
  assign n84814 = ~n84811 & n84813;
  assign n84815 = ~n83519 & n84814;
  assign n84816 = ~n84800 & n84814;
  assign n15321 = ~n84815 & ~n84816;
  assign n84818 = P2_P1_INSTQUEUE_REG_3__6_ & ~n84806;
  assign n84819 = n83536 & n84809;
  assign n84820 = n83538 & n84793;
  assign n84821 = n83552 & n84802;
  assign n84822 = n83566 & n84800;
  assign n84823 = ~n84818 & ~n84819;
  assign n84824 = ~n84820 & n84823;
  assign n84825 = ~n84821 & n84824;
  assign n15326 = n84822 | ~n84825;
  assign n84827 = P2_P1_INSTQUEUE_REG_3__5_ & ~n84806;
  assign n84828 = n83583 & n84809;
  assign n84829 = n83585 & n84793;
  assign n84830 = n83596 & n84802;
  assign n84831 = n83608 & n84800;
  assign n84832 = ~n84827 & ~n84828;
  assign n84833 = ~n84829 & n84832;
  assign n84834 = ~n84830 & n84833;
  assign n15331 = n84831 | ~n84834;
  assign n84836 = P2_P1_INSTQUEUE_REG_3__4_ & ~n84806;
  assign n84837 = n83627 & n84809;
  assign n84838 = n83629 & n84793;
  assign n84839 = n83642 & n84802;
  assign n84840 = n83654 & n84800;
  assign n84841 = ~n84836 & ~n84837;
  assign n84842 = ~n84838 & n84841;
  assign n84843 = ~n84839 & n84842;
  assign n15336 = n84840 | ~n84843;
  assign n84845 = P2_P1_INSTQUEUE_REG_3__3_ & ~n84806;
  assign n84846 = n83671 & n84809;
  assign n84847 = n83673 & n84793;
  assign n84848 = n83685 & n84802;
  assign n84849 = n83695 & n84800;
  assign n84850 = ~n84845 & ~n84846;
  assign n84851 = ~n84847 & n84850;
  assign n84852 = ~n84848 & n84851;
  assign n15341 = n84849 | ~n84852;
  assign n84854 = P2_P1_INSTQUEUE_REG_3__2_ & ~n84806;
  assign n84855 = n83713 & n84809;
  assign n84856 = n83715 & n84793;
  assign n84857 = n83729 & n84802;
  assign n84858 = n83743 & n84800;
  assign n84859 = ~n84854 & ~n84855;
  assign n84860 = ~n84856 & n84859;
  assign n84861 = ~n84857 & n84860;
  assign n15346 = n84858 | ~n84861;
  assign n84863 = P2_P1_INSTQUEUE_REG_3__1_ & ~n84806;
  assign n84864 = n83758 & n84809;
  assign n84865 = n83760 & n84793;
  assign n84866 = n83769 & n84802;
  assign n84867 = n83781 & n84800;
  assign n84868 = ~n84863 & ~n84864;
  assign n84869 = ~n84865 & n84868;
  assign n84870 = ~n84866 & n84869;
  assign n15351 = n84867 | ~n84870;
  assign n84872 = P2_P1_INSTQUEUE_REG_3__0_ & ~n84806;
  assign n84873 = n83791 & n84809;
  assign n84874 = n83793 & n84793;
  assign n84875 = n83806 & n84802;
  assign n84876 = n83820 & n84800;
  assign n84877 = ~n84872 & ~n84873;
  assign n84878 = ~n84874 & n84877;
  assign n84879 = ~n84875 & n84878;
  assign n15356 = n84876 | ~n84879;
  assign n84881 = n84184 & n84530;
  assign n84882 = P2_P1_STATE2_REG_3_ & ~n84881;
  assign n84883 = n77374 & ~n84882;
  assign n84884 = n77392 & n84796;
  assign n84885 = ~n84881 & ~n84884;
  assign n84886 = n83833 & n84799;
  assign n84887 = n77395 & n84801;
  assign n84888 = ~n84886 & ~n84887;
  assign n84889 = n77391 & ~n84888;
  assign n84890 = n84885 & ~n84889;
  assign n84891 = n84883 & ~n84890;
  assign n84892 = P2_P1_INSTQUEUE_REG_2__7_ & ~n84891;
  assign n84893 = n77427 & n84881;
  assign n84894 = ~n84719 & ~n84885;
  assign n84895 = n77701 & n84894;
  assign n84896 = n80593 & n84887;
  assign n84897 = ~n84892 & ~n84893;
  assign n84898 = ~n84895 & n84897;
  assign n84899 = ~n84896 & n84898;
  assign n84900 = ~n83519 & n84899;
  assign n84901 = ~n84886 & n84899;
  assign n15361 = ~n84900 & ~n84901;
  assign n84903 = P2_P1_INSTQUEUE_REG_2__6_ & ~n84891;
  assign n84904 = n83536 & n84894;
  assign n84905 = n83538 & n84881;
  assign n84906 = n83552 & n84887;
  assign n84907 = n83566 & n84886;
  assign n84908 = ~n84903 & ~n84904;
  assign n84909 = ~n84905 & n84908;
  assign n84910 = ~n84906 & n84909;
  assign n15366 = n84907 | ~n84910;
  assign n84912 = P2_P1_INSTQUEUE_REG_2__5_ & ~n84891;
  assign n84913 = n83583 & n84894;
  assign n84914 = n83585 & n84881;
  assign n84915 = n83596 & n84887;
  assign n84916 = n83608 & n84886;
  assign n84917 = ~n84912 & ~n84913;
  assign n84918 = ~n84914 & n84917;
  assign n84919 = ~n84915 & n84918;
  assign n15371 = n84916 | ~n84919;
  assign n84921 = P2_P1_INSTQUEUE_REG_2__4_ & ~n84891;
  assign n84922 = n83627 & n84894;
  assign n84923 = n83629 & n84881;
  assign n84924 = n83642 & n84887;
  assign n84925 = n83654 & n84886;
  assign n84926 = ~n84921 & ~n84922;
  assign n84927 = ~n84923 & n84926;
  assign n84928 = ~n84924 & n84927;
  assign n15376 = n84925 | ~n84928;
  assign n84930 = P2_P1_INSTQUEUE_REG_2__3_ & ~n84891;
  assign n84931 = n83671 & n84894;
  assign n84932 = n83673 & n84881;
  assign n84933 = n83685 & n84887;
  assign n84934 = n83695 & n84886;
  assign n84935 = ~n84930 & ~n84931;
  assign n84936 = ~n84932 & n84935;
  assign n84937 = ~n84933 & n84936;
  assign n15381 = n84934 | ~n84937;
  assign n84939 = P2_P1_INSTQUEUE_REG_2__2_ & ~n84891;
  assign n84940 = n83713 & n84894;
  assign n84941 = n83715 & n84881;
  assign n84942 = n83729 & n84887;
  assign n84943 = n83743 & n84886;
  assign n84944 = ~n84939 & ~n84940;
  assign n84945 = ~n84941 & n84944;
  assign n84946 = ~n84942 & n84945;
  assign n15386 = n84943 | ~n84946;
  assign n84948 = P2_P1_INSTQUEUE_REG_2__1_ & ~n84891;
  assign n84949 = n83758 & n84894;
  assign n84950 = n83760 & n84881;
  assign n84951 = n83769 & n84887;
  assign n84952 = n83781 & n84886;
  assign n84953 = ~n84948 & ~n84949;
  assign n84954 = ~n84950 & n84953;
  assign n84955 = ~n84951 & n84954;
  assign n15391 = n84952 | ~n84955;
  assign n84957 = P2_P1_INSTQUEUE_REG_2__0_ & ~n84891;
  assign n84958 = n83791 & n84894;
  assign n84959 = n83793 & n84881;
  assign n84960 = n83806 & n84887;
  assign n84961 = n83820 & n84886;
  assign n84962 = ~n84957 & ~n84958;
  assign n84963 = ~n84959 & n84962;
  assign n84964 = ~n84960 & n84963;
  assign n15396 = n84961 | ~n84964;
  assign n84966 = n77383 & n84792;
  assign n84967 = P2_P1_STATE2_REG_3_ & ~n84966;
  assign n84968 = n77374 & ~n84967;
  assign n84969 = n77393 & n84796;
  assign n84970 = ~n84966 & ~n84969;
  assign n84971 = n83922 & n84799;
  assign n84972 = n77396 & n84801;
  assign n84973 = ~n84971 & ~n84972;
  assign n84974 = n77391 & ~n84973;
  assign n84975 = n84970 & ~n84974;
  assign n84976 = n84968 & ~n84975;
  assign n84977 = P2_P1_INSTQUEUE_REG_1__7_ & ~n84976;
  assign n84978 = n77427 & n84966;
  assign n84979 = ~n84719 & ~n84970;
  assign n84980 = n77701 & n84979;
  assign n84981 = n80593 & n84972;
  assign n84982 = ~n84977 & ~n84978;
  assign n84983 = ~n84980 & n84982;
  assign n84984 = ~n84981 & n84983;
  assign n84985 = ~n83519 & n84984;
  assign n84986 = ~n84971 & n84984;
  assign n15401 = ~n84985 & ~n84986;
  assign n84988 = P2_P1_INSTQUEUE_REG_1__6_ & ~n84976;
  assign n84989 = n83536 & n84979;
  assign n84990 = n83538 & n84966;
  assign n84991 = n83552 & n84972;
  assign n84992 = n83566 & n84971;
  assign n84993 = ~n84988 & ~n84989;
  assign n84994 = ~n84990 & n84993;
  assign n84995 = ~n84991 & n84994;
  assign n15406 = n84992 | ~n84995;
  assign n84997 = P2_P1_INSTQUEUE_REG_1__5_ & ~n84976;
  assign n84998 = n83583 & n84979;
  assign n84999 = n83585 & n84966;
  assign n85000 = n83596 & n84972;
  assign n85001 = n83608 & n84971;
  assign n85002 = ~n84997 & ~n84998;
  assign n85003 = ~n84999 & n85002;
  assign n85004 = ~n85000 & n85003;
  assign n15411 = n85001 | ~n85004;
  assign n85006 = P2_P1_INSTQUEUE_REG_1__4_ & ~n84976;
  assign n85007 = n83627 & n84979;
  assign n85008 = n83629 & n84966;
  assign n85009 = n83642 & n84972;
  assign n85010 = n83654 & n84971;
  assign n85011 = ~n85006 & ~n85007;
  assign n85012 = ~n85008 & n85011;
  assign n85013 = ~n85009 & n85012;
  assign n15416 = n85010 | ~n85013;
  assign n85015 = P2_P1_INSTQUEUE_REG_1__3_ & ~n84976;
  assign n85016 = n83671 & n84979;
  assign n85017 = n83673 & n84966;
  assign n85018 = n83685 & n84972;
  assign n85019 = n83695 & n84971;
  assign n85020 = ~n85015 & ~n85016;
  assign n85021 = ~n85017 & n85020;
  assign n85022 = ~n85018 & n85021;
  assign n15421 = n85019 | ~n85022;
  assign n85024 = P2_P1_INSTQUEUE_REG_1__2_ & ~n84976;
  assign n85025 = n83713 & n84979;
  assign n85026 = n83715 & n84966;
  assign n85027 = n83729 & n84972;
  assign n85028 = n83743 & n84971;
  assign n85029 = ~n85024 & ~n85025;
  assign n85030 = ~n85026 & n85029;
  assign n85031 = ~n85027 & n85030;
  assign n15426 = n85028 | ~n85031;
  assign n85033 = P2_P1_INSTQUEUE_REG_1__1_ & ~n84976;
  assign n85034 = n83758 & n84979;
  assign n85035 = n83760 & n84966;
  assign n85036 = n83769 & n84972;
  assign n85037 = n83781 & n84971;
  assign n85038 = ~n85033 & ~n85034;
  assign n85039 = ~n85035 & n85038;
  assign n85040 = ~n85036 & n85039;
  assign n15431 = n85037 | ~n85040;
  assign n85042 = P2_P1_INSTQUEUE_REG_1__0_ & ~n84976;
  assign n85043 = n83791 & n84979;
  assign n85044 = n83793 & n84966;
  assign n85045 = n83806 & n84972;
  assign n85046 = n83820 & n84971;
  assign n85047 = ~n85042 & ~n85043;
  assign n85048 = ~n85044 & n85047;
  assign n85049 = ~n85045 & n85048;
  assign n15436 = n85046 | ~n85049;
  assign n85051 = n84184 & n84706;
  assign n85052 = P2_P1_STATE2_REG_3_ & ~n85051;
  assign n85053 = n77374 & ~n85052;
  assign n85054 = n84009 & n84799;
  assign n85055 = n84011 & n84801;
  assign n85056 = ~n85054 & ~n85055;
  assign n85057 = n77391 & ~n85056;
  assign n85058 = n77385 & n84796;
  assign n85059 = ~n85057 & ~n85058;
  assign n85060 = n85053 & ~n85059;
  assign n85061 = P2_P1_INSTQUEUE_REG_0__7_ & ~n85060;
  assign n85062 = n77427 & n85051;
  assign n85063 = ~n84719 & n85058;
  assign n85064 = n77701 & n85063;
  assign n85065 = n80593 & n85055;
  assign n85066 = ~n85061 & ~n85062;
  assign n85067 = ~n85064 & n85066;
  assign n85068 = ~n85065 & n85067;
  assign n85069 = ~n83519 & n85068;
  assign n85070 = ~n85054 & n85068;
  assign n15441 = ~n85069 & ~n85070;
  assign n85072 = P2_P1_INSTQUEUE_REG_0__6_ & ~n85060;
  assign n85073 = n83536 & n85063;
  assign n85074 = n83538 & n85051;
  assign n85075 = n83552 & n85055;
  assign n85076 = n83566 & n85054;
  assign n85077 = ~n85072 & ~n85073;
  assign n85078 = ~n85074 & n85077;
  assign n85079 = ~n85075 & n85078;
  assign n15446 = n85076 | ~n85079;
  assign n85081 = P2_P1_INSTQUEUE_REG_0__5_ & ~n85060;
  assign n85082 = n83583 & n85063;
  assign n85083 = n83585 & n85051;
  assign n85084 = n83596 & n85055;
  assign n85085 = n83608 & n85054;
  assign n85086 = ~n85081 & ~n85082;
  assign n85087 = ~n85083 & n85086;
  assign n85088 = ~n85084 & n85087;
  assign n15451 = n85085 | ~n85088;
  assign n85090 = P2_P1_INSTQUEUE_REG_0__4_ & ~n85060;
  assign n85091 = n83627 & n85063;
  assign n85092 = n83629 & n85051;
  assign n85093 = n83642 & n85055;
  assign n85094 = n83654 & n85054;
  assign n85095 = ~n85090 & ~n85091;
  assign n85096 = ~n85092 & n85095;
  assign n85097 = ~n85093 & n85096;
  assign n15456 = n85094 | ~n85097;
  assign n85099 = P2_P1_INSTQUEUE_REG_0__3_ & ~n85060;
  assign n85100 = n83671 & n85063;
  assign n85101 = n83673 & n85051;
  assign n85102 = n83685 & n85055;
  assign n85103 = n83695 & n85054;
  assign n85104 = ~n85099 & ~n85100;
  assign n85105 = ~n85101 & n85104;
  assign n85106 = ~n85102 & n85105;
  assign n15461 = n85103 | ~n85106;
  assign n85108 = P2_P1_INSTQUEUE_REG_0__2_ & ~n85060;
  assign n85109 = n83713 & n85063;
  assign n85110 = n83715 & n85051;
  assign n85111 = n83729 & n85055;
  assign n85112 = n83743 & n85054;
  assign n85113 = ~n85108 & ~n85109;
  assign n85114 = ~n85110 & n85113;
  assign n85115 = ~n85111 & n85114;
  assign n15466 = n85112 | ~n85115;
  assign n85117 = P2_P1_INSTQUEUE_REG_0__1_ & ~n85060;
  assign n85118 = n83758 & n85063;
  assign n85119 = n83760 & n85051;
  assign n85120 = n83769 & n85055;
  assign n85121 = n83781 & n85054;
  assign n85122 = ~n85117 & ~n85118;
  assign n85123 = ~n85119 & n85122;
  assign n85124 = ~n85120 & n85123;
  assign n15471 = n85121 | ~n85124;
  assign n85126 = P2_P1_INSTQUEUE_REG_0__0_ & ~n85060;
  assign n85127 = n83791 & n85063;
  assign n85128 = n83793 & n85051;
  assign n85129 = n83806 & n85055;
  assign n85130 = n83820 & n85054;
  assign n85131 = ~n85126 & ~n85127;
  assign n85132 = ~n85128 & n85131;
  assign n85133 = ~n85129 & n85132;
  assign n15476 = n85130 | ~n85133;
  assign n85135 = P2_P1_STATE2_REG_3_ & ~P2_P1_STATE2_REG_0_;
  assign n85136 = P2_P1_STATE2_REG_0_ & P2_P1_FLUSH_REG;
  assign n85137 = n76669 & n85136;
  assign n85138 = ~n85135 & ~n85137;
  assign n85139 = ~n77201 & n77311;
  assign n85140 = n85138 & ~n85139;
  assign n85141 = P2_P1_INSTQUEUERD_ADDR_REG_4_ & n85140;
  assign n85142 = ~n77244 & n77317;
  assign n85143 = n77036 & n85142;
  assign n85144 = ~n85140 & n85143;
  assign n15481 = n85141 | n85144;
  assign n85146 = ~n77235 & n77317;
  assign n85147 = ~n76708 & ~n77208;
  assign n85148 = n77326 & ~n85147;
  assign n85149 = ~n85146 & ~n85148;
  assign n85150 = ~n85140 & ~n85149;
  assign n85151 = P2_P1_INSTQUEUERD_ADDR_REG_3_ & n85140;
  assign n15486 = n85150 | n85151;
  assign n85153 = ~n77159 & n77326;
  assign n85154 = P2_P1_STATE2_REG_1_ & ~n77333;
  assign n85155 = ~n77342 & n85154;
  assign n85156 = ~n85153 & ~n85155;
  assign n85157 = ~n77175 & n77317;
  assign n85158 = n85156 & ~n85157;
  assign n85159 = ~n85140 & ~n85158;
  assign n85160 = P2_P1_INSTQUEUERD_ADDR_REG_2_ & n85140;
  assign n15491 = n85159 | n85160;
  assign n85162 = n77271 & n77326;
  assign n85163 = n77342 & n85154;
  assign n85164 = ~n85162 & ~n85163;
  assign n85165 = ~n77276 & n77317;
  assign n85166 = n85164 & ~n85165;
  assign n85167 = ~n85140 & ~n85166;
  assign n85168 = P2_P1_INSTQUEUERD_ADDR_REG_1_ & n85140;
  assign n15496 = n85167 | n85168;
  assign n85170 = P2_P1_STATE2_REG_1_ & n77333;
  assign n85171 = ~P2_P1_INSTQUEUERD_ADDR_REG_0_ & n77326;
  assign n85172 = ~n85170 & ~n85171;
  assign n85173 = ~n77262 & n77317;
  assign n85174 = n85172 & ~n85173;
  assign n85175 = ~n85140 & ~n85174;
  assign n85176 = P2_P1_INSTQUEUERD_ADDR_REG_0_ & n85140;
  assign n15501 = n85175 | n85176;
  assign n85178 = P2_P1_STATE2_REG_0_ & n76669;
  assign n85179 = ~n77356 & n85178;
  assign n85180 = ~n77374 & ~n85137;
  assign n85181 = ~n85179 & n85180;
  assign n15506 = P2_P1_INSTQUEUEWR_ADDR_REG_4_ & n85181;
  assign n85183 = P2_P1_STATE2_REG_3_ & ~n77368;
  assign n85184 = ~n85181 & ~n85183;
  assign n85185 = P2_P1_INSTQUEUEWR_ADDR_REG_3_ & ~n85184;
  assign n85186 = ~n77317 & ~n77390;
  assign n85187 = ~n77410 & ~n85186;
  assign n85188 = P2_P1_STATE2_REG_3_ & n77379;
  assign n85189 = ~n85187 & ~n85188;
  assign n85190 = n77398 & ~n77405;
  assign n85191 = ~n77416 & ~n85190;
  assign n85192 = ~n84449 & ~n85191;
  assign n85193 = n77429 & ~n85192;
  assign n85194 = n85189 & ~n85193;
  assign n85195 = ~n85181 & ~n85194;
  assign n15511 = n85185 | n85195;
  assign n85197 = ~n77401 & ~n85186;
  assign n85198 = P2_P1_STATE2_REG_3_ & ~P2_P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n85199 = n77367 & n85198;
  assign n85200 = ~n85197 & ~n85199;
  assign n85201 = ~n77398 & ~n77405;
  assign n85202 = n77398 & n77405;
  assign n85203 = ~n85201 & ~n85202;
  assign n85204 = n77429 & ~n85203;
  assign n85205 = n85200 & ~n85204;
  assign n85206 = ~n85181 & ~n85205;
  assign n85207 = P2_P1_STATE2_REG_3_ & ~n77367;
  assign n85208 = ~n85181 & ~n85207;
  assign n85209 = P2_P1_INSTQUEUEWR_ADDR_REG_2_ & ~n85208;
  assign n15516 = n85206 | n85209;
  assign n85211 = ~n77394 & ~n85186;
  assign n85212 = P2_P1_STATE2_REG_3_ & ~P2_P1_INSTQUEUEWR_ADDR_REG_1_;
  assign n85213 = ~n77397 & n77429;
  assign n85214 = ~n85212 & ~n85213;
  assign n85215 = P2_P1_INSTQUEUEWR_ADDR_REG_0_ & ~n85214;
  assign n85216 = n77429 & n83922;
  assign n85217 = ~n85211 & ~n85215;
  assign n85218 = ~n85216 & n85217;
  assign n85219 = ~n85181 & ~n85218;
  assign n85220 = P2_P1_STATE2_REG_3_ & ~P2_P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n85221 = ~n85181 & ~n85220;
  assign n85222 = P2_P1_INSTQUEUEWR_ADDR_REG_1_ & ~n85221;
  assign n15521 = n85219 | n85222;
  assign n85224 = ~n77317 & ~n77389;
  assign n85225 = ~n85181 & n85224;
  assign n85226 = P2_P1_INSTQUEUEWR_ADDR_REG_0_ & ~n85225;
  assign n85227 = ~n77357 & ~n85220;
  assign n85228 = ~n85181 & ~n85227;
  assign n15526 = n85226 | n85228;
  assign n85230 = ~P2_P1_STATE2_REG_1_ & n77389;
  assign n85231 = ~P2_P1_STATE2_REG_0_ & n85230;
  assign n85232 = n76965 & n77009;
  assign n85233 = ~n76797 & ~n76956;
  assign n85234 = n77054 & n85233;
  assign n85235 = n76963 & n77009;
  assign n85236 = ~n77193 & ~n85234;
  assign n85237 = ~n85235 & n85236;
  assign n85238 = n77014 & n77062;
  assign n85239 = n76766 & n76961;
  assign n85240 = n77009 & n85239;
  assign n85241 = ~n85238 & ~n85240;
  assign n85242 = n76925 & ~n85241;
  assign n85243 = ~n76765 & n77068;
  assign n85244 = ~n76584 & n76734;
  assign n85245 = n77009 & n85244;
  assign n85246 = ~n85243 & ~n85245;
  assign n85247 = ~n76925 & ~n85246;
  assign n85248 = n76956 & n77054;
  assign n85249 = ~n85242 & ~n85247;
  assign n85250 = ~n85248 & n85249;
  assign n85251 = n76890 & ~n85250;
  assign n85252 = n77185 & ~n85232;
  assign n85253 = n85237 & n85252;
  assign n85254 = ~n85251 & n85253;
  assign n85255 = n77311 & ~n85254;
  assign n85256 = ~n85231 & ~n85255;
  assign n85257 = P2_P1_STATE2_REG_2_ & ~n85256;
  assign n85258 = ~P2_P1_INSTADDRPOINTER_REG_0_ & n77255;
  assign n85259 = ~P2_P1_INSTADDRPOINTER_REG_0_ & n77098;
  assign n85260 = ~n85258 & ~n85259;
  assign n85261 = ~P2_P1_INSTADDRPOINTER_REG_0_ & ~n77145;
  assign n85262 = P2_P1_INSTADDRPOINTER_REG_0_ & n77216;
  assign n85263 = P2_P1_INSTADDRPOINTER_REG_0_ & n77217;
  assign n85264 = n76957 & n77088;
  assign n85265 = n77094 & n85264;
  assign n85266 = ~P2_P1_INSTADDRPOINTER_REG_0_ & n85265;
  assign n85267 = n77034 & n77088;
  assign n85268 = n77094 & n85267;
  assign n85269 = ~P2_P1_INSTADDRPOINTER_REG_0_ & n85268;
  assign n85270 = ~n85266 & ~n85269;
  assign n85271 = P2_P1_INSTADDRPOINTER_REG_0_ & n77032;
  assign n85272 = n85270 & ~n85271;
  assign n85273 = n77159 & n85147;
  assign n85274 = P2_P1_INSTQUEUERD_ADDR_REG_0_ & ~n77271;
  assign n85275 = n85273 & n85274;
  assign n85276 = P2_P1_INSTQUEUE_REG_0__0_ & n85275;
  assign n85277 = ~P2_P1_INSTQUEUERD_ADDR_REG_0_ & ~n77271;
  assign n85278 = n85273 & n85277;
  assign n85279 = P2_P1_INSTQUEUE_REG_1__0_ & n85278;
  assign n85280 = P2_P1_INSTQUEUERD_ADDR_REG_0_ & n77271;
  assign n85281 = n85273 & n85280;
  assign n85282 = P2_P1_INSTQUEUE_REG_2__0_ & n85281;
  assign n85283 = ~P2_P1_INSTQUEUERD_ADDR_REG_0_ & n77271;
  assign n85284 = n85273 & n85283;
  assign n85285 = P2_P1_INSTQUEUE_REG_3__0_ & n85284;
  assign n85286 = ~n85276 & ~n85279;
  assign n85287 = ~n85282 & n85286;
  assign n85288 = ~n85285 & n85287;
  assign n85289 = ~n77159 & n85147;
  assign n85290 = n85274 & n85289;
  assign n85291 = P2_P1_INSTQUEUE_REG_4__0_ & n85290;
  assign n85292 = n85277 & n85289;
  assign n85293 = P2_P1_INSTQUEUE_REG_5__0_ & n85292;
  assign n85294 = n85280 & n85289;
  assign n85295 = P2_P1_INSTQUEUE_REG_6__0_ & n85294;
  assign n85296 = n85283 & n85289;
  assign n85297 = P2_P1_INSTQUEUE_REG_7__0_ & n85296;
  assign n85298 = ~n85291 & ~n85293;
  assign n85299 = ~n85295 & n85298;
  assign n85300 = ~n85297 & n85299;
  assign n85301 = n77159 & ~n85147;
  assign n85302 = n85274 & n85301;
  assign n85303 = P2_P1_INSTQUEUE_REG_8__0_ & n85302;
  assign n85304 = n85277 & n85301;
  assign n85305 = P2_P1_INSTQUEUE_REG_9__0_ & n85304;
  assign n85306 = n85280 & n85301;
  assign n85307 = P2_P1_INSTQUEUE_REG_10__0_ & n85306;
  assign n85308 = n85283 & n85301;
  assign n85309 = P2_P1_INSTQUEUE_REG_11__0_ & n85308;
  assign n85310 = ~n85303 & ~n85305;
  assign n85311 = ~n85307 & n85310;
  assign n85312 = ~n85309 & n85311;
  assign n85313 = ~n77159 & ~n85147;
  assign n85314 = n85274 & n85313;
  assign n85315 = P2_P1_INSTQUEUE_REG_12__0_ & n85314;
  assign n85316 = n85277 & n85313;
  assign n85317 = P2_P1_INSTQUEUE_REG_13__0_ & n85316;
  assign n85318 = n85280 & n85313;
  assign n85319 = P2_P1_INSTQUEUE_REG_14__0_ & n85318;
  assign n85320 = n85283 & n85313;
  assign n85321 = P2_P1_INSTQUEUE_REG_15__0_ & n85320;
  assign n85322 = ~n85315 & ~n85317;
  assign n85323 = ~n85319 & n85322;
  assign n85324 = ~n85321 & n85323;
  assign n85325 = n85288 & n85300;
  assign n85326 = n85312 & n85325;
  assign n85327 = n85324 & n85326;
  assign n85328 = P2_P1_INSTADDRPOINTER_REG_0_ & n85327;
  assign n85329 = ~P2_P1_INSTADDRPOINTER_REG_0_ & ~n85327;
  assign n85330 = ~n85328 & ~n85329;
  assign n85331 = P2_P1_INSTQUEUE_REG_0__7_ & n85275;
  assign n85332 = P2_P1_INSTQUEUE_REG_1__7_ & n85278;
  assign n85333 = P2_P1_INSTQUEUE_REG_2__7_ & n85281;
  assign n85334 = P2_P1_INSTQUEUE_REG_3__7_ & n85284;
  assign n85335 = ~n85331 & ~n85332;
  assign n85336 = ~n85333 & n85335;
  assign n85337 = ~n85334 & n85336;
  assign n85338 = P2_P1_INSTQUEUE_REG_4__7_ & n85290;
  assign n85339 = P2_P1_INSTQUEUE_REG_5__7_ & n85292;
  assign n85340 = P2_P1_INSTQUEUE_REG_6__7_ & n85294;
  assign n85341 = P2_P1_INSTQUEUE_REG_7__7_ & n85296;
  assign n85342 = ~n85338 & ~n85339;
  assign n85343 = ~n85340 & n85342;
  assign n85344 = ~n85341 & n85343;
  assign n85345 = P2_P1_INSTQUEUE_REG_8__7_ & n85302;
  assign n85346 = P2_P1_INSTQUEUE_REG_9__7_ & n85304;
  assign n85347 = P2_P1_INSTQUEUE_REG_10__7_ & n85306;
  assign n85348 = P2_P1_INSTQUEUE_REG_11__7_ & n85308;
  assign n85349 = ~n85345 & ~n85346;
  assign n85350 = ~n85347 & n85349;
  assign n85351 = ~n85348 & n85350;
  assign n85352 = P2_P1_INSTQUEUE_REG_12__7_ & n85314;
  assign n85353 = P2_P1_INSTQUEUE_REG_13__7_ & n85316;
  assign n85354 = P2_P1_INSTQUEUE_REG_14__7_ & n85318;
  assign n85355 = P2_P1_INSTQUEUE_REG_15__7_ & n85320;
  assign n85356 = ~n85352 & ~n85353;
  assign n85357 = ~n85354 & n85356;
  assign n85358 = ~n85355 & n85357;
  assign n85359 = n85337 & n85344;
  assign n85360 = n85351 & n85359;
  assign n85361 = n85358 & n85360;
  assign n85362 = n77064 & ~n85361;
  assign n85363 = ~n85330 & n85362;
  assign n85364 = n77064 & n85361;
  assign n85365 = ~n85330 & n85364;
  assign n85366 = ~n85262 & ~n85263;
  assign n85367 = n85272 & n85366;
  assign n85368 = ~n85363 & n85367;
  assign n85369 = ~n85365 & n85368;
  assign n85370 = n77030 & n77058;
  assign n85371 = ~P2_P1_INSTADDRPOINTER_REG_0_ & n85370;
  assign n85372 = ~P2_P1_INSTADDRPOINTER_REG_0_ & n77102;
  assign n85373 = n76859 & n77045;
  assign n85374 = n77091 & n85373;
  assign n85375 = ~P2_P1_INSTADDRPOINTER_REG_0_ & n85374;
  assign n85376 = ~P2_P1_INSTADDRPOINTER_REG_0_ & n85327;
  assign n85377 = P2_P1_INSTADDRPOINTER_REG_0_ & ~n85327;
  assign n85378 = ~n85376 & ~n85377;
  assign n85379 = n77059 & ~n85378;
  assign n85380 = n76734 & n77088;
  assign n85381 = n77091 & n85380;
  assign n85382 = ~P2_P1_INSTADDRPOINTER_REG_0_ & n85381;
  assign n85383 = ~n85371 & ~n85372;
  assign n85384 = ~n85375 & n85383;
  assign n85385 = ~n85379 & n85384;
  assign n85386 = ~n85382 & n85385;
  assign n85387 = P2_P1_INSTADDRPOINTER_REG_0_ & n76958;
  assign n85388 = P2_P1_INSTADDRPOINTER_REG_0_ & n77036;
  assign n85389 = P2_P1_INSTADDRPOINTER_REG_0_ & n77040;
  assign n85390 = ~P2_P1_INSTADDRPOINTER_REG_0_ & n77056;
  assign n85391 = ~P2_P1_INSTADDRPOINTER_REG_0_ & n77048;
  assign n85392 = ~n85387 & ~n85388;
  assign n85393 = ~n85389 & n85392;
  assign n85394 = ~n85390 & n85393;
  assign n85395 = ~n85391 & n85394;
  assign n85396 = n85386 & n85395;
  assign n85397 = n85260 & ~n85261;
  assign n85398 = n85369 & n85397;
  assign n85399 = n85396 & n85398;
  assign n85400 = n85257 & ~n85399;
  assign n85401 = ~P2_P1_STATE2_REG_2_ & ~n85256;
  assign n85402 = P2_P1_REIP_REG_0_ & n85401;
  assign n85403 = P2_P1_INSTADDRPOINTER_REG_0_ & n85256;
  assign n85404 = ~n85400 & ~n85402;
  assign n15531 = n85403 | ~n85404;
  assign n85406 = P2_P1_INSTADDRPOINTER_REG_1_ & n85256;
  assign n85407 = P2_P1_REIP_REG_1_ & n85401;
  assign n85408 = ~n77145 & ~n77339;
  assign n85409 = n77255 & ~n77339;
  assign n85410 = n77098 & ~n77339;
  assign n85411 = ~n85409 & ~n85410;
  assign n85412 = ~P2_P1_INSTADDRPOINTER_REG_1_ & n85377;
  assign n85413 = P2_P1_INSTADDRPOINTER_REG_1_ & ~n85377;
  assign n85414 = ~n85412 & ~n85413;
  assign n85415 = P2_P1_INSTQUEUE_REG_0__1_ & n85275;
  assign n85416 = P2_P1_INSTQUEUE_REG_1__1_ & n85278;
  assign n85417 = P2_P1_INSTQUEUE_REG_2__1_ & n85281;
  assign n85418 = P2_P1_INSTQUEUE_REG_3__1_ & n85284;
  assign n85419 = ~n85415 & ~n85416;
  assign n85420 = ~n85417 & n85419;
  assign n85421 = ~n85418 & n85420;
  assign n85422 = P2_P1_INSTQUEUE_REG_4__1_ & n85290;
  assign n85423 = P2_P1_INSTQUEUE_REG_5__1_ & n85292;
  assign n85424 = P2_P1_INSTQUEUE_REG_6__1_ & n85294;
  assign n85425 = P2_P1_INSTQUEUE_REG_7__1_ & n85296;
  assign n85426 = ~n85422 & ~n85423;
  assign n85427 = ~n85424 & n85426;
  assign n85428 = ~n85425 & n85427;
  assign n85429 = P2_P1_INSTQUEUE_REG_8__1_ & n85302;
  assign n85430 = P2_P1_INSTQUEUE_REG_9__1_ & n85304;
  assign n85431 = P2_P1_INSTQUEUE_REG_10__1_ & n85306;
  assign n85432 = P2_P1_INSTQUEUE_REG_11__1_ & n85308;
  assign n85433 = ~n85429 & ~n85430;
  assign n85434 = ~n85431 & n85433;
  assign n85435 = ~n85432 & n85434;
  assign n85436 = P2_P1_INSTQUEUE_REG_12__1_ & n85314;
  assign n85437 = P2_P1_INSTQUEUE_REG_13__1_ & n85316;
  assign n85438 = P2_P1_INSTQUEUE_REG_14__1_ & n85318;
  assign n85439 = P2_P1_INSTQUEUE_REG_15__1_ & n85320;
  assign n85440 = ~n85436 & ~n85437;
  assign n85441 = ~n85438 & n85440;
  assign n85442 = ~n85439 & n85441;
  assign n85443 = n85421 & n85428;
  assign n85444 = n85435 & n85443;
  assign n85445 = n85442 & n85444;
  assign n85446 = ~n85414 & ~n85445;
  assign n85447 = ~P2_P1_INSTADDRPOINTER_REG_1_ & ~n85377;
  assign n85448 = n85445 & n85447;
  assign n85449 = n85377 & n85445;
  assign n85450 = P2_P1_INSTADDRPOINTER_REG_1_ & n85449;
  assign n85451 = ~n85446 & ~n85448;
  assign n85452 = ~n85450 & n85451;
  assign n85453 = n85364 & ~n85452;
  assign n85454 = ~n77339 & n85381;
  assign n85455 = ~n77339 & n85374;
  assign n85456 = ~n77339 & n85370;
  assign n85457 = n77102 & ~n77339;
  assign n85458 = ~n85454 & ~n85455;
  assign n85459 = ~n85456 & n85458;
  assign n85460 = ~n85457 & n85459;
  assign n85461 = ~P2_P1_INSTADDRPOINTER_REG_1_ & n76958;
  assign n85462 = ~P2_P1_INSTADDRPOINTER_REG_1_ & n77036;
  assign n85463 = ~P2_P1_INSTADDRPOINTER_REG_1_ & n77040;
  assign n85464 = n77056 & ~n77339;
  assign n85465 = n77048 & ~n77339;
  assign n85466 = ~n85461 & ~n85462;
  assign n85467 = ~n85463 & n85466;
  assign n85468 = ~n85464 & n85467;
  assign n85469 = ~n85465 & n85468;
  assign n85470 = ~P2_P1_INSTADDRPOINTER_REG_1_ & n85328;
  assign n85471 = P2_P1_INSTADDRPOINTER_REG_1_ & ~n85328;
  assign n85472 = ~n85470 & ~n85471;
  assign n85473 = ~n85327 & n85445;
  assign n85474 = n85327 & ~n85445;
  assign n85475 = ~n85473 & ~n85474;
  assign n85476 = ~n85472 & n85475;
  assign n85477 = ~P2_P1_INSTADDRPOINTER_REG_1_ & ~n85328;
  assign n85478 = ~n85475 & n85477;
  assign n85479 = n85328 & ~n85475;
  assign n85480 = P2_P1_INSTADDRPOINTER_REG_1_ & n85479;
  assign n85481 = ~n85476 & ~n85478;
  assign n85482 = ~n85480 & n85481;
  assign n85483 = n77059 & ~n85482;
  assign n85484 = n85460 & n85469;
  assign n85485 = ~n85483 & n85484;
  assign n85486 = ~P2_P1_INSTADDRPOINTER_REG_1_ & n77216;
  assign n85487 = ~P2_P1_INSTADDRPOINTER_REG_1_ & n77217;
  assign n85488 = ~n77339 & n85265;
  assign n85489 = ~n77339 & n85268;
  assign n85490 = ~n85488 & ~n85489;
  assign n85491 = ~P2_P1_INSTADDRPOINTER_REG_1_ & n77032;
  assign n85492 = n85490 & ~n85491;
  assign n85493 = n85377 & ~n85445;
  assign n85494 = ~n85377 & n85445;
  assign n85495 = ~n85493 & ~n85494;
  assign n85496 = ~P2_P1_INSTADDRPOINTER_REG_1_ & ~n85495;
  assign n85497 = ~n85377 & ~n85445;
  assign n85498 = P2_P1_INSTADDRPOINTER_REG_1_ & n85497;
  assign n85499 = P2_P1_INSTADDRPOINTER_REG_1_ & n85377;
  assign n85500 = n85445 & n85499;
  assign n85501 = ~n85496 & ~n85498;
  assign n85502 = ~n85500 & n85501;
  assign n85503 = n85362 & ~n85502;
  assign n85504 = ~n85486 & ~n85487;
  assign n85505 = n85492 & n85504;
  assign n85506 = ~n85503 & n85505;
  assign n85507 = ~n85408 & n85411;
  assign n85508 = ~n85453 & n85507;
  assign n85509 = n85485 & n85508;
  assign n85510 = n85506 & n85509;
  assign n85511 = n85257 & ~n85510;
  assign n85512 = ~n85406 & ~n85407;
  assign n15536 = n85511 | ~n85512;
  assign n85514 = P2_P1_INSTADDRPOINTER_REG_2_ & n85256;
  assign n85515 = P2_P1_REIP_REG_2_ & n85401;
  assign n85516 = P2_P1_INSTADDRPOINTER_REG_0_ & P2_P1_INSTADDRPOINTER_REG_1_;
  assign n85517 = ~P2_P1_INSTADDRPOINTER_REG_2_ & n85516;
  assign n85518 = P2_P1_INSTADDRPOINTER_REG_2_ & ~n85516;
  assign n85519 = ~n85517 & ~n85518;
  assign n85520 = ~n77145 & ~n85519;
  assign n85521 = P2_P1_INSTADDRPOINTER_REG_1_ & ~P2_P1_INSTADDRPOINTER_REG_2_;
  assign n85522 = ~P2_P1_INSTADDRPOINTER_REG_1_ & P2_P1_INSTADDRPOINTER_REG_2_;
  assign n85523 = ~n85521 & ~n85522;
  assign n85524 = n77216 & ~n85523;
  assign n85525 = n77217 & ~n85523;
  assign n85526 = n85265 & ~n85519;
  assign n85527 = n85268 & ~n85519;
  assign n85528 = ~n85526 & ~n85527;
  assign n85529 = n77032 & ~n85523;
  assign n85530 = n85528 & ~n85529;
  assign n85531 = ~n85524 & ~n85525;
  assign n85532 = n85530 & n85531;
  assign n85533 = P2_P1_INSTADDRPOINTER_REG_1_ & ~n85497;
  assign n85534 = ~n85449 & ~n85533;
  assign n85535 = P2_P1_INSTQUEUE_REG_0__2_ & n85275;
  assign n85536 = P2_P1_INSTQUEUE_REG_1__2_ & n85278;
  assign n85537 = P2_P1_INSTQUEUE_REG_2__2_ & n85281;
  assign n85538 = P2_P1_INSTQUEUE_REG_3__2_ & n85284;
  assign n85539 = ~n85535 & ~n85536;
  assign n85540 = ~n85537 & n85539;
  assign n85541 = ~n85538 & n85540;
  assign n85542 = P2_P1_INSTQUEUE_REG_4__2_ & n85290;
  assign n85543 = P2_P1_INSTQUEUE_REG_5__2_ & n85292;
  assign n85544 = P2_P1_INSTQUEUE_REG_6__2_ & n85294;
  assign n85545 = P2_P1_INSTQUEUE_REG_7__2_ & n85296;
  assign n85546 = ~n85542 & ~n85543;
  assign n85547 = ~n85544 & n85546;
  assign n85548 = ~n85545 & n85547;
  assign n85549 = P2_P1_INSTQUEUE_REG_8__2_ & n85302;
  assign n85550 = P2_P1_INSTQUEUE_REG_9__2_ & n85304;
  assign n85551 = P2_P1_INSTQUEUE_REG_10__2_ & n85306;
  assign n85552 = P2_P1_INSTQUEUE_REG_11__2_ & n85308;
  assign n85553 = ~n85549 & ~n85550;
  assign n85554 = ~n85551 & n85553;
  assign n85555 = ~n85552 & n85554;
  assign n85556 = P2_P1_INSTQUEUE_REG_12__2_ & n85314;
  assign n85557 = P2_P1_INSTQUEUE_REG_13__2_ & n85316;
  assign n85558 = P2_P1_INSTQUEUE_REG_14__2_ & n85318;
  assign n85559 = P2_P1_INSTQUEUE_REG_15__2_ & n85320;
  assign n85560 = ~n85556 & ~n85557;
  assign n85561 = ~n85558 & n85560;
  assign n85562 = ~n85559 & n85561;
  assign n85563 = n85541 & n85548;
  assign n85564 = n85555 & n85563;
  assign n85565 = n85562 & n85564;
  assign n85566 = ~n85445 & n85565;
  assign n85567 = n85445 & ~n85565;
  assign n85568 = ~n85566 & ~n85567;
  assign n85569 = ~P2_P1_INSTADDRPOINTER_REG_2_ & ~n85568;
  assign n85570 = P2_P1_INSTADDRPOINTER_REG_2_ & n85568;
  assign n85571 = ~n85569 & ~n85570;
  assign n85572 = n85534 & ~n85571;
  assign n85573 = ~n85534 & n85571;
  assign n85574 = ~n85572 & ~n85573;
  assign n85575 = n85364 & ~n85574;
  assign n85576 = n77255 & ~n85519;
  assign n85577 = n77098 & ~n85519;
  assign n85578 = ~n85576 & ~n85577;
  assign n85579 = P2_P1_INSTADDRPOINTER_REG_1_ & n85445;
  assign n85580 = ~n85449 & ~n85499;
  assign n85581 = ~n85579 & n85580;
  assign n85582 = ~n85571 & n85581;
  assign n85583 = ~P2_P1_INSTADDRPOINTER_REG_2_ & n85568;
  assign n85584 = P2_P1_INSTADDRPOINTER_REG_2_ & ~n85568;
  assign n85585 = ~n85583 & ~n85584;
  assign n85586 = ~n85581 & ~n85585;
  assign n85587 = ~n85582 & ~n85586;
  assign n85588 = n85362 & ~n85587;
  assign n85589 = n85578 & ~n85588;
  assign n85590 = n85381 & ~n85519;
  assign n85591 = n85374 & ~n85519;
  assign n85592 = n85370 & ~n85519;
  assign n85593 = n77102 & ~n85519;
  assign n85594 = ~n85590 & ~n85591;
  assign n85595 = ~n85592 & n85594;
  assign n85596 = ~n85593 & n85595;
  assign n85597 = n76958 & ~n85523;
  assign n85598 = n77036 & ~n85523;
  assign n85599 = n77040 & ~n85523;
  assign n85600 = ~P2_P1_INSTADDRPOINTER_REG_2_ & ~n85516;
  assign n85601 = P2_P1_INSTADDRPOINTER_REG_2_ & n85516;
  assign n85602 = ~n85600 & ~n85601;
  assign n85603 = n77056 & ~n85602;
  assign n85604 = n77048 & ~n85602;
  assign n85605 = ~n85597 & ~n85598;
  assign n85606 = ~n85599 & n85605;
  assign n85607 = ~n85603 & n85606;
  assign n85608 = ~n85604 & n85607;
  assign n85609 = ~n85327 & ~n85445;
  assign n85610 = n85565 & ~n85609;
  assign n85611 = ~n85565 & n85609;
  assign n85612 = ~n85610 & ~n85611;
  assign n85613 = ~P2_P1_INSTADDRPOINTER_REG_2_ & ~n85612;
  assign n85614 = P2_P1_INSTADDRPOINTER_REG_2_ & n85612;
  assign n85615 = ~n85613 & ~n85614;
  assign n85616 = ~n85328 & n85475;
  assign n85617 = P2_P1_INSTADDRPOINTER_REG_1_ & ~n85616;
  assign n85618 = ~n85479 & ~n85617;
  assign n85619 = ~n85615 & n85618;
  assign n85620 = ~P2_P1_INSTADDRPOINTER_REG_2_ & n85612;
  assign n85621 = P2_P1_INSTADDRPOINTER_REG_2_ & ~n85612;
  assign n85622 = ~n85620 & ~n85621;
  assign n85623 = ~n85618 & ~n85622;
  assign n85624 = ~n85619 & ~n85623;
  assign n85625 = n77059 & ~n85624;
  assign n85626 = n85596 & n85608;
  assign n85627 = ~n85625 & n85626;
  assign n85628 = ~n85520 & n85532;
  assign n85629 = ~n85575 & n85628;
  assign n85630 = n85589 & n85629;
  assign n85631 = n85627 & n85630;
  assign n85632 = n85257 & ~n85631;
  assign n85633 = ~n85514 & ~n85515;
  assign n15541 = n85632 | ~n85633;
  assign n85635 = P2_P1_INSTADDRPOINTER_REG_3_ & n85256;
  assign n85636 = P2_P1_REIP_REG_3_ & n85401;
  assign n85637 = ~P2_P1_INSTADDRPOINTER_REG_3_ & n85601;
  assign n85638 = P2_P1_INSTADDRPOINTER_REG_3_ & ~n85601;
  assign n85639 = ~n85637 & ~n85638;
  assign n85640 = n77255 & ~n85639;
  assign n85641 = n77098 & ~n85639;
  assign n85642 = ~n85640 & ~n85641;
  assign n85643 = ~n77145 & ~n85639;
  assign n85644 = P2_P1_INSTADDRPOINTER_REG_1_ & P2_P1_INSTADDRPOINTER_REG_2_;
  assign n85645 = ~P2_P1_INSTADDRPOINTER_REG_3_ & n85644;
  assign n85646 = P2_P1_INSTADDRPOINTER_REG_3_ & ~n85644;
  assign n85647 = ~n85645 & ~n85646;
  assign n85648 = n77216 & ~n85647;
  assign n85649 = n77217 & ~n85647;
  assign n85650 = n85265 & ~n85639;
  assign n85651 = n85268 & ~n85639;
  assign n85652 = ~n85650 & ~n85651;
  assign n85653 = n77032 & ~n85647;
  assign n85654 = n85652 & ~n85653;
  assign n85655 = ~n85648 & ~n85649;
  assign n85656 = n85654 & n85655;
  assign n85657 = ~n85581 & ~n85583;
  assign n85658 = ~n85584 & ~n85657;
  assign n85659 = P2_P1_INSTQUEUE_REG_0__3_ & n85275;
  assign n85660 = P2_P1_INSTQUEUE_REG_1__3_ & n85278;
  assign n85661 = P2_P1_INSTQUEUE_REG_2__3_ & n85281;
  assign n85662 = P2_P1_INSTQUEUE_REG_3__3_ & n85284;
  assign n85663 = ~n85659 & ~n85660;
  assign n85664 = ~n85661 & n85663;
  assign n85665 = ~n85662 & n85664;
  assign n85666 = P2_P1_INSTQUEUE_REG_4__3_ & n85290;
  assign n85667 = P2_P1_INSTQUEUE_REG_5__3_ & n85292;
  assign n85668 = P2_P1_INSTQUEUE_REG_6__3_ & n85294;
  assign n85669 = P2_P1_INSTQUEUE_REG_7__3_ & n85296;
  assign n85670 = ~n85666 & ~n85667;
  assign n85671 = ~n85668 & n85670;
  assign n85672 = ~n85669 & n85671;
  assign n85673 = P2_P1_INSTQUEUE_REG_8__3_ & n85302;
  assign n85674 = P2_P1_INSTQUEUE_REG_9__3_ & n85304;
  assign n85675 = P2_P1_INSTQUEUE_REG_10__3_ & n85306;
  assign n85676 = P2_P1_INSTQUEUE_REG_11__3_ & n85308;
  assign n85677 = ~n85673 & ~n85674;
  assign n85678 = ~n85675 & n85677;
  assign n85679 = ~n85676 & n85678;
  assign n85680 = P2_P1_INSTQUEUE_REG_12__3_ & n85314;
  assign n85681 = P2_P1_INSTQUEUE_REG_13__3_ & n85316;
  assign n85682 = P2_P1_INSTQUEUE_REG_14__3_ & n85318;
  assign n85683 = P2_P1_INSTQUEUE_REG_15__3_ & n85320;
  assign n85684 = ~n85680 & ~n85681;
  assign n85685 = ~n85682 & n85684;
  assign n85686 = ~n85683 & n85685;
  assign n85687 = n85665 & n85672;
  assign n85688 = n85679 & n85687;
  assign n85689 = n85686 & n85688;
  assign n85690 = ~n85445 & ~n85565;
  assign n85691 = n85689 & ~n85690;
  assign n85692 = ~n85689 & n85690;
  assign n85693 = ~n85691 & ~n85692;
  assign n85694 = P2_P1_INSTADDRPOINTER_REG_3_ & ~n85693;
  assign n85695 = ~P2_P1_INSTADDRPOINTER_REG_3_ & n85693;
  assign n85696 = ~n85694 & ~n85695;
  assign n85697 = n85658 & ~n85696;
  assign n85698 = P2_P1_INSTADDRPOINTER_REG_3_ & n85693;
  assign n85699 = ~P2_P1_INSTADDRPOINTER_REG_3_ & ~n85693;
  assign n85700 = ~n85698 & ~n85699;
  assign n85701 = ~n85658 & ~n85700;
  assign n85702 = ~n85697 & ~n85701;
  assign n85703 = n85362 & ~n85702;
  assign n85704 = ~n85534 & ~n85583;
  assign n85705 = ~n85584 & ~n85704;
  assign n85706 = n85689 & n85690;
  assign n85707 = ~n85689 & ~n85690;
  assign n85708 = ~n85706 & ~n85707;
  assign n85709 = ~P2_P1_INSTADDRPOINTER_REG_3_ & n85708;
  assign n85710 = ~n85705 & ~n85709;
  assign n85711 = P2_P1_INSTADDRPOINTER_REG_3_ & ~n85708;
  assign n85712 = n85710 & ~n85711;
  assign n85713 = ~P2_P1_INSTADDRPOINTER_REG_3_ & ~n85708;
  assign n85714 = P2_P1_INSTADDRPOINTER_REG_3_ & n85708;
  assign n85715 = ~n85713 & ~n85714;
  assign n85716 = n85705 & n85715;
  assign n85717 = ~n85712 & ~n85716;
  assign n85718 = n85364 & n85717;
  assign n85719 = ~n85703 & ~n85718;
  assign n85720 = n85381 & ~n85639;
  assign n85721 = n85374 & ~n85639;
  assign n85722 = n85370 & ~n85639;
  assign n85723 = n77102 & ~n85639;
  assign n85724 = ~n85720 & ~n85721;
  assign n85725 = ~n85722 & n85724;
  assign n85726 = ~n85723 & n85725;
  assign n85727 = n76958 & ~n85647;
  assign n85728 = n77036 & ~n85647;
  assign n85729 = n77040 & ~n85647;
  assign n85730 = ~P2_P1_INSTADDRPOINTER_REG_3_ & n85600;
  assign n85731 = P2_P1_INSTADDRPOINTER_REG_3_ & ~n85600;
  assign n85732 = ~n85730 & ~n85731;
  assign n85733 = n77056 & n85732;
  assign n85734 = n77048 & n85732;
  assign n85735 = ~n85727 & ~n85728;
  assign n85736 = ~n85729 & n85735;
  assign n85737 = ~n85733 & n85736;
  assign n85738 = ~n85734 & n85737;
  assign n85739 = n85618 & ~n85621;
  assign n85740 = n85610 & n85689;
  assign n85741 = ~n85610 & ~n85689;
  assign n85742 = ~n85740 & ~n85741;
  assign n85743 = P2_P1_INSTADDRPOINTER_REG_3_ & n85742;
  assign n85744 = ~n85620 & n85742;
  assign n85745 = P2_P1_INSTADDRPOINTER_REG_3_ & ~n85620;
  assign n85746 = ~n85744 & ~n85745;
  assign n85747 = ~n85739 & ~n85743;
  assign n85748 = ~n85746 & n85747;
  assign n85749 = ~P2_P1_INSTADDRPOINTER_REG_3_ & n85742;
  assign n85750 = P2_P1_INSTADDRPOINTER_REG_3_ & ~n85742;
  assign n85751 = ~n85749 & ~n85750;
  assign n85752 = ~n85621 & n85751;
  assign n85753 = ~n85618 & ~n85620;
  assign n85754 = n85752 & ~n85753;
  assign n85755 = ~n85748 & ~n85754;
  assign n85756 = n77059 & n85755;
  assign n85757 = n85726 & n85738;
  assign n85758 = ~n85756 & n85757;
  assign n85759 = n85642 & ~n85643;
  assign n85760 = n85656 & n85759;
  assign n85761 = n85719 & n85760;
  assign n85762 = n85758 & n85761;
  assign n85763 = n85257 & ~n85762;
  assign n85764 = ~n85635 & ~n85636;
  assign n15546 = n85763 | ~n85764;
  assign n85766 = P2_P1_INSTADDRPOINTER_REG_4_ & n85256;
  assign n85767 = P2_P1_REIP_REG_4_ & n85401;
  assign n85768 = P2_P1_INSTADDRPOINTER_REG_3_ & n85601;
  assign n85769 = ~P2_P1_INSTADDRPOINTER_REG_4_ & n85768;
  assign n85770 = P2_P1_INSTADDRPOINTER_REG_4_ & ~n85768;
  assign n85771 = ~n85769 & ~n85770;
  assign n85772 = ~n77145 & ~n85771;
  assign n85773 = P2_P1_INSTADDRPOINTER_REG_3_ & n85644;
  assign n85774 = ~P2_P1_INSTADDRPOINTER_REG_4_ & n85773;
  assign n85775 = P2_P1_INSTADDRPOINTER_REG_4_ & ~n85773;
  assign n85776 = ~n85774 & ~n85775;
  assign n85777 = n77216 & ~n85776;
  assign n85778 = n77217 & ~n85776;
  assign n85779 = n85265 & ~n85771;
  assign n85780 = n85268 & ~n85771;
  assign n85781 = ~n85779 & ~n85780;
  assign n85782 = n77032 & ~n85776;
  assign n85783 = n85781 & ~n85782;
  assign n85784 = ~n85777 & ~n85778;
  assign n85785 = n85783 & n85784;
  assign n85786 = P2_P1_INSTQUEUE_REG_0__4_ & n85275;
  assign n85787 = P2_P1_INSTQUEUE_REG_1__4_ & n85278;
  assign n85788 = P2_P1_INSTQUEUE_REG_2__4_ & n85281;
  assign n85789 = P2_P1_INSTQUEUE_REG_3__4_ & n85284;
  assign n85790 = ~n85786 & ~n85787;
  assign n85791 = ~n85788 & n85790;
  assign n85792 = ~n85789 & n85791;
  assign n85793 = P2_P1_INSTQUEUE_REG_4__4_ & n85290;
  assign n85794 = P2_P1_INSTQUEUE_REG_5__4_ & n85292;
  assign n85795 = P2_P1_INSTQUEUE_REG_6__4_ & n85294;
  assign n85796 = P2_P1_INSTQUEUE_REG_7__4_ & n85296;
  assign n85797 = ~n85793 & ~n85794;
  assign n85798 = ~n85795 & n85797;
  assign n85799 = ~n85796 & n85798;
  assign n85800 = P2_P1_INSTQUEUE_REG_8__4_ & n85302;
  assign n85801 = P2_P1_INSTQUEUE_REG_9__4_ & n85304;
  assign n85802 = P2_P1_INSTQUEUE_REG_10__4_ & n85306;
  assign n85803 = P2_P1_INSTQUEUE_REG_11__4_ & n85308;
  assign n85804 = ~n85800 & ~n85801;
  assign n85805 = ~n85802 & n85804;
  assign n85806 = ~n85803 & n85805;
  assign n85807 = P2_P1_INSTQUEUE_REG_12__4_ & n85314;
  assign n85808 = P2_P1_INSTQUEUE_REG_13__4_ & n85316;
  assign n85809 = P2_P1_INSTQUEUE_REG_14__4_ & n85318;
  assign n85810 = P2_P1_INSTQUEUE_REG_15__4_ & n85320;
  assign n85811 = ~n85807 & ~n85808;
  assign n85812 = ~n85809 & n85811;
  assign n85813 = ~n85810 & n85812;
  assign n85814 = n85792 & n85799;
  assign n85815 = n85806 & n85814;
  assign n85816 = n85813 & n85815;
  assign n85817 = n85692 & n85816;
  assign n85818 = ~n85692 & ~n85816;
  assign n85819 = ~n85817 & ~n85818;
  assign n85820 = P2_P1_INSTADDRPOINTER_REG_4_ & ~n85819;
  assign n85821 = ~P2_P1_INSTADDRPOINTER_REG_4_ & n85819;
  assign n85822 = ~n85820 & ~n85821;
  assign n85823 = ~n85710 & ~n85711;
  assign n85824 = n85822 & ~n85823;
  assign n85825 = ~P2_P1_INSTADDRPOINTER_REG_4_ & ~n85819;
  assign n85826 = P2_P1_INSTADDRPOINTER_REG_4_ & n85819;
  assign n85827 = ~n85825 & ~n85826;
  assign n85828 = ~n85711 & n85827;
  assign n85829 = ~n85710 & n85828;
  assign n85830 = ~n85824 & ~n85829;
  assign n85831 = n85364 & n85830;
  assign n85832 = n77255 & ~n85771;
  assign n85833 = n77098 & ~n85771;
  assign n85834 = ~n85832 & ~n85833;
  assign n85835 = ~n85583 & ~n85699;
  assign n85836 = ~n85449 & ~n85579;
  assign n85837 = ~n85584 & n85836;
  assign n85838 = ~n85499 & n85837;
  assign n85839 = n85835 & ~n85838;
  assign n85840 = ~n85698 & ~n85839;
  assign n85841 = n85692 & ~n85816;
  assign n85842 = ~n85692 & n85816;
  assign n85843 = ~n85841 & ~n85842;
  assign n85844 = P2_P1_INSTADDRPOINTER_REG_4_ & ~n85843;
  assign n85845 = ~P2_P1_INSTADDRPOINTER_REG_4_ & n85843;
  assign n85846 = ~n85844 & ~n85845;
  assign n85847 = n85840 & ~n85846;
  assign n85848 = P2_P1_INSTADDRPOINTER_REG_4_ & n85843;
  assign n85849 = ~P2_P1_INSTADDRPOINTER_REG_4_ & ~n85843;
  assign n85850 = ~n85848 & ~n85849;
  assign n85851 = ~n85840 & ~n85850;
  assign n85852 = ~n85847 & ~n85851;
  assign n85853 = n85362 & ~n85852;
  assign n85854 = n85834 & ~n85853;
  assign n85855 = n85381 & ~n85771;
  assign n85856 = n85374 & ~n85771;
  assign n85857 = n85370 & ~n85771;
  assign n85858 = n77102 & ~n85771;
  assign n85859 = ~n85855 & ~n85856;
  assign n85860 = ~n85857 & n85859;
  assign n85861 = ~n85858 & n85860;
  assign n85862 = n76958 & ~n85776;
  assign n85863 = n77036 & ~n85776;
  assign n85864 = n77040 & ~n85776;
  assign n85865 = ~P2_P1_INSTADDRPOINTER_REG_4_ & n85731;
  assign n85866 = P2_P1_INSTADDRPOINTER_REG_4_ & ~n85731;
  assign n85867 = ~n85865 & ~n85866;
  assign n85868 = n77056 & ~n85867;
  assign n85869 = n77048 & ~n85867;
  assign n85870 = ~n85862 & ~n85863;
  assign n85871 = ~n85864 & n85870;
  assign n85872 = ~n85868 & n85871;
  assign n85873 = ~n85869 & n85872;
  assign n85874 = n85741 & n85816;
  assign n85875 = ~n85741 & ~n85816;
  assign n85876 = ~n85874 & ~n85875;
  assign n85877 = ~P2_P1_INSTADDRPOINTER_REG_4_ & ~n85876;
  assign n85878 = P2_P1_INSTADDRPOINTER_REG_4_ & n85876;
  assign n85879 = ~n85877 & ~n85878;
  assign n85880 = n85621 & n85742;
  assign n85881 = ~n85621 & ~n85742;
  assign n85882 = P2_P1_INSTADDRPOINTER_REG_3_ & ~n85881;
  assign n85883 = ~n85880 & ~n85882;
  assign n85884 = ~n85618 & ~n85746;
  assign n85885 = n85883 & ~n85884;
  assign n85886 = ~n85879 & n85885;
  assign n85887 = ~P2_P1_INSTADDRPOINTER_REG_4_ & n85876;
  assign n85888 = P2_P1_INSTADDRPOINTER_REG_4_ & ~n85876;
  assign n85889 = ~n85887 & ~n85888;
  assign n85890 = ~n85885 & ~n85889;
  assign n85891 = ~n85886 & ~n85890;
  assign n85892 = n77059 & ~n85891;
  assign n85893 = n85861 & n85873;
  assign n85894 = ~n85892 & n85893;
  assign n85895 = ~n85772 & n85785;
  assign n85896 = ~n85831 & n85895;
  assign n85897 = n85854 & n85896;
  assign n85898 = n85894 & n85897;
  assign n85899 = n85257 & ~n85898;
  assign n85900 = ~n85766 & ~n85767;
  assign n15551 = n85899 | ~n85900;
  assign n85902 = P2_P1_INSTADDRPOINTER_REG_5_ & n85256;
  assign n85903 = P2_P1_REIP_REG_5_ & n85401;
  assign n85904 = P2_P1_INSTADDRPOINTER_REG_4_ & n85773;
  assign n85905 = ~P2_P1_INSTADDRPOINTER_REG_5_ & n85904;
  assign n85906 = P2_P1_INSTADDRPOINTER_REG_5_ & ~n85904;
  assign n85907 = ~n85905 & ~n85906;
  assign n85908 = n77216 & ~n85907;
  assign n85909 = n77217 & ~n85907;
  assign n85910 = P2_P1_INSTADDRPOINTER_REG_4_ & n85768;
  assign n85911 = ~P2_P1_INSTADDRPOINTER_REG_5_ & n85910;
  assign n85912 = P2_P1_INSTADDRPOINTER_REG_5_ & ~n85910;
  assign n85913 = ~n85911 & ~n85912;
  assign n85914 = n85265 & ~n85913;
  assign n85915 = n85268 & ~n85913;
  assign n85916 = ~n85914 & ~n85915;
  assign n85917 = n77032 & ~n85907;
  assign n85918 = n85916 & ~n85917;
  assign n85919 = ~n85908 & ~n85909;
  assign n85920 = n85918 & n85919;
  assign n85921 = ~n77145 & ~n85913;
  assign n85922 = n85698 & ~n85849;
  assign n85923 = ~n85848 & ~n85922;
  assign n85924 = n85835 & ~n85849;
  assign n85925 = ~n85838 & n85924;
  assign n85926 = n85923 & ~n85925;
  assign n85927 = P2_P1_INSTQUEUE_REG_0__5_ & n85275;
  assign n85928 = P2_P1_INSTQUEUE_REG_1__5_ & n85278;
  assign n85929 = P2_P1_INSTQUEUE_REG_2__5_ & n85281;
  assign n85930 = P2_P1_INSTQUEUE_REG_3__5_ & n85284;
  assign n85931 = ~n85927 & ~n85928;
  assign n85932 = ~n85929 & n85931;
  assign n85933 = ~n85930 & n85932;
  assign n85934 = P2_P1_INSTQUEUE_REG_4__5_ & n85290;
  assign n85935 = P2_P1_INSTQUEUE_REG_5__5_ & n85292;
  assign n85936 = P2_P1_INSTQUEUE_REG_6__5_ & n85294;
  assign n85937 = P2_P1_INSTQUEUE_REG_7__5_ & n85296;
  assign n85938 = ~n85934 & ~n85935;
  assign n85939 = ~n85936 & n85938;
  assign n85940 = ~n85937 & n85939;
  assign n85941 = P2_P1_INSTQUEUE_REG_8__5_ & n85302;
  assign n85942 = P2_P1_INSTQUEUE_REG_9__5_ & n85304;
  assign n85943 = P2_P1_INSTQUEUE_REG_10__5_ & n85306;
  assign n85944 = P2_P1_INSTQUEUE_REG_11__5_ & n85308;
  assign n85945 = ~n85941 & ~n85942;
  assign n85946 = ~n85943 & n85945;
  assign n85947 = ~n85944 & n85946;
  assign n85948 = P2_P1_INSTQUEUE_REG_12__5_ & n85314;
  assign n85949 = P2_P1_INSTQUEUE_REG_13__5_ & n85316;
  assign n85950 = P2_P1_INSTQUEUE_REG_14__5_ & n85318;
  assign n85951 = P2_P1_INSTQUEUE_REG_15__5_ & n85320;
  assign n85952 = ~n85948 & ~n85949;
  assign n85953 = ~n85950 & n85952;
  assign n85954 = ~n85951 & n85953;
  assign n85955 = n85933 & n85940;
  assign n85956 = n85947 & n85955;
  assign n85957 = n85954 & n85956;
  assign n85958 = ~n85841 & n85957;
  assign n85959 = ~n85816 & ~n85957;
  assign n85960 = n85692 & n85959;
  assign n85961 = ~n85958 & ~n85960;
  assign n85962 = P2_P1_INSTADDRPOINTER_REG_5_ & ~n85961;
  assign n85963 = ~P2_P1_INSTADDRPOINTER_REG_5_ & n85961;
  assign n85964 = ~n85962 & ~n85963;
  assign n85965 = n85926 & ~n85964;
  assign n85966 = ~n85926 & n85964;
  assign n85967 = ~n85965 & ~n85966;
  assign n85968 = n85362 & ~n85967;
  assign n85969 = n77255 & ~n85913;
  assign n85970 = n77098 & ~n85913;
  assign n85971 = ~n85969 & ~n85970;
  assign n85972 = n85711 & ~n85821;
  assign n85973 = ~n85820 & ~n85972;
  assign n85974 = ~n85709 & ~n85821;
  assign n85975 = ~n85705 & n85974;
  assign n85976 = n85973 & ~n85975;
  assign n85977 = n85841 & n85957;
  assign n85978 = ~n85841 & ~n85957;
  assign n85979 = ~n85977 & ~n85978;
  assign n85980 = ~P2_P1_INSTADDRPOINTER_REG_5_ & ~n85979;
  assign n85981 = P2_P1_INSTADDRPOINTER_REG_5_ & n85979;
  assign n85982 = ~n85980 & ~n85981;
  assign n85983 = n85976 & ~n85982;
  assign n85984 = ~n85976 & n85982;
  assign n85985 = ~n85983 & ~n85984;
  assign n85986 = n85364 & ~n85985;
  assign n85987 = n85971 & ~n85986;
  assign n85988 = n85381 & ~n85913;
  assign n85989 = n85374 & ~n85913;
  assign n85990 = n85370 & ~n85913;
  assign n85991 = n77102 & ~n85913;
  assign n85992 = ~n85988 & ~n85989;
  assign n85993 = ~n85990 & n85992;
  assign n85994 = ~n85991 & n85993;
  assign n85995 = n76958 & ~n85907;
  assign n85996 = n77036 & ~n85907;
  assign n85997 = n77040 & ~n85907;
  assign n85998 = P2_P1_INSTADDRPOINTER_REG_4_ & n85731;
  assign n85999 = ~P2_P1_INSTADDRPOINTER_REG_5_ & n85998;
  assign n86000 = P2_P1_INSTADDRPOINTER_REG_5_ & ~n85998;
  assign n86001 = ~n85999 & ~n86000;
  assign n86002 = n77056 & ~n86001;
  assign n86003 = n77048 & ~n86001;
  assign n86004 = ~n85995 & ~n85996;
  assign n86005 = ~n85997 & n86004;
  assign n86006 = ~n86002 & n86005;
  assign n86007 = ~n86003 & n86006;
  assign n86008 = n85741 & ~n85816;
  assign n86009 = n85957 & n86008;
  assign n86010 = ~n85957 & ~n86008;
  assign n86011 = ~n86009 & ~n86010;
  assign n86012 = P2_P1_INSTADDRPOINTER_REG_5_ & ~n86011;
  assign n86013 = ~P2_P1_INSTADDRPOINTER_REG_5_ & n86011;
  assign n86014 = ~n85887 & ~n86013;
  assign n86015 = ~n86012 & n86014;
  assign n86016 = n85885 & ~n85888;
  assign n86017 = n86015 & ~n86016;
  assign n86018 = ~P2_P1_INSTADDRPOINTER_REG_5_ & ~n86011;
  assign n86019 = P2_P1_INSTADDRPOINTER_REG_5_ & n86011;
  assign n86020 = ~n86018 & ~n86019;
  assign n86021 = ~n85888 & n86020;
  assign n86022 = ~n85885 & ~n85887;
  assign n86023 = n86021 & ~n86022;
  assign n86024 = ~n86017 & ~n86023;
  assign n86025 = n77059 & n86024;
  assign n86026 = n85994 & n86007;
  assign n86027 = ~n86025 & n86026;
  assign n86028 = n85920 & ~n85921;
  assign n86029 = ~n85968 & n86028;
  assign n86030 = n85987 & n86029;
  assign n86031 = n86027 & n86030;
  assign n86032 = n85257 & ~n86031;
  assign n86033 = ~n85902 & ~n85903;
  assign n15556 = n86032 | ~n86033;
  assign n86035 = P2_P1_INSTADDRPOINTER_REG_6_ & n85256;
  assign n86036 = P2_P1_REIP_REG_6_ & n85401;
  assign n86037 = P2_P1_INSTADDRPOINTER_REG_5_ & n85904;
  assign n86038 = ~P2_P1_INSTADDRPOINTER_REG_6_ & n86037;
  assign n86039 = P2_P1_INSTADDRPOINTER_REG_6_ & ~n86037;
  assign n86040 = ~n86038 & ~n86039;
  assign n86041 = n77216 & ~n86040;
  assign n86042 = n77217 & ~n86040;
  assign n86043 = P2_P1_INSTADDRPOINTER_REG_5_ & n85910;
  assign n86044 = ~P2_P1_INSTADDRPOINTER_REG_6_ & n86043;
  assign n86045 = P2_P1_INSTADDRPOINTER_REG_6_ & ~n86043;
  assign n86046 = ~n86044 & ~n86045;
  assign n86047 = n85265 & ~n86046;
  assign n86048 = n85268 & ~n86046;
  assign n86049 = ~n86047 & ~n86048;
  assign n86050 = n77032 & ~n86040;
  assign n86051 = n86049 & ~n86050;
  assign n86052 = ~n86041 & ~n86042;
  assign n86053 = n86051 & n86052;
  assign n86054 = ~n77145 & ~n86046;
  assign n86055 = ~P2_P1_INSTADDRPOINTER_REG_5_ & ~n85961;
  assign n86056 = ~n85926 & ~n86055;
  assign n86057 = P2_P1_INSTADDRPOINTER_REG_5_ & n85961;
  assign n86058 = ~n86056 & ~n86057;
  assign n86059 = P2_P1_INSTQUEUE_REG_0__6_ & n85275;
  assign n86060 = P2_P1_INSTQUEUE_REG_1__6_ & n85278;
  assign n86061 = P2_P1_INSTQUEUE_REG_2__6_ & n85281;
  assign n86062 = P2_P1_INSTQUEUE_REG_3__6_ & n85284;
  assign n86063 = ~n86059 & ~n86060;
  assign n86064 = ~n86061 & n86063;
  assign n86065 = ~n86062 & n86064;
  assign n86066 = P2_P1_INSTQUEUE_REG_4__6_ & n85290;
  assign n86067 = P2_P1_INSTQUEUE_REG_5__6_ & n85292;
  assign n86068 = P2_P1_INSTQUEUE_REG_6__6_ & n85294;
  assign n86069 = P2_P1_INSTQUEUE_REG_7__6_ & n85296;
  assign n86070 = ~n86066 & ~n86067;
  assign n86071 = ~n86068 & n86070;
  assign n86072 = ~n86069 & n86071;
  assign n86073 = P2_P1_INSTQUEUE_REG_8__6_ & n85302;
  assign n86074 = P2_P1_INSTQUEUE_REG_9__6_ & n85304;
  assign n86075 = P2_P1_INSTQUEUE_REG_10__6_ & n85306;
  assign n86076 = P2_P1_INSTQUEUE_REG_11__6_ & n85308;
  assign n86077 = ~n86073 & ~n86074;
  assign n86078 = ~n86075 & n86077;
  assign n86079 = ~n86076 & n86078;
  assign n86080 = P2_P1_INSTQUEUE_REG_12__6_ & n85314;
  assign n86081 = P2_P1_INSTQUEUE_REG_13__6_ & n85316;
  assign n86082 = P2_P1_INSTQUEUE_REG_14__6_ & n85318;
  assign n86083 = P2_P1_INSTQUEUE_REG_15__6_ & n85320;
  assign n86084 = ~n86080 & ~n86081;
  assign n86085 = ~n86082 & n86084;
  assign n86086 = ~n86083 & n86085;
  assign n86087 = n86065 & n86072;
  assign n86088 = n86079 & n86087;
  assign n86089 = n86086 & n86088;
  assign n86090 = n85960 & ~n86089;
  assign n86091 = ~n85960 & n86089;
  assign n86092 = ~n86090 & ~n86091;
  assign n86093 = P2_P1_INSTADDRPOINTER_REG_6_ & ~n86092;
  assign n86094 = ~P2_P1_INSTADDRPOINTER_REG_6_ & n86092;
  assign n86095 = ~n86093 & ~n86094;
  assign n86096 = n86058 & ~n86095;
  assign n86097 = ~n86058 & n86095;
  assign n86098 = ~n86096 & ~n86097;
  assign n86099 = n85362 & ~n86098;
  assign n86100 = n77255 & ~n86046;
  assign n86101 = n77098 & ~n86046;
  assign n86102 = ~n86100 & ~n86101;
  assign n86103 = ~n85976 & ~n85979;
  assign n86104 = P2_P1_INSTADDRPOINTER_REG_5_ & ~n85976;
  assign n86105 = P2_P1_INSTADDRPOINTER_REG_5_ & ~n85979;
  assign n86106 = ~n86103 & ~n86104;
  assign n86107 = ~n86105 & n86106;
  assign n86108 = n85841 & ~n85957;
  assign n86109 = n86089 & n86108;
  assign n86110 = ~n86089 & ~n86108;
  assign n86111 = ~n86109 & ~n86110;
  assign n86112 = ~P2_P1_INSTADDRPOINTER_REG_6_ & ~n86111;
  assign n86113 = P2_P1_INSTADDRPOINTER_REG_6_ & n86111;
  assign n86114 = ~n86112 & ~n86113;
  assign n86115 = n86107 & ~n86114;
  assign n86116 = ~n86107 & n86114;
  assign n86117 = ~n86115 & ~n86116;
  assign n86118 = n85364 & ~n86117;
  assign n86119 = n86102 & ~n86118;
  assign n86120 = n85381 & ~n86046;
  assign n86121 = n85374 & ~n86046;
  assign n86122 = n85370 & ~n86046;
  assign n86123 = n77102 & ~n86046;
  assign n86124 = ~n86120 & ~n86121;
  assign n86125 = ~n86122 & n86124;
  assign n86126 = ~n86123 & n86125;
  assign n86127 = n76958 & ~n86040;
  assign n86128 = n77036 & ~n86040;
  assign n86129 = n77040 & ~n86040;
  assign n86130 = P2_P1_INSTADDRPOINTER_REG_5_ & n85998;
  assign n86131 = ~P2_P1_INSTADDRPOINTER_REG_6_ & n86130;
  assign n86132 = P2_P1_INSTADDRPOINTER_REG_6_ & ~n86130;
  assign n86133 = ~n86131 & ~n86132;
  assign n86134 = n77056 & ~n86133;
  assign n86135 = n77048 & ~n86133;
  assign n86136 = ~n86127 & ~n86128;
  assign n86137 = ~n86129 & n86136;
  assign n86138 = ~n86134 & n86137;
  assign n86139 = ~n86135 & n86138;
  assign n86140 = n85888 & ~n86011;
  assign n86141 = ~n85888 & n86011;
  assign n86142 = P2_P1_INSTADDRPOINTER_REG_5_ & ~n86141;
  assign n86143 = ~n86140 & ~n86142;
  assign n86144 = ~n85885 & n86014;
  assign n86145 = n86143 & ~n86144;
  assign n86146 = ~n85957 & n86008;
  assign n86147 = n86089 & n86146;
  assign n86148 = ~n86089 & ~n86146;
  assign n86149 = ~n86147 & ~n86148;
  assign n86150 = ~P2_P1_INSTADDRPOINTER_REG_6_ & ~n86149;
  assign n86151 = P2_P1_INSTADDRPOINTER_REG_6_ & n86149;
  assign n86152 = ~n86150 & ~n86151;
  assign n86153 = n86145 & ~n86152;
  assign n86154 = ~n86145 & n86152;
  assign n86155 = ~n86153 & ~n86154;
  assign n86156 = n77059 & ~n86155;
  assign n86157 = n86126 & n86139;
  assign n86158 = ~n86156 & n86157;
  assign n86159 = n86053 & ~n86054;
  assign n86160 = ~n86099 & n86159;
  assign n86161 = n86119 & n86160;
  assign n86162 = n86158 & n86161;
  assign n86163 = n85257 & ~n86162;
  assign n86164 = ~n86035 & ~n86036;
  assign n15561 = n86163 | ~n86164;
  assign n86166 = P2_P1_INSTADDRPOINTER_REG_7_ & n85256;
  assign n86167 = P2_P1_REIP_REG_7_ & n85401;
  assign n86168 = P2_P1_INSTADDRPOINTER_REG_6_ & n86037;
  assign n86169 = ~P2_P1_INSTADDRPOINTER_REG_7_ & n86168;
  assign n86170 = P2_P1_INSTADDRPOINTER_REG_7_ & ~n86168;
  assign n86171 = ~n86169 & ~n86170;
  assign n86172 = n77216 & ~n86171;
  assign n86173 = n77217 & ~n86171;
  assign n86174 = P2_P1_INSTADDRPOINTER_REG_6_ & n86043;
  assign n86175 = ~P2_P1_INSTADDRPOINTER_REG_7_ & n86174;
  assign n86176 = P2_P1_INSTADDRPOINTER_REG_7_ & ~n86174;
  assign n86177 = ~n86175 & ~n86176;
  assign n86178 = n85265 & ~n86177;
  assign n86179 = n85268 & ~n86177;
  assign n86180 = ~n86178 & ~n86179;
  assign n86181 = n77032 & ~n86171;
  assign n86182 = n86180 & ~n86181;
  assign n86183 = ~n86172 & ~n86173;
  assign n86184 = n86182 & n86183;
  assign n86185 = ~n77145 & ~n86177;
  assign n86186 = P2_P1_INSTADDRPOINTER_REG_6_ & n86092;
  assign n86187 = ~P2_P1_INSTADDRPOINTER_REG_6_ & ~n86092;
  assign n86188 = ~n86058 & ~n86187;
  assign n86189 = ~n86186 & ~n86188;
  assign n86190 = n85361 & ~n86090;
  assign n86191 = ~n85361 & ~n86089;
  assign n86192 = n85960 & n86191;
  assign n86193 = ~n86190 & ~n86192;
  assign n86194 = P2_P1_INSTADDRPOINTER_REG_7_ & ~n86193;
  assign n86195 = ~P2_P1_INSTADDRPOINTER_REG_7_ & n86193;
  assign n86196 = ~n86194 & ~n86195;
  assign n86197 = n86189 & ~n86196;
  assign n86198 = ~n86189 & n86196;
  assign n86199 = ~n86197 & ~n86198;
  assign n86200 = n85362 & ~n86199;
  assign n86201 = n77255 & ~n86177;
  assign n86202 = n77098 & ~n86177;
  assign n86203 = ~n86201 & ~n86202;
  assign n86204 = P2_P1_INSTADDRPOINTER_REG_6_ & ~n86111;
  assign n86205 = ~P2_P1_INSTADDRPOINTER_REG_6_ & n86111;
  assign n86206 = ~n86107 & ~n86205;
  assign n86207 = ~n86204 & ~n86206;
  assign n86208 = ~n86089 & n86108;
  assign n86209 = n85361 & n86208;
  assign n86210 = ~n85361 & ~n86208;
  assign n86211 = ~n86209 & ~n86210;
  assign n86212 = ~P2_P1_INSTADDRPOINTER_REG_7_ & ~n86211;
  assign n86213 = P2_P1_INSTADDRPOINTER_REG_7_ & n86211;
  assign n86214 = ~n86212 & ~n86213;
  assign n86215 = n86207 & ~n86214;
  assign n86216 = ~n86207 & n86214;
  assign n86217 = ~n86215 & ~n86216;
  assign n86218 = n85364 & ~n86217;
  assign n86219 = n86203 & ~n86218;
  assign n86220 = n85381 & ~n86177;
  assign n86221 = n85374 & ~n86177;
  assign n86222 = n85370 & ~n86177;
  assign n86223 = n77102 & ~n86177;
  assign n86224 = ~n86220 & ~n86221;
  assign n86225 = ~n86222 & n86224;
  assign n86226 = ~n86223 & n86225;
  assign n86227 = n76958 & ~n86171;
  assign n86228 = n77036 & ~n86171;
  assign n86229 = n77040 & ~n86171;
  assign n86230 = P2_P1_INSTADDRPOINTER_REG_6_ & n86130;
  assign n86231 = ~P2_P1_INSTADDRPOINTER_REG_7_ & n86230;
  assign n86232 = P2_P1_INSTADDRPOINTER_REG_7_ & ~n86230;
  assign n86233 = ~n86231 & ~n86232;
  assign n86234 = n77056 & ~n86233;
  assign n86235 = n77048 & ~n86233;
  assign n86236 = ~n86227 & ~n86228;
  assign n86237 = ~n86229 & n86236;
  assign n86238 = ~n86234 & n86237;
  assign n86239 = ~n86235 & n86238;
  assign n86240 = P2_P1_INSTADDRPOINTER_REG_6_ & ~n86149;
  assign n86241 = ~P2_P1_INSTADDRPOINTER_REG_6_ & n86149;
  assign n86242 = ~n86145 & ~n86241;
  assign n86243 = ~n86240 & ~n86242;
  assign n86244 = ~n86089 & n86146;
  assign n86245 = n85361 & n86244;
  assign n86246 = ~n85361 & ~n86244;
  assign n86247 = ~n86245 & ~n86246;
  assign n86248 = ~P2_P1_INSTADDRPOINTER_REG_7_ & ~n86247;
  assign n86249 = P2_P1_INSTADDRPOINTER_REG_7_ & n86247;
  assign n86250 = ~n86248 & ~n86249;
  assign n86251 = n86243 & ~n86250;
  assign n86252 = ~n86243 & n86250;
  assign n86253 = ~n86251 & ~n86252;
  assign n86254 = n77059 & ~n86253;
  assign n86255 = n86226 & n86239;
  assign n86256 = ~n86254 & n86255;
  assign n86257 = n86184 & ~n86185;
  assign n86258 = ~n86200 & n86257;
  assign n86259 = n86219 & n86258;
  assign n86260 = n86256 & n86259;
  assign n86261 = n85257 & ~n86260;
  assign n86262 = ~n86166 & ~n86167;
  assign n15566 = n86261 | ~n86262;
  assign n86264 = P2_P1_INSTADDRPOINTER_REG_8_ & n85256;
  assign n86265 = P2_P1_REIP_REG_8_ & n85401;
  assign n86266 = P2_P1_INSTADDRPOINTER_REG_7_ & n86168;
  assign n86267 = ~P2_P1_INSTADDRPOINTER_REG_8_ & n86266;
  assign n86268 = P2_P1_INSTADDRPOINTER_REG_8_ & ~n86266;
  assign n86269 = ~n86267 & ~n86268;
  assign n86270 = n77216 & ~n86269;
  assign n86271 = n77217 & ~n86269;
  assign n86272 = n77032 & ~n86269;
  assign n86273 = P2_P1_INSTADDRPOINTER_REG_7_ & n86174;
  assign n86274 = ~P2_P1_INSTADDRPOINTER_REG_8_ & n86273;
  assign n86275 = P2_P1_INSTADDRPOINTER_REG_8_ & ~n86273;
  assign n86276 = ~n86274 & ~n86275;
  assign n86277 = n85268 & ~n86276;
  assign n86278 = n85265 & ~n86276;
  assign n86279 = ~n86272 & ~n86277;
  assign n86280 = ~n86278 & n86279;
  assign n86281 = ~n86270 & ~n86271;
  assign n86282 = n86280 & n86281;
  assign n86283 = ~n77145 & ~n86276;
  assign n86284 = ~P2_P1_INSTADDRPOINTER_REG_7_ & ~n86193;
  assign n86285 = ~n86189 & ~n86284;
  assign n86286 = P2_P1_INSTADDRPOINTER_REG_7_ & n86193;
  assign n86287 = ~n86285 & ~n86286;
  assign n86288 = ~P2_P1_INSTADDRPOINTER_REG_8_ & ~n86192;
  assign n86289 = P2_P1_INSTADDRPOINTER_REG_8_ & n86192;
  assign n86290 = ~n86288 & ~n86289;
  assign n86291 = n86287 & ~n86290;
  assign n86292 = ~n86287 & n86290;
  assign n86293 = ~n86291 & ~n86292;
  assign n86294 = n85362 & ~n86293;
  assign n86295 = n77255 & ~n86276;
  assign n86296 = n77098 & ~n86276;
  assign n86297 = ~n86295 & ~n86296;
  assign n86298 = ~n86207 & ~n86211;
  assign n86299 = P2_P1_INSTADDRPOINTER_REG_7_ & ~n86207;
  assign n86300 = P2_P1_INSTADDRPOINTER_REG_7_ & ~n86211;
  assign n86301 = ~n86298 & ~n86299;
  assign n86302 = ~n86300 & n86301;
  assign n86303 = n86108 & n86191;
  assign n86304 = ~P2_P1_INSTADDRPOINTER_REG_8_ & n86303;
  assign n86305 = P2_P1_INSTADDRPOINTER_REG_8_ & ~n86303;
  assign n86306 = ~n86304 & ~n86305;
  assign n86307 = n86302 & ~n86306;
  assign n86308 = ~n86302 & n86306;
  assign n86309 = ~n86307 & ~n86308;
  assign n86310 = n85364 & ~n86309;
  assign n86311 = n86297 & ~n86310;
  assign n86312 = n85381 & ~n86276;
  assign n86313 = n77102 & ~n86276;
  assign n86314 = n85370 & ~n86276;
  assign n86315 = n85374 & ~n86276;
  assign n86316 = ~n86312 & ~n86313;
  assign n86317 = ~n86314 & n86316;
  assign n86318 = ~n86315 & n86317;
  assign n86319 = n76958 & ~n86269;
  assign n86320 = n77036 & ~n86269;
  assign n86321 = n77040 & ~n86269;
  assign n86322 = P2_P1_INSTADDRPOINTER_REG_7_ & n86230;
  assign n86323 = ~P2_P1_INSTADDRPOINTER_REG_8_ & n86322;
  assign n86324 = P2_P1_INSTADDRPOINTER_REG_8_ & ~n86322;
  assign n86325 = ~n86323 & ~n86324;
  assign n86326 = n77056 & ~n86325;
  assign n86327 = n77048 & ~n86325;
  assign n86328 = ~n86319 & ~n86320;
  assign n86329 = ~n86321 & n86328;
  assign n86330 = ~n86326 & n86329;
  assign n86331 = ~n86327 & n86330;
  assign n86332 = ~n86243 & ~n86247;
  assign n86333 = P2_P1_INSTADDRPOINTER_REG_7_ & ~n86243;
  assign n86334 = P2_P1_INSTADDRPOINTER_REG_7_ & ~n86247;
  assign n86335 = ~n86332 & ~n86333;
  assign n86336 = ~n86334 & n86335;
  assign n86337 = n86146 & n86191;
  assign n86338 = ~P2_P1_INSTADDRPOINTER_REG_8_ & n86337;
  assign n86339 = P2_P1_INSTADDRPOINTER_REG_8_ & ~n86337;
  assign n86340 = ~n86338 & ~n86339;
  assign n86341 = n86336 & ~n86340;
  assign n86342 = ~n86336 & n86340;
  assign n86343 = ~n86341 & ~n86342;
  assign n86344 = n77059 & ~n86343;
  assign n86345 = n86318 & n86331;
  assign n86346 = ~n86344 & n86345;
  assign n86347 = n86282 & ~n86283;
  assign n86348 = ~n86294 & n86347;
  assign n86349 = n86311 & n86348;
  assign n86350 = n86346 & n86349;
  assign n86351 = n85257 & ~n86350;
  assign n86352 = ~n86264 & ~n86265;
  assign n15571 = n86351 | ~n86352;
  assign n86354 = P2_P1_INSTADDRPOINTER_REG_9_ & n85256;
  assign n86355 = P2_P1_REIP_REG_9_ & n85401;
  assign n86356 = P2_P1_INSTADDRPOINTER_REG_8_ & n86266;
  assign n86357 = ~P2_P1_INSTADDRPOINTER_REG_9_ & n86356;
  assign n86358 = P2_P1_INSTADDRPOINTER_REG_9_ & ~n86356;
  assign n86359 = ~n86357 & ~n86358;
  assign n86360 = n77216 & ~n86359;
  assign n86361 = n77217 & ~n86359;
  assign n86362 = P2_P1_INSTADDRPOINTER_REG_8_ & n86273;
  assign n86363 = ~P2_P1_INSTADDRPOINTER_REG_9_ & n86362;
  assign n86364 = P2_P1_INSTADDRPOINTER_REG_9_ & ~n86362;
  assign n86365 = ~n86363 & ~n86364;
  assign n86366 = n85265 & ~n86365;
  assign n86367 = n77032 & ~n86359;
  assign n86368 = n85268 & ~n86365;
  assign n86369 = ~n86367 & ~n86368;
  assign n86370 = ~n86360 & ~n86361;
  assign n86371 = ~n86366 & n86370;
  assign n86372 = n86369 & n86371;
  assign n86373 = ~n77145 & ~n86365;
  assign n86374 = ~P2_P1_INSTADDRPOINTER_REG_8_ & n86192;
  assign n86375 = ~n86287 & ~n86374;
  assign n86376 = P2_P1_INSTADDRPOINTER_REG_8_ & ~n86192;
  assign n86377 = ~n86375 & ~n86376;
  assign n86378 = P2_P1_INSTADDRPOINTER_REG_9_ & n86192;
  assign n86379 = ~P2_P1_INSTADDRPOINTER_REG_9_ & ~n86192;
  assign n86380 = ~n86378 & ~n86379;
  assign n86381 = n86377 & ~n86380;
  assign n86382 = P2_P1_INSTADDRPOINTER_REG_9_ & ~n86192;
  assign n86383 = ~P2_P1_INSTADDRPOINTER_REG_9_ & n86192;
  assign n86384 = ~n86382 & ~n86383;
  assign n86385 = ~n86377 & ~n86384;
  assign n86386 = ~n86381 & ~n86385;
  assign n86387 = n85362 & ~n86386;
  assign n86388 = n77255 & ~n86365;
  assign n86389 = n77098 & ~n86365;
  assign n86390 = ~n86388 & ~n86389;
  assign n86391 = P2_P1_INSTADDRPOINTER_REG_8_ & n86303;
  assign n86392 = ~P2_P1_INSTADDRPOINTER_REG_8_ & ~n86303;
  assign n86393 = ~n86302 & ~n86392;
  assign n86394 = ~n86391 & ~n86393;
  assign n86395 = ~P2_P1_INSTADDRPOINTER_REG_9_ & n86394;
  assign n86396 = P2_P1_INSTADDRPOINTER_REG_9_ & ~n86394;
  assign n86397 = ~n86395 & ~n86396;
  assign n86398 = n85364 & n86397;
  assign n86399 = n86390 & ~n86398;
  assign n86400 = n85381 & ~n86365;
  assign n86401 = n77102 & ~n86365;
  assign n86402 = n85370 & ~n86365;
  assign n86403 = n85374 & ~n86365;
  assign n86404 = ~n86400 & ~n86401;
  assign n86405 = ~n86402 & n86404;
  assign n86406 = ~n86403 & n86405;
  assign n86407 = n76958 & ~n86359;
  assign n86408 = n77036 & ~n86359;
  assign n86409 = n77040 & ~n86359;
  assign n86410 = P2_P1_INSTADDRPOINTER_REG_8_ & n86322;
  assign n86411 = ~P2_P1_INSTADDRPOINTER_REG_9_ & n86410;
  assign n86412 = P2_P1_INSTADDRPOINTER_REG_9_ & ~n86410;
  assign n86413 = ~n86411 & ~n86412;
  assign n86414 = n77056 & ~n86413;
  assign n86415 = n77048 & ~n86413;
  assign n86416 = ~n86407 & ~n86408;
  assign n86417 = ~n86409 & n86416;
  assign n86418 = ~n86414 & n86417;
  assign n86419 = ~n86415 & n86418;
  assign n86420 = P2_P1_INSTADDRPOINTER_REG_8_ & n86337;
  assign n86421 = ~P2_P1_INSTADDRPOINTER_REG_8_ & ~n86337;
  assign n86422 = ~n86336 & ~n86421;
  assign n86423 = ~n86420 & ~n86422;
  assign n86424 = ~P2_P1_INSTADDRPOINTER_REG_9_ & n86423;
  assign n86425 = P2_P1_INSTADDRPOINTER_REG_9_ & ~n86423;
  assign n86426 = ~n86424 & ~n86425;
  assign n86427 = n77059 & n86426;
  assign n86428 = n86406 & n86419;
  assign n86429 = ~n86427 & n86428;
  assign n86430 = n86372 & ~n86373;
  assign n86431 = ~n86387 & n86430;
  assign n86432 = n86399 & n86431;
  assign n86433 = n86429 & n86432;
  assign n86434 = n85257 & ~n86433;
  assign n86435 = ~n86354 & ~n86355;
  assign n15576 = n86434 | ~n86435;
  assign n86437 = P2_P1_INSTADDRPOINTER_REG_10_ & n85256;
  assign n86438 = P2_P1_REIP_REG_10_ & n85401;
  assign n86439 = P2_P1_INSTADDRPOINTER_REG_9_ & n86356;
  assign n86440 = ~P2_P1_INSTADDRPOINTER_REG_10_ & n86439;
  assign n86441 = P2_P1_INSTADDRPOINTER_REG_10_ & ~n86439;
  assign n86442 = ~n86440 & ~n86441;
  assign n86443 = n77216 & ~n86442;
  assign n86444 = n77217 & ~n86442;
  assign n86445 = P2_P1_INSTADDRPOINTER_REG_9_ & n86362;
  assign n86446 = ~P2_P1_INSTADDRPOINTER_REG_10_ & n86445;
  assign n86447 = P2_P1_INSTADDRPOINTER_REG_10_ & ~n86445;
  assign n86448 = ~n86446 & ~n86447;
  assign n86449 = n85265 & ~n86448;
  assign n86450 = n77032 & ~n86442;
  assign n86451 = n85268 & ~n86448;
  assign n86452 = ~n86450 & ~n86451;
  assign n86453 = ~n86443 & ~n86444;
  assign n86454 = ~n86449 & n86453;
  assign n86455 = n86452 & n86454;
  assign n86456 = ~n77145 & ~n86448;
  assign n86457 = ~n86374 & ~n86383;
  assign n86458 = ~n86287 & n86457;
  assign n86459 = ~n86376 & ~n86382;
  assign n86460 = ~n86458 & n86459;
  assign n86461 = ~P2_P1_INSTADDRPOINTER_REG_10_ & ~n86192;
  assign n86462 = P2_P1_INSTADDRPOINTER_REG_10_ & n86192;
  assign n86463 = ~n86461 & ~n86462;
  assign n86464 = n86460 & ~n86463;
  assign n86465 = P2_P1_INSTADDRPOINTER_REG_10_ & ~n86192;
  assign n86466 = ~P2_P1_INSTADDRPOINTER_REG_10_ & n86192;
  assign n86467 = ~n86465 & ~n86466;
  assign n86468 = ~n86460 & ~n86467;
  assign n86469 = ~n86464 & ~n86468;
  assign n86470 = n85362 & ~n86469;
  assign n86471 = n77255 & ~n86448;
  assign n86472 = n77098 & ~n86448;
  assign n86473 = ~n86471 & ~n86472;
  assign n86474 = ~P2_P1_INSTADDRPOINTER_REG_10_ & ~n86396;
  assign n86475 = P2_P1_INSTADDRPOINTER_REG_9_ & P2_P1_INSTADDRPOINTER_REG_10_;
  assign n86476 = ~n86394 & n86475;
  assign n86477 = ~n86474 & ~n86476;
  assign n86478 = n85364 & n86477;
  assign n86479 = n86473 & ~n86478;
  assign n86480 = n85381 & ~n86448;
  assign n86481 = n77102 & ~n86448;
  assign n86482 = n85370 & ~n86448;
  assign n86483 = n85374 & ~n86448;
  assign n86484 = ~n86480 & ~n86481;
  assign n86485 = ~n86482 & n86484;
  assign n86486 = ~n86483 & n86485;
  assign n86487 = n76958 & ~n86442;
  assign n86488 = n77036 & ~n86442;
  assign n86489 = n77040 & ~n86442;
  assign n86490 = P2_P1_INSTADDRPOINTER_REG_9_ & n86410;
  assign n86491 = ~P2_P1_INSTADDRPOINTER_REG_10_ & n86490;
  assign n86492 = P2_P1_INSTADDRPOINTER_REG_10_ & ~n86490;
  assign n86493 = ~n86491 & ~n86492;
  assign n86494 = n77056 & ~n86493;
  assign n86495 = n77048 & ~n86493;
  assign n86496 = ~n86487 & ~n86488;
  assign n86497 = ~n86489 & n86496;
  assign n86498 = ~n86494 & n86497;
  assign n86499 = ~n86495 & n86498;
  assign n86500 = ~P2_P1_INSTADDRPOINTER_REG_10_ & ~n86425;
  assign n86501 = ~n86423 & n86475;
  assign n86502 = ~n86500 & ~n86501;
  assign n86503 = n77059 & n86502;
  assign n86504 = n86486 & n86499;
  assign n86505 = ~n86503 & n86504;
  assign n86506 = n86455 & ~n86456;
  assign n86507 = ~n86470 & n86506;
  assign n86508 = n86479 & n86507;
  assign n86509 = n86505 & n86508;
  assign n86510 = n85257 & ~n86509;
  assign n86511 = ~n86437 & ~n86438;
  assign n15581 = n86510 | ~n86511;
  assign n86513 = P2_P1_INSTADDRPOINTER_REG_11_ & n85256;
  assign n86514 = P2_P1_REIP_REG_11_ & n85401;
  assign n86515 = ~n86513 & ~n86514;
  assign n86516 = P2_P1_INSTADDRPOINTER_REG_10_ & n86445;
  assign n86517 = ~P2_P1_INSTADDRPOINTER_REG_11_ & n86516;
  assign n86518 = P2_P1_INSTADDRPOINTER_REG_11_ & ~n86516;
  assign n86519 = ~n86517 & ~n86518;
  assign n86520 = n85381 & ~n86519;
  assign n86521 = n77102 & ~n86519;
  assign n86522 = n85370 & ~n86519;
  assign n86523 = n85374 & ~n86519;
  assign n86524 = ~n86520 & ~n86521;
  assign n86525 = ~n86522 & n86524;
  assign n86526 = ~n86523 & n86525;
  assign n86527 = P2_P1_INSTADDRPOINTER_REG_10_ & n86439;
  assign n86528 = ~P2_P1_INSTADDRPOINTER_REG_11_ & n86527;
  assign n86529 = P2_P1_INSTADDRPOINTER_REG_11_ & ~n86527;
  assign n86530 = ~n86528 & ~n86529;
  assign n86531 = n76958 & ~n86530;
  assign n86532 = n77036 & ~n86530;
  assign n86533 = n77040 & ~n86530;
  assign n86534 = P2_P1_INSTADDRPOINTER_REG_10_ & n86490;
  assign n86535 = ~P2_P1_INSTADDRPOINTER_REG_11_ & n86534;
  assign n86536 = P2_P1_INSTADDRPOINTER_REG_11_ & ~n86534;
  assign n86537 = ~n86535 & ~n86536;
  assign n86538 = n77056 & ~n86537;
  assign n86539 = n77048 & ~n86537;
  assign n86540 = ~n86531 & ~n86532;
  assign n86541 = ~n86533 & n86540;
  assign n86542 = ~n86538 & n86541;
  assign n86543 = ~n86539 & n86542;
  assign n86544 = P2_P1_INSTADDRPOINTER_REG_11_ & ~n86501;
  assign n86545 = ~P2_P1_INSTADDRPOINTER_REG_11_ & n86501;
  assign n86546 = ~n86544 & ~n86545;
  assign n86547 = n77059 & ~n86546;
  assign n86548 = n86526 & n86543;
  assign n86549 = ~n86547 & n86548;
  assign n86550 = n77255 & ~n86519;
  assign n86551 = n77098 & ~n86519;
  assign n86552 = ~n86550 & ~n86551;
  assign n86553 = ~n77145 & ~n86519;
  assign n86554 = n86459 & ~n86465;
  assign n86555 = n86457 & ~n86466;
  assign n86556 = ~n86287 & n86555;
  assign n86557 = n86554 & ~n86556;
  assign n86558 = ~P2_P1_INSTADDRPOINTER_REG_11_ & ~n86192;
  assign n86559 = P2_P1_INSTADDRPOINTER_REG_11_ & n86192;
  assign n86560 = ~n86558 & ~n86559;
  assign n86561 = n86557 & ~n86560;
  assign n86562 = ~n86557 & n86560;
  assign n86563 = ~n86561 & ~n86562;
  assign n86564 = n85362 & ~n86563;
  assign n86565 = n77216 & ~n86530;
  assign n86566 = n77217 & ~n86530;
  assign n86567 = n85265 & ~n86519;
  assign n86568 = n77032 & ~n86530;
  assign n86569 = n85268 & ~n86519;
  assign n86570 = ~n86568 & ~n86569;
  assign n86571 = ~n86565 & ~n86566;
  assign n86572 = ~n86567 & n86571;
  assign n86573 = n86570 & n86572;
  assign n86574 = P2_P1_INSTADDRPOINTER_REG_11_ & ~n86476;
  assign n86575 = ~P2_P1_INSTADDRPOINTER_REG_11_ & n86476;
  assign n86576 = ~n86574 & ~n86575;
  assign n86577 = n85364 & ~n86576;
  assign n86578 = n86552 & ~n86553;
  assign n86579 = ~n86564 & n86578;
  assign n86580 = n86573 & n86579;
  assign n86581 = ~n86577 & n86580;
  assign n86582 = n86549 & n86581;
  assign n86583 = n85257 & ~n86582;
  assign n15586 = ~n86515 | n86583;
  assign n86585 = P2_P1_INSTADDRPOINTER_REG_12_ & n85256;
  assign n86586 = P2_P1_REIP_REG_12_ & n85401;
  assign n86587 = P2_P1_INSTADDRPOINTER_REG_11_ & n86527;
  assign n86588 = ~P2_P1_INSTADDRPOINTER_REG_12_ & n86587;
  assign n86589 = P2_P1_INSTADDRPOINTER_REG_12_ & ~n86587;
  assign n86590 = ~n86588 & ~n86589;
  assign n86591 = n77216 & ~n86590;
  assign n86592 = n77217 & ~n86590;
  assign n86593 = P2_P1_INSTADDRPOINTER_REG_11_ & n86516;
  assign n86594 = ~P2_P1_INSTADDRPOINTER_REG_12_ & n86593;
  assign n86595 = P2_P1_INSTADDRPOINTER_REG_12_ & ~n86593;
  assign n86596 = ~n86594 & ~n86595;
  assign n86597 = n85265 & ~n86596;
  assign n86598 = n77032 & ~n86590;
  assign n86599 = n85268 & ~n86596;
  assign n86600 = ~n86598 & ~n86599;
  assign n86601 = ~n86591 & ~n86592;
  assign n86602 = ~n86597 & n86601;
  assign n86603 = n86600 & n86602;
  assign n86604 = ~n77145 & ~n86596;
  assign n86605 = ~P2_P1_INSTADDRPOINTER_REG_12_ & ~n86192;
  assign n86606 = P2_P1_INSTADDRPOINTER_REG_12_ & n86192;
  assign n86607 = ~n86605 & ~n86606;
  assign n86608 = P2_P1_INSTADDRPOINTER_REG_11_ & ~n86192;
  assign n86609 = ~P2_P1_INSTADDRPOINTER_REG_11_ & n86192;
  assign n86610 = ~n86557 & ~n86609;
  assign n86611 = ~n86608 & ~n86610;
  assign n86612 = ~n86607 & n86611;
  assign n86613 = ~P2_P1_INSTADDRPOINTER_REG_12_ & n86192;
  assign n86614 = P2_P1_INSTADDRPOINTER_REG_12_ & ~n86192;
  assign n86615 = ~n86613 & ~n86614;
  assign n86616 = ~n86611 & ~n86615;
  assign n86617 = ~n86612 & ~n86616;
  assign n86618 = n85362 & ~n86617;
  assign n86619 = n77255 & ~n86596;
  assign n86620 = n77098 & ~n86596;
  assign n86621 = ~n86619 & ~n86620;
  assign n86622 = P2_P1_INSTADDRPOINTER_REG_11_ & n86476;
  assign n86623 = ~P2_P1_INSTADDRPOINTER_REG_12_ & ~n86622;
  assign n86624 = P2_P1_INSTADDRPOINTER_REG_11_ & P2_P1_INSTADDRPOINTER_REG_12_;
  assign n86625 = n86476 & n86624;
  assign n86626 = ~n86623 & ~n86625;
  assign n86627 = n85364 & n86626;
  assign n86628 = n86621 & ~n86627;
  assign n86629 = n85381 & ~n86596;
  assign n86630 = n77102 & ~n86596;
  assign n86631 = n85370 & ~n86596;
  assign n86632 = n85374 & ~n86596;
  assign n86633 = ~n86629 & ~n86630;
  assign n86634 = ~n86631 & n86633;
  assign n86635 = ~n86632 & n86634;
  assign n86636 = n76958 & ~n86590;
  assign n86637 = n77036 & ~n86590;
  assign n86638 = n77040 & ~n86590;
  assign n86639 = P2_P1_INSTADDRPOINTER_REG_11_ & n86534;
  assign n86640 = ~P2_P1_INSTADDRPOINTER_REG_12_ & n86639;
  assign n86641 = P2_P1_INSTADDRPOINTER_REG_12_ & ~n86639;
  assign n86642 = ~n86640 & ~n86641;
  assign n86643 = n77056 & ~n86642;
  assign n86644 = n77048 & ~n86642;
  assign n86645 = ~n86636 & ~n86637;
  assign n86646 = ~n86638 & n86645;
  assign n86647 = ~n86643 & n86646;
  assign n86648 = ~n86644 & n86647;
  assign n86649 = P2_P1_INSTADDRPOINTER_REG_11_ & n86501;
  assign n86650 = ~P2_P1_INSTADDRPOINTER_REG_12_ & ~n86649;
  assign n86651 = n86501 & n86624;
  assign n86652 = ~n86650 & ~n86651;
  assign n86653 = n77059 & n86652;
  assign n86654 = n86635 & n86648;
  assign n86655 = ~n86653 & n86654;
  assign n86656 = n86603 & ~n86604;
  assign n86657 = ~n86618 & n86656;
  assign n86658 = n86628 & n86657;
  assign n86659 = n86655 & n86658;
  assign n86660 = n85257 & ~n86659;
  assign n86661 = ~n86585 & ~n86586;
  assign n15591 = n86660 | ~n86661;
  assign n86663 = P2_P1_INSTADDRPOINTER_REG_13_ & n85256;
  assign n86664 = P2_P1_REIP_REG_13_ & n85401;
  assign n86665 = P2_P1_INSTADDRPOINTER_REG_12_ & n86587;
  assign n86666 = ~P2_P1_INSTADDRPOINTER_REG_13_ & n86665;
  assign n86667 = P2_P1_INSTADDRPOINTER_REG_13_ & ~n86665;
  assign n86668 = ~n86666 & ~n86667;
  assign n86669 = n77216 & ~n86668;
  assign n86670 = n77217 & ~n86668;
  assign n86671 = P2_P1_INSTADDRPOINTER_REG_12_ & n86593;
  assign n86672 = ~P2_P1_INSTADDRPOINTER_REG_13_ & n86671;
  assign n86673 = P2_P1_INSTADDRPOINTER_REG_13_ & ~n86671;
  assign n86674 = ~n86672 & ~n86673;
  assign n86675 = n85265 & ~n86674;
  assign n86676 = n77032 & ~n86668;
  assign n86677 = n85268 & ~n86674;
  assign n86678 = ~n86676 & ~n86677;
  assign n86679 = ~n86669 & ~n86670;
  assign n86680 = ~n86675 & n86679;
  assign n86681 = n86678 & n86680;
  assign n86682 = ~n77145 & ~n86674;
  assign n86683 = P2_P1_INSTADDRPOINTER_REG_13_ & ~n86192;
  assign n86684 = P2_P1_INSTADDRPOINTER_REG_12_ & P2_P1_INSTADDRPOINTER_REG_13_;
  assign n86685 = n86192 & ~n86684;
  assign n86686 = ~n86683 & ~n86685;
  assign n86687 = n86611 & ~n86614;
  assign n86688 = n86686 & ~n86687;
  assign n86689 = ~P2_P1_INSTADDRPOINTER_REG_13_ & ~n86192;
  assign n86690 = P2_P1_INSTADDRPOINTER_REG_13_ & n86192;
  assign n86691 = ~n86689 & ~n86690;
  assign n86692 = ~n86614 & n86691;
  assign n86693 = ~n86611 & ~n86613;
  assign n86694 = n86692 & ~n86693;
  assign n86695 = ~n86688 & ~n86694;
  assign n86696 = n85362 & n86695;
  assign n86697 = n77255 & ~n86674;
  assign n86698 = n77098 & ~n86674;
  assign n86699 = ~n86697 & ~n86698;
  assign n86700 = ~P2_P1_INSTADDRPOINTER_REG_13_ & ~n86625;
  assign n86701 = P2_P1_INSTADDRPOINTER_REG_13_ & n86625;
  assign n86702 = ~n86700 & ~n86701;
  assign n86703 = n85364 & n86702;
  assign n86704 = n86699 & ~n86703;
  assign n86705 = n85381 & ~n86674;
  assign n86706 = n77102 & ~n86674;
  assign n86707 = n85370 & ~n86674;
  assign n86708 = n85374 & ~n86674;
  assign n86709 = ~n86705 & ~n86706;
  assign n86710 = ~n86707 & n86709;
  assign n86711 = ~n86708 & n86710;
  assign n86712 = n76958 & ~n86668;
  assign n86713 = n77036 & ~n86668;
  assign n86714 = n77040 & ~n86668;
  assign n86715 = P2_P1_INSTADDRPOINTER_REG_12_ & n86639;
  assign n86716 = ~P2_P1_INSTADDRPOINTER_REG_13_ & n86715;
  assign n86717 = P2_P1_INSTADDRPOINTER_REG_13_ & ~n86715;
  assign n86718 = ~n86716 & ~n86717;
  assign n86719 = n77056 & ~n86718;
  assign n86720 = n77048 & ~n86718;
  assign n86721 = ~n86712 & ~n86713;
  assign n86722 = ~n86714 & n86721;
  assign n86723 = ~n86719 & n86722;
  assign n86724 = ~n86720 & n86723;
  assign n86725 = ~P2_P1_INSTADDRPOINTER_REG_13_ & ~n86651;
  assign n86726 = P2_P1_INSTADDRPOINTER_REG_13_ & n86651;
  assign n86727 = ~n86725 & ~n86726;
  assign n86728 = n77059 & n86727;
  assign n86729 = n86711 & n86724;
  assign n86730 = ~n86728 & n86729;
  assign n86731 = n86681 & ~n86682;
  assign n86732 = ~n86696 & n86731;
  assign n86733 = n86704 & n86732;
  assign n86734 = n86730 & n86733;
  assign n86735 = n85257 & ~n86734;
  assign n86736 = ~n86663 & ~n86664;
  assign n15596 = n86735 | ~n86736;
  assign n86738 = P2_P1_INSTADDRPOINTER_REG_14_ & n85256;
  assign n86739 = P2_P1_REIP_REG_14_ & n85401;
  assign n86740 = ~n86738 & ~n86739;
  assign n86741 = P2_P1_INSTADDRPOINTER_REG_13_ & n86671;
  assign n86742 = ~P2_P1_INSTADDRPOINTER_REG_14_ & n86741;
  assign n86743 = P2_P1_INSTADDRPOINTER_REG_14_ & ~n86741;
  assign n86744 = ~n86742 & ~n86743;
  assign n86745 = n85381 & ~n86744;
  assign n86746 = n77102 & ~n86744;
  assign n86747 = n85370 & ~n86744;
  assign n86748 = n85374 & ~n86744;
  assign n86749 = ~n86745 & ~n86746;
  assign n86750 = ~n86747 & n86749;
  assign n86751 = ~n86748 & n86750;
  assign n86752 = P2_P1_INSTADDRPOINTER_REG_13_ & n86665;
  assign n86753 = ~P2_P1_INSTADDRPOINTER_REG_14_ & n86752;
  assign n86754 = P2_P1_INSTADDRPOINTER_REG_14_ & ~n86752;
  assign n86755 = ~n86753 & ~n86754;
  assign n86756 = n76958 & ~n86755;
  assign n86757 = n77036 & ~n86755;
  assign n86758 = n77040 & ~n86755;
  assign n86759 = P2_P1_INSTADDRPOINTER_REG_13_ & n86715;
  assign n86760 = ~P2_P1_INSTADDRPOINTER_REG_14_ & n86759;
  assign n86761 = P2_P1_INSTADDRPOINTER_REG_14_ & ~n86759;
  assign n86762 = ~n86760 & ~n86761;
  assign n86763 = n77056 & ~n86762;
  assign n86764 = n77048 & ~n86762;
  assign n86765 = ~n86756 & ~n86757;
  assign n86766 = ~n86758 & n86765;
  assign n86767 = ~n86763 & n86766;
  assign n86768 = ~n86764 & n86767;
  assign n86769 = ~P2_P1_INSTADDRPOINTER_REG_14_ & n86726;
  assign n86770 = P2_P1_INSTADDRPOINTER_REG_14_ & ~n86726;
  assign n86771 = ~n86769 & ~n86770;
  assign n86772 = n77059 & ~n86771;
  assign n86773 = n86751 & n86768;
  assign n86774 = ~n86772 & n86773;
  assign n86775 = n77255 & ~n86744;
  assign n86776 = n77098 & ~n86744;
  assign n86777 = ~n86775 & ~n86776;
  assign n86778 = ~n77145 & ~n86744;
  assign n86779 = n77216 & ~n86755;
  assign n86780 = n77217 & ~n86755;
  assign n86781 = n85265 & ~n86744;
  assign n86782 = n77032 & ~n86755;
  assign n86783 = n85268 & ~n86744;
  assign n86784 = ~n86782 & ~n86783;
  assign n86785 = ~n86779 & ~n86780;
  assign n86786 = ~n86781 & n86785;
  assign n86787 = n86784 & n86786;
  assign n86788 = ~n86614 & ~n86683;
  assign n86789 = ~n86608 & n86788;
  assign n86790 = ~n86609 & ~n86685;
  assign n86791 = ~n86557 & n86790;
  assign n86792 = n86789 & ~n86791;
  assign n86793 = ~P2_P1_INSTADDRPOINTER_REG_14_ & ~n86192;
  assign n86794 = P2_P1_INSTADDRPOINTER_REG_14_ & n86192;
  assign n86795 = ~n86793 & ~n86794;
  assign n86796 = n86792 & ~n86795;
  assign n86797 = ~n86792 & n86795;
  assign n86798 = ~n86796 & ~n86797;
  assign n86799 = n85362 & ~n86798;
  assign n86800 = ~P2_P1_INSTADDRPOINTER_REG_14_ & n86701;
  assign n86801 = P2_P1_INSTADDRPOINTER_REG_14_ & ~n86701;
  assign n86802 = ~n86800 & ~n86801;
  assign n86803 = n85364 & ~n86802;
  assign n86804 = n86777 & ~n86778;
  assign n86805 = n86787 & n86804;
  assign n86806 = ~n86799 & n86805;
  assign n86807 = ~n86803 & n86806;
  assign n86808 = n86774 & n86807;
  assign n86809 = n85257 & ~n86808;
  assign n15601 = ~n86740 | n86809;
  assign n86811 = P2_P1_INSTADDRPOINTER_REG_15_ & n85256;
  assign n86812 = P2_P1_REIP_REG_15_ & n85401;
  assign n86813 = ~n86811 & ~n86812;
  assign n86814 = P2_P1_INSTADDRPOINTER_REG_14_ & n86741;
  assign n86815 = ~P2_P1_INSTADDRPOINTER_REG_15_ & n86814;
  assign n86816 = P2_P1_INSTADDRPOINTER_REG_15_ & ~n86814;
  assign n86817 = ~n86815 & ~n86816;
  assign n86818 = n85381 & ~n86817;
  assign n86819 = n77102 & ~n86817;
  assign n86820 = n85370 & ~n86817;
  assign n86821 = n85374 & ~n86817;
  assign n86822 = ~n86818 & ~n86819;
  assign n86823 = ~n86820 & n86822;
  assign n86824 = ~n86821 & n86823;
  assign n86825 = P2_P1_INSTADDRPOINTER_REG_14_ & n86752;
  assign n86826 = ~P2_P1_INSTADDRPOINTER_REG_15_ & n86825;
  assign n86827 = P2_P1_INSTADDRPOINTER_REG_15_ & ~n86825;
  assign n86828 = ~n86826 & ~n86827;
  assign n86829 = n76958 & ~n86828;
  assign n86830 = n77036 & ~n86828;
  assign n86831 = n77040 & ~n86828;
  assign n86832 = P2_P1_INSTADDRPOINTER_REG_14_ & n86759;
  assign n86833 = ~P2_P1_INSTADDRPOINTER_REG_15_ & n86832;
  assign n86834 = P2_P1_INSTADDRPOINTER_REG_15_ & ~n86832;
  assign n86835 = ~n86833 & ~n86834;
  assign n86836 = n77056 & ~n86835;
  assign n86837 = n77048 & ~n86835;
  assign n86838 = ~n86829 & ~n86830;
  assign n86839 = ~n86831 & n86838;
  assign n86840 = ~n86836 & n86839;
  assign n86841 = ~n86837 & n86840;
  assign n86842 = P2_P1_INSTADDRPOINTER_REG_14_ & n86726;
  assign n86843 = ~P2_P1_INSTADDRPOINTER_REG_15_ & ~n86842;
  assign n86844 = P2_P1_INSTADDRPOINTER_REG_14_ & P2_P1_INSTADDRPOINTER_REG_15_;
  assign n86845 = P2_P1_INSTADDRPOINTER_REG_13_ & n86844;
  assign n86846 = n86651 & n86845;
  assign n86847 = ~n86843 & ~n86846;
  assign n86848 = n77059 & n86847;
  assign n86849 = n86824 & n86841;
  assign n86850 = ~n86848 & n86849;
  assign n86851 = n77255 & ~n86817;
  assign n86852 = n77098 & ~n86817;
  assign n86853 = ~n86851 & ~n86852;
  assign n86854 = ~n77145 & ~n86817;
  assign n86855 = n77216 & ~n86828;
  assign n86856 = n77217 & ~n86828;
  assign n86857 = n85265 & ~n86817;
  assign n86858 = n77032 & ~n86828;
  assign n86859 = n85268 & ~n86817;
  assign n86860 = ~n86858 & ~n86859;
  assign n86861 = ~n86855 & ~n86856;
  assign n86862 = ~n86857 & n86861;
  assign n86863 = n86860 & n86862;
  assign n86864 = P2_P1_INSTADDRPOINTER_REG_14_ & ~n86192;
  assign n86865 = n86789 & ~n86864;
  assign n86866 = ~P2_P1_INSTADDRPOINTER_REG_14_ & n86192;
  assign n86867 = n86790 & ~n86866;
  assign n86868 = ~n86557 & n86867;
  assign n86869 = n86865 & ~n86868;
  assign n86870 = ~P2_P1_INSTADDRPOINTER_REG_15_ & ~n86192;
  assign n86871 = P2_P1_INSTADDRPOINTER_REG_15_ & n86192;
  assign n86872 = ~n86870 & ~n86871;
  assign n86873 = n86869 & ~n86872;
  assign n86874 = ~n86869 & n86872;
  assign n86875 = ~n86873 & ~n86874;
  assign n86876 = n85362 & ~n86875;
  assign n86877 = P2_P1_INSTADDRPOINTER_REG_14_ & n86701;
  assign n86878 = ~P2_P1_INSTADDRPOINTER_REG_15_ & ~n86877;
  assign n86879 = n86625 & n86845;
  assign n86880 = ~n86878 & ~n86879;
  assign n86881 = n85364 & n86880;
  assign n86882 = n86853 & ~n86854;
  assign n86883 = n86863 & n86882;
  assign n86884 = ~n86876 & n86883;
  assign n86885 = ~n86881 & n86884;
  assign n86886 = n86850 & n86885;
  assign n86887 = n85257 & ~n86886;
  assign n15606 = ~n86813 | n86887;
  assign n86889 = P2_P1_INSTADDRPOINTER_REG_16_ & n85256;
  assign n86890 = P2_P1_REIP_REG_16_ & n85401;
  assign n86891 = ~n86889 & ~n86890;
  assign n86892 = P2_P1_INSTADDRPOINTER_REG_15_ & n86814;
  assign n86893 = ~P2_P1_INSTADDRPOINTER_REG_16_ & n86892;
  assign n86894 = P2_P1_INSTADDRPOINTER_REG_16_ & ~n86892;
  assign n86895 = ~n86893 & ~n86894;
  assign n86896 = n85381 & ~n86895;
  assign n86897 = n77102 & ~n86895;
  assign n86898 = n85370 & ~n86895;
  assign n86899 = n85374 & ~n86895;
  assign n86900 = ~n86896 & ~n86897;
  assign n86901 = ~n86898 & n86900;
  assign n86902 = ~n86899 & n86901;
  assign n86903 = P2_P1_INSTADDRPOINTER_REG_15_ & n86825;
  assign n86904 = ~P2_P1_INSTADDRPOINTER_REG_16_ & n86903;
  assign n86905 = P2_P1_INSTADDRPOINTER_REG_16_ & ~n86903;
  assign n86906 = ~n86904 & ~n86905;
  assign n86907 = n76958 & ~n86906;
  assign n86908 = n77036 & ~n86906;
  assign n86909 = n77040 & ~n86906;
  assign n86910 = P2_P1_INSTADDRPOINTER_REG_15_ & n86832;
  assign n86911 = ~P2_P1_INSTADDRPOINTER_REG_16_ & n86910;
  assign n86912 = P2_P1_INSTADDRPOINTER_REG_16_ & ~n86910;
  assign n86913 = ~n86911 & ~n86912;
  assign n86914 = n77056 & ~n86913;
  assign n86915 = n77048 & ~n86913;
  assign n86916 = ~n86907 & ~n86908;
  assign n86917 = ~n86909 & n86916;
  assign n86918 = ~n86914 & n86917;
  assign n86919 = ~n86915 & n86918;
  assign n86920 = ~P2_P1_INSTADDRPOINTER_REG_16_ & n86846;
  assign n86921 = P2_P1_INSTADDRPOINTER_REG_16_ & ~n86846;
  assign n86922 = ~n86920 & ~n86921;
  assign n86923 = n77059 & ~n86922;
  assign n86924 = n86902 & n86919;
  assign n86925 = ~n86923 & n86924;
  assign n86926 = n77255 & ~n86895;
  assign n86927 = n77098 & ~n86895;
  assign n86928 = ~n86926 & ~n86927;
  assign n86929 = ~n77145 & ~n86895;
  assign n86930 = P2_P1_INSTADDRPOINTER_REG_15_ & ~n86192;
  assign n86931 = ~P2_P1_INSTADDRPOINTER_REG_15_ & n86192;
  assign n86932 = ~n86869 & ~n86931;
  assign n86933 = ~n86930 & ~n86932;
  assign n86934 = ~P2_P1_INSTADDRPOINTER_REG_16_ & ~n86192;
  assign n86935 = P2_P1_INSTADDRPOINTER_REG_16_ & n86192;
  assign n86936 = ~n86934 & ~n86935;
  assign n86937 = n86933 & ~n86936;
  assign n86938 = ~n86933 & n86936;
  assign n86939 = ~n86937 & ~n86938;
  assign n86940 = n85362 & ~n86939;
  assign n86941 = n77216 & ~n86906;
  assign n86942 = n77217 & ~n86906;
  assign n86943 = n85265 & ~n86895;
  assign n86944 = n77032 & ~n86906;
  assign n86945 = n85268 & ~n86895;
  assign n86946 = ~n86944 & ~n86945;
  assign n86947 = ~n86941 & ~n86942;
  assign n86948 = ~n86943 & n86947;
  assign n86949 = n86946 & n86948;
  assign n86950 = ~P2_P1_INSTADDRPOINTER_REG_16_ & n86879;
  assign n86951 = P2_P1_INSTADDRPOINTER_REG_16_ & ~n86879;
  assign n86952 = ~n86950 & ~n86951;
  assign n86953 = n85364 & ~n86952;
  assign n86954 = n86928 & ~n86929;
  assign n86955 = ~n86940 & n86954;
  assign n86956 = n86949 & n86955;
  assign n86957 = ~n86953 & n86956;
  assign n86958 = n86925 & n86957;
  assign n86959 = n85257 & ~n86958;
  assign n15611 = ~n86891 | n86959;
  assign n86961 = P2_P1_INSTADDRPOINTER_REG_17_ & n85256;
  assign n86962 = P2_P1_REIP_REG_17_ & n85401;
  assign n86963 = P2_P1_INSTADDRPOINTER_REG_16_ & n86903;
  assign n86964 = ~P2_P1_INSTADDRPOINTER_REG_17_ & n86963;
  assign n86965 = P2_P1_INSTADDRPOINTER_REG_17_ & ~n86963;
  assign n86966 = ~n86964 & ~n86965;
  assign n86967 = n77216 & ~n86966;
  assign n86968 = n77217 & ~n86966;
  assign n86969 = P2_P1_INSTADDRPOINTER_REG_16_ & n86892;
  assign n86970 = ~P2_P1_INSTADDRPOINTER_REG_17_ & n86969;
  assign n86971 = P2_P1_INSTADDRPOINTER_REG_17_ & ~n86969;
  assign n86972 = ~n86970 & ~n86971;
  assign n86973 = n85265 & ~n86972;
  assign n86974 = n77032 & ~n86966;
  assign n86975 = n85268 & ~n86972;
  assign n86976 = ~n86974 & ~n86975;
  assign n86977 = ~n86967 & ~n86968;
  assign n86978 = ~n86973 & n86977;
  assign n86979 = n86976 & n86978;
  assign n86980 = ~n77145 & ~n86972;
  assign n86981 = P2_P1_INSTADDRPOINTER_REG_16_ & P2_P1_INSTADDRPOINTER_REG_17_;
  assign n86982 = ~n86933 & n86981;
  assign n86983 = n86192 & ~n86982;
  assign n86984 = P2_P1_INSTADDRPOINTER_REG_17_ & ~n86192;
  assign n86985 = ~P2_P1_INSTADDRPOINTER_REG_16_ & ~n86930;
  assign n86986 = ~n86932 & n86985;
  assign n86987 = ~n86983 & ~n86984;
  assign n86988 = ~n86986 & n86987;
  assign n86989 = P2_P1_INSTADDRPOINTER_REG_17_ & n86986;
  assign n86990 = ~n86192 & ~n86989;
  assign n86991 = P2_P1_INSTADDRPOINTER_REG_17_ & n86192;
  assign n86992 = P2_P1_INSTADDRPOINTER_REG_16_ & ~n86933;
  assign n86993 = ~n86990 & ~n86991;
  assign n86994 = ~n86992 & n86993;
  assign n86995 = ~n86988 & ~n86994;
  assign n86996 = n85362 & n86995;
  assign n86997 = n77255 & ~n86972;
  assign n86998 = n77098 & ~n86972;
  assign n86999 = ~n86997 & ~n86998;
  assign n87000 = P2_P1_INSTADDRPOINTER_REG_16_ & n86879;
  assign n87001 = ~P2_P1_INSTADDRPOINTER_REG_17_ & ~n87000;
  assign n87002 = n86879 & n86981;
  assign n87003 = ~n87001 & ~n87002;
  assign n87004 = n85364 & n87003;
  assign n87005 = n86999 & ~n87004;
  assign n87006 = n85381 & ~n86972;
  assign n87007 = n77102 & ~n86972;
  assign n87008 = n85370 & ~n86972;
  assign n87009 = n85374 & ~n86972;
  assign n87010 = ~n87006 & ~n87007;
  assign n87011 = ~n87008 & n87010;
  assign n87012 = ~n87009 & n87011;
  assign n87013 = n76958 & ~n86966;
  assign n87014 = n77036 & ~n86966;
  assign n87015 = n77040 & ~n86966;
  assign n87016 = P2_P1_INSTADDRPOINTER_REG_16_ & n86910;
  assign n87017 = ~P2_P1_INSTADDRPOINTER_REG_17_ & n87016;
  assign n87018 = P2_P1_INSTADDRPOINTER_REG_17_ & ~n87016;
  assign n87019 = ~n87017 & ~n87018;
  assign n87020 = n77056 & ~n87019;
  assign n87021 = n77048 & ~n87019;
  assign n87022 = ~n87013 & ~n87014;
  assign n87023 = ~n87015 & n87022;
  assign n87024 = ~n87020 & n87023;
  assign n87025 = ~n87021 & n87024;
  assign n87026 = P2_P1_INSTADDRPOINTER_REG_16_ & n86846;
  assign n87027 = ~P2_P1_INSTADDRPOINTER_REG_17_ & ~n87026;
  assign n87028 = n86846 & n86981;
  assign n87029 = ~n87027 & ~n87028;
  assign n87030 = n77059 & n87029;
  assign n87031 = n87012 & n87025;
  assign n87032 = ~n87030 & n87031;
  assign n87033 = n86979 & ~n86980;
  assign n87034 = ~n86996 & n87033;
  assign n87035 = n87005 & n87034;
  assign n87036 = n87032 & n87035;
  assign n87037 = n85257 & ~n87036;
  assign n87038 = ~n86961 & ~n86962;
  assign n15616 = n87037 | ~n87038;
  assign n87040 = P2_P1_INSTADDRPOINTER_REG_18_ & n85256;
  assign n87041 = P2_P1_REIP_REG_18_ & n85401;
  assign n87042 = ~n87040 & ~n87041;
  assign n87043 = P2_P1_INSTADDRPOINTER_REG_17_ & n86969;
  assign n87044 = ~P2_P1_INSTADDRPOINTER_REG_18_ & n87043;
  assign n87045 = P2_P1_INSTADDRPOINTER_REG_18_ & ~n87043;
  assign n87046 = ~n87044 & ~n87045;
  assign n87047 = n85381 & ~n87046;
  assign n87048 = n77102 & ~n87046;
  assign n87049 = n85370 & ~n87046;
  assign n87050 = n85374 & ~n87046;
  assign n87051 = ~n87047 & ~n87048;
  assign n87052 = ~n87049 & n87051;
  assign n87053 = ~n87050 & n87052;
  assign n87054 = P2_P1_INSTADDRPOINTER_REG_17_ & n86963;
  assign n87055 = ~P2_P1_INSTADDRPOINTER_REG_18_ & n87054;
  assign n87056 = P2_P1_INSTADDRPOINTER_REG_18_ & ~n87054;
  assign n87057 = ~n87055 & ~n87056;
  assign n87058 = n76958 & ~n87057;
  assign n87059 = n77036 & ~n87057;
  assign n87060 = n77040 & ~n87057;
  assign n87061 = P2_P1_INSTADDRPOINTER_REG_17_ & n87016;
  assign n87062 = ~P2_P1_INSTADDRPOINTER_REG_18_ & n87061;
  assign n87063 = P2_P1_INSTADDRPOINTER_REG_18_ & ~n87061;
  assign n87064 = ~n87062 & ~n87063;
  assign n87065 = n77056 & ~n87064;
  assign n87066 = n77048 & ~n87064;
  assign n87067 = ~n87058 & ~n87059;
  assign n87068 = ~n87060 & n87067;
  assign n87069 = ~n87065 & n87068;
  assign n87070 = ~n87066 & n87069;
  assign n87071 = ~P2_P1_INSTADDRPOINTER_REG_18_ & n87028;
  assign n87072 = P2_P1_INSTADDRPOINTER_REG_18_ & ~n87028;
  assign n87073 = ~n87071 & ~n87072;
  assign n87074 = n77059 & ~n87073;
  assign n87075 = n87053 & n87070;
  assign n87076 = ~n87074 & n87075;
  assign n87077 = n77255 & ~n87046;
  assign n87078 = n77098 & ~n87046;
  assign n87079 = ~n87077 & ~n87078;
  assign n87080 = ~n77145 & ~n87046;
  assign n87081 = ~n86192 & ~n86986;
  assign n87082 = ~n86982 & ~n87081;
  assign n87083 = ~n86984 & n87082;
  assign n87084 = ~P2_P1_INSTADDRPOINTER_REG_18_ & ~n86192;
  assign n87085 = P2_P1_INSTADDRPOINTER_REG_18_ & n86192;
  assign n87086 = ~n87084 & ~n87085;
  assign n87087 = n87083 & ~n87086;
  assign n87088 = ~n87083 & n87086;
  assign n87089 = ~n87087 & ~n87088;
  assign n87090 = n85362 & ~n87089;
  assign n87091 = n77216 & ~n87057;
  assign n87092 = n77217 & ~n87057;
  assign n87093 = n85265 & ~n87046;
  assign n87094 = n77032 & ~n87057;
  assign n87095 = n85268 & ~n87046;
  assign n87096 = ~n87094 & ~n87095;
  assign n87097 = ~n87091 & ~n87092;
  assign n87098 = ~n87093 & n87097;
  assign n87099 = n87096 & n87098;
  assign n87100 = ~P2_P1_INSTADDRPOINTER_REG_18_ & n87002;
  assign n87101 = P2_P1_INSTADDRPOINTER_REG_18_ & ~n87002;
  assign n87102 = ~n87100 & ~n87101;
  assign n87103 = n85364 & ~n87102;
  assign n87104 = n87079 & ~n87080;
  assign n87105 = ~n87090 & n87104;
  assign n87106 = n87099 & n87105;
  assign n87107 = ~n87103 & n87106;
  assign n87108 = n87076 & n87107;
  assign n87109 = n85257 & ~n87108;
  assign n15621 = ~n87042 | n87109;
  assign n87111 = P2_P1_INSTADDRPOINTER_REG_19_ & n85256;
  assign n87112 = P2_P1_REIP_REG_19_ & n85401;
  assign n87113 = P2_P1_INSTADDRPOINTER_REG_18_ & n87054;
  assign n87114 = ~P2_P1_INSTADDRPOINTER_REG_19_ & n87113;
  assign n87115 = P2_P1_INSTADDRPOINTER_REG_19_ & ~n87113;
  assign n87116 = ~n87114 & ~n87115;
  assign n87117 = n77216 & ~n87116;
  assign n87118 = n77217 & ~n87116;
  assign n87119 = P2_P1_INSTADDRPOINTER_REG_18_ & n87043;
  assign n87120 = ~P2_P1_INSTADDRPOINTER_REG_19_ & n87119;
  assign n87121 = P2_P1_INSTADDRPOINTER_REG_19_ & ~n87119;
  assign n87122 = ~n87120 & ~n87121;
  assign n87123 = n85265 & ~n87122;
  assign n87124 = n77032 & ~n87116;
  assign n87125 = n85268 & ~n87122;
  assign n87126 = ~n87124 & ~n87125;
  assign n87127 = ~n87117 & ~n87118;
  assign n87128 = ~n87123 & n87127;
  assign n87129 = n87126 & n87128;
  assign n87130 = ~n77145 & ~n87122;
  assign n87131 = ~P2_P1_INSTADDRPOINTER_REG_19_ & ~n86192;
  assign n87132 = P2_P1_INSTADDRPOINTER_REG_19_ & n86192;
  assign n87133 = ~n87131 & ~n87132;
  assign n87134 = ~P2_P1_INSTADDRPOINTER_REG_18_ & n86192;
  assign n87135 = ~n87083 & ~n87134;
  assign n87136 = P2_P1_INSTADDRPOINTER_REG_18_ & ~n86192;
  assign n87137 = ~n87135 & ~n87136;
  assign n87138 = ~n87133 & n87137;
  assign n87139 = ~P2_P1_INSTADDRPOINTER_REG_19_ & n86192;
  assign n87140 = P2_P1_INSTADDRPOINTER_REG_19_ & ~n86192;
  assign n87141 = ~n87139 & ~n87140;
  assign n87142 = ~n87137 & ~n87141;
  assign n87143 = ~n87138 & ~n87142;
  assign n87144 = n85362 & ~n87143;
  assign n87145 = n77255 & ~n87122;
  assign n87146 = n77098 & ~n87122;
  assign n87147 = ~n87145 & ~n87146;
  assign n87148 = P2_P1_INSTADDRPOINTER_REG_18_ & n87002;
  assign n87149 = ~P2_P1_INSTADDRPOINTER_REG_19_ & ~n87148;
  assign n87150 = P2_P1_INSTADDRPOINTER_REG_18_ & P2_P1_INSTADDRPOINTER_REG_19_;
  assign n87151 = n87002 & n87150;
  assign n87152 = ~n87149 & ~n87151;
  assign n87153 = n85364 & n87152;
  assign n87154 = n87147 & ~n87153;
  assign n87155 = n85381 & ~n87122;
  assign n87156 = n77102 & ~n87122;
  assign n87157 = n85370 & ~n87122;
  assign n87158 = n85374 & ~n87122;
  assign n87159 = ~n87155 & ~n87156;
  assign n87160 = ~n87157 & n87159;
  assign n87161 = ~n87158 & n87160;
  assign n87162 = n76958 & ~n87116;
  assign n87163 = n77036 & ~n87116;
  assign n87164 = n77040 & ~n87116;
  assign n87165 = P2_P1_INSTADDRPOINTER_REG_18_ & n87061;
  assign n87166 = ~P2_P1_INSTADDRPOINTER_REG_19_ & n87165;
  assign n87167 = P2_P1_INSTADDRPOINTER_REG_19_ & ~n87165;
  assign n87168 = ~n87166 & ~n87167;
  assign n87169 = n77056 & ~n87168;
  assign n87170 = n77048 & ~n87168;
  assign n87171 = ~n87162 & ~n87163;
  assign n87172 = ~n87164 & n87171;
  assign n87173 = ~n87169 & n87172;
  assign n87174 = ~n87170 & n87173;
  assign n87175 = P2_P1_INSTADDRPOINTER_REG_18_ & n87028;
  assign n87176 = ~P2_P1_INSTADDRPOINTER_REG_19_ & ~n87175;
  assign n87177 = n87028 & n87150;
  assign n87178 = ~n87176 & ~n87177;
  assign n87179 = n77059 & n87178;
  assign n87180 = n87161 & n87174;
  assign n87181 = ~n87179 & n87180;
  assign n87182 = n87129 & ~n87130;
  assign n87183 = ~n87144 & n87182;
  assign n87184 = n87154 & n87183;
  assign n87185 = n87181 & n87184;
  assign n87186 = n85257 & ~n87185;
  assign n87187 = ~n87111 & ~n87112;
  assign n15626 = n87186 | ~n87187;
  assign n87189 = P2_P1_INSTADDRPOINTER_REG_20_ & n85256;
  assign n87190 = P2_P1_REIP_REG_20_ & n85401;
  assign n87191 = ~n87189 & ~n87190;
  assign n87192 = P2_P1_INSTADDRPOINTER_REG_19_ & P2_P1_INSTADDRPOINTER_REG_20_;
  assign n87193 = n86192 & ~n87192;
  assign n87194 = P2_P1_INSTADDRPOINTER_REG_20_ & ~n86192;
  assign n87195 = ~n87193 & ~n87194;
  assign n87196 = n87137 & ~n87140;
  assign n87197 = n87195 & ~n87196;
  assign n87198 = ~P2_P1_INSTADDRPOINTER_REG_19_ & n87137;
  assign n87199 = P2_P1_INSTADDRPOINTER_REG_20_ & n87198;
  assign n87200 = ~n86192 & ~n87199;
  assign n87201 = P2_P1_INSTADDRPOINTER_REG_20_ & n86192;
  assign n87202 = P2_P1_INSTADDRPOINTER_REG_19_ & ~n87137;
  assign n87203 = ~n87200 & ~n87201;
  assign n87204 = ~n87202 & n87203;
  assign n87205 = ~n87197 & ~n87204;
  assign n87206 = n85362 & n87205;
  assign n87207 = P2_P1_INSTADDRPOINTER_REG_19_ & n87119;
  assign n87208 = ~P2_P1_INSTADDRPOINTER_REG_20_ & n87207;
  assign n87209 = P2_P1_INSTADDRPOINTER_REG_20_ & ~n87207;
  assign n87210 = ~n87208 & ~n87209;
  assign n87211 = ~n77145 & ~n87210;
  assign n87212 = n77255 & ~n87210;
  assign n87213 = n77098 & ~n87210;
  assign n87214 = ~n87212 & ~n87213;
  assign n87215 = P2_P1_INSTADDRPOINTER_REG_19_ & n87113;
  assign n87216 = ~P2_P1_INSTADDRPOINTER_REG_20_ & n87215;
  assign n87217 = P2_P1_INSTADDRPOINTER_REG_20_ & ~n87215;
  assign n87218 = ~n87216 & ~n87217;
  assign n87219 = n77216 & ~n87218;
  assign n87220 = n77217 & ~n87218;
  assign n87221 = n85265 & ~n87210;
  assign n87222 = n77032 & ~n87218;
  assign n87223 = n85268 & ~n87210;
  assign n87224 = ~n87222 & ~n87223;
  assign n87225 = ~n87219 & ~n87220;
  assign n87226 = ~n87221 & n87225;
  assign n87227 = n87224 & n87226;
  assign n87228 = ~P2_P1_INSTADDRPOINTER_REG_20_ & ~n87151;
  assign n87229 = P2_P1_INSTADDRPOINTER_REG_20_ & n87151;
  assign n87230 = ~n87228 & ~n87229;
  assign n87231 = n85364 & n87230;
  assign n87232 = n85381 & ~n87210;
  assign n87233 = n77102 & ~n87210;
  assign n87234 = n85370 & ~n87210;
  assign n87235 = n85374 & ~n87210;
  assign n87236 = ~n87232 & ~n87233;
  assign n87237 = ~n87234 & n87236;
  assign n87238 = ~n87235 & n87237;
  assign n87239 = n76958 & ~n87218;
  assign n87240 = n77036 & ~n87218;
  assign n87241 = n77040 & ~n87218;
  assign n87242 = P2_P1_INSTADDRPOINTER_REG_19_ & n87165;
  assign n87243 = ~P2_P1_INSTADDRPOINTER_REG_20_ & n87242;
  assign n87244 = P2_P1_INSTADDRPOINTER_REG_20_ & ~n87242;
  assign n87245 = ~n87243 & ~n87244;
  assign n87246 = n77056 & ~n87245;
  assign n87247 = n77048 & ~n87245;
  assign n87248 = ~n87239 & ~n87240;
  assign n87249 = ~n87241 & n87248;
  assign n87250 = ~n87246 & n87249;
  assign n87251 = ~n87247 & n87250;
  assign n87252 = ~P2_P1_INSTADDRPOINTER_REG_20_ & ~n87177;
  assign n87253 = P2_P1_INSTADDRPOINTER_REG_20_ & n87177;
  assign n87254 = ~n87252 & ~n87253;
  assign n87255 = n77059 & n87254;
  assign n87256 = n87238 & n87251;
  assign n87257 = ~n87255 & n87256;
  assign n87258 = ~n87211 & n87214;
  assign n87259 = n87227 & n87258;
  assign n87260 = ~n87231 & n87259;
  assign n87261 = n87257 & n87260;
  assign n87262 = ~n87206 & n87261;
  assign n87263 = n85257 & ~n87262;
  assign n15631 = ~n87191 | n87263;
  assign n87265 = P2_P1_INSTADDRPOINTER_REG_21_ & n85256;
  assign n87266 = P2_P1_REIP_REG_21_ & n85401;
  assign n87267 = P2_P1_INSTADDRPOINTER_REG_20_ & n87207;
  assign n87268 = ~P2_P1_INSTADDRPOINTER_REG_21_ & n87267;
  assign n87269 = P2_P1_INSTADDRPOINTER_REG_21_ & ~n87267;
  assign n87270 = ~n87268 & ~n87269;
  assign n87271 = ~n77145 & ~n87270;
  assign n87272 = P2_P1_INSTADDRPOINTER_REG_20_ & n87215;
  assign n87273 = ~P2_P1_INSTADDRPOINTER_REG_21_ & n87272;
  assign n87274 = P2_P1_INSTADDRPOINTER_REG_21_ & ~n87272;
  assign n87275 = ~n87273 & ~n87274;
  assign n87276 = n77216 & ~n87275;
  assign n87277 = n77217 & ~n87275;
  assign n87278 = n85265 & ~n87270;
  assign n87279 = n77032 & ~n87275;
  assign n87280 = n85268 & ~n87270;
  assign n87281 = ~n87279 & ~n87280;
  assign n87282 = ~n87276 & ~n87277;
  assign n87283 = ~n87278 & n87282;
  assign n87284 = n87281 & n87283;
  assign n87285 = ~P2_P1_INSTADDRPOINTER_REG_21_ & ~n87229;
  assign n87286 = P2_P1_INSTADDRPOINTER_REG_21_ & n87229;
  assign n87287 = ~n87285 & ~n87286;
  assign n87288 = n85364 & n87287;
  assign n87289 = n76958 & ~n87275;
  assign n87290 = n77036 & ~n87275;
  assign n87291 = n77040 & ~n87275;
  assign n87292 = P2_P1_INSTADDRPOINTER_REG_20_ & n87242;
  assign n87293 = ~P2_P1_INSTADDRPOINTER_REG_21_ & n87292;
  assign n87294 = P2_P1_INSTADDRPOINTER_REG_21_ & ~n87292;
  assign n87295 = ~n87293 & ~n87294;
  assign n87296 = n77056 & ~n87295;
  assign n87297 = n77048 & ~n87295;
  assign n87298 = ~n87289 & ~n87290;
  assign n87299 = ~n87291 & n87298;
  assign n87300 = ~n87296 & n87299;
  assign n87301 = ~n87297 & n87300;
  assign n87302 = n85381 & ~n87270;
  assign n87303 = n77102 & ~n87270;
  assign n87304 = n85370 & ~n87270;
  assign n87305 = n85374 & ~n87270;
  assign n87306 = ~n87302 & ~n87303;
  assign n87307 = ~n87304 & n87306;
  assign n87308 = ~n87305 & n87307;
  assign n87309 = ~P2_P1_INSTADDRPOINTER_REG_21_ & ~n87253;
  assign n87310 = P2_P1_INSTADDRPOINTER_REG_20_ & P2_P1_INSTADDRPOINTER_REG_21_;
  assign n87311 = n87177 & n87310;
  assign n87312 = ~n87309 & ~n87311;
  assign n87313 = n77059 & n87312;
  assign n87314 = n87301 & n87308;
  assign n87315 = ~n87313 & n87314;
  assign n87316 = n77255 & ~n87270;
  assign n87317 = n77098 & ~n87270;
  assign n87318 = ~n87316 & ~n87317;
  assign n87319 = ~n87137 & n87192;
  assign n87320 = ~n87194 & ~n87319;
  assign n87321 = ~n86192 & ~n87198;
  assign n87322 = n87320 & ~n87321;
  assign n87323 = ~P2_P1_INSTADDRPOINTER_REG_21_ & ~n86192;
  assign n87324 = P2_P1_INSTADDRPOINTER_REG_21_ & n86192;
  assign n87325 = ~n87323 & ~n87324;
  assign n87326 = n87322 & ~n87325;
  assign n87327 = ~n87322 & n87325;
  assign n87328 = ~n87326 & ~n87327;
  assign n87329 = n85362 & ~n87328;
  assign n87330 = n87318 & ~n87329;
  assign n87331 = ~n87271 & n87284;
  assign n87332 = ~n87288 & n87331;
  assign n87333 = n87315 & n87332;
  assign n87334 = n87330 & n87333;
  assign n87335 = n85257 & ~n87334;
  assign n87336 = ~n87265 & ~n87266;
  assign n15636 = n87335 | ~n87336;
  assign n87338 = P2_P1_INSTADDRPOINTER_REG_22_ & n85256;
  assign n87339 = P2_P1_REIP_REG_22_ & n85401;
  assign n87340 = ~n87338 & ~n87339;
  assign n87341 = P2_P1_INSTADDRPOINTER_REG_21_ & n87292;
  assign n87342 = ~P2_P1_INSTADDRPOINTER_REG_22_ & n87341;
  assign n87343 = P2_P1_INSTADDRPOINTER_REG_22_ & ~n87341;
  assign n87344 = ~n87342 & ~n87343;
  assign n87345 = n77056 & ~n87344;
  assign n87346 = n77048 & ~n87344;
  assign n87347 = ~n87345 & ~n87346;
  assign n87348 = P2_P1_INSTADDRPOINTER_REG_21_ & n87272;
  assign n87349 = ~P2_P1_INSTADDRPOINTER_REG_22_ & n87348;
  assign n87350 = P2_P1_INSTADDRPOINTER_REG_22_ & ~n87348;
  assign n87351 = ~n87349 & ~n87350;
  assign n87352 = n76958 & ~n87351;
  assign n87353 = n77036 & ~n87351;
  assign n87354 = n77040 & ~n87351;
  assign n87355 = ~n87352 & ~n87353;
  assign n87356 = ~n87354 & n87355;
  assign n87357 = P2_P1_INSTADDRPOINTER_REG_21_ & n87267;
  assign n87358 = ~P2_P1_INSTADDRPOINTER_REG_22_ & n87357;
  assign n87359 = P2_P1_INSTADDRPOINTER_REG_22_ & ~n87357;
  assign n87360 = ~n87358 & ~n87359;
  assign n87361 = n85370 & ~n87360;
  assign n87362 = n85374 & ~n87360;
  assign n87363 = n77102 & ~n87360;
  assign n87364 = ~n87361 & ~n87362;
  assign n87365 = ~n87363 & n87364;
  assign n87366 = ~P2_P1_INSTADDRPOINTER_REG_22_ & n87311;
  assign n87367 = P2_P1_INSTADDRPOINTER_REG_22_ & ~n87311;
  assign n87368 = ~n87366 & ~n87367;
  assign n87369 = n77059 & ~n87368;
  assign n87370 = n85381 & ~n87360;
  assign n87371 = ~n87369 & ~n87370;
  assign n87372 = n87347 & n87356;
  assign n87373 = n87365 & n87372;
  assign n87374 = n87371 & n87373;
  assign n87375 = P2_P1_INSTADDRPOINTER_REG_21_ & n87192;
  assign n87376 = n86192 & ~n87375;
  assign n87377 = ~n87134 & ~n87376;
  assign n87378 = ~n87083 & n87377;
  assign n87379 = P2_P1_INSTADDRPOINTER_REG_21_ & ~n86192;
  assign n87380 = ~n87136 & ~n87379;
  assign n87381 = ~n87140 & n87380;
  assign n87382 = ~n87194 & n87381;
  assign n87383 = ~n87378 & n87382;
  assign n87384 = ~P2_P1_INSTADDRPOINTER_REG_22_ & ~n86192;
  assign n87385 = P2_P1_INSTADDRPOINTER_REG_22_ & n86192;
  assign n87386 = ~n87384 & ~n87385;
  assign n87387 = n87383 & ~n87386;
  assign n87388 = ~n87383 & n87386;
  assign n87389 = ~n87387 & ~n87388;
  assign n87390 = n85362 & ~n87389;
  assign n87391 = ~n77145 & ~n87360;
  assign n87392 = n77255 & ~n87360;
  assign n87393 = n77098 & ~n87360;
  assign n87394 = ~n87392 & ~n87393;
  assign n87395 = n77216 & ~n87351;
  assign n87396 = n77217 & ~n87351;
  assign n87397 = n85265 & ~n87360;
  assign n87398 = n77032 & ~n87351;
  assign n87399 = n85268 & ~n87360;
  assign n87400 = ~n87398 & ~n87399;
  assign n87401 = ~n87395 & ~n87396;
  assign n87402 = ~n87397 & n87401;
  assign n87403 = n87400 & n87402;
  assign n87404 = ~P2_P1_INSTADDRPOINTER_REG_22_ & n87286;
  assign n87405 = P2_P1_INSTADDRPOINTER_REG_22_ & ~n87286;
  assign n87406 = ~n87404 & ~n87405;
  assign n87407 = n85364 & ~n87406;
  assign n87408 = ~n87390 & ~n87391;
  assign n87409 = n87394 & n87408;
  assign n87410 = n87403 & n87409;
  assign n87411 = ~n87407 & n87410;
  assign n87412 = n87374 & n87411;
  assign n87413 = n85257 & ~n87412;
  assign n15641 = ~n87340 | n87413;
  assign n87415 = P2_P1_INSTADDRPOINTER_REG_23_ & n85256;
  assign n87416 = P2_P1_REIP_REG_23_ & n85401;
  assign n87417 = ~n87415 & ~n87416;
  assign n87418 = P2_P1_INSTADDRPOINTER_REG_22_ & n87341;
  assign n87419 = ~P2_P1_INSTADDRPOINTER_REG_23_ & n87418;
  assign n87420 = P2_P1_INSTADDRPOINTER_REG_23_ & ~n87418;
  assign n87421 = ~n87419 & ~n87420;
  assign n87422 = n77056 & ~n87421;
  assign n87423 = n77048 & ~n87421;
  assign n87424 = ~n87422 & ~n87423;
  assign n87425 = P2_P1_INSTADDRPOINTER_REG_22_ & n87348;
  assign n87426 = ~P2_P1_INSTADDRPOINTER_REG_23_ & n87425;
  assign n87427 = P2_P1_INSTADDRPOINTER_REG_23_ & ~n87425;
  assign n87428 = ~n87426 & ~n87427;
  assign n87429 = n76958 & ~n87428;
  assign n87430 = n77036 & ~n87428;
  assign n87431 = n77040 & ~n87428;
  assign n87432 = ~n87429 & ~n87430;
  assign n87433 = ~n87431 & n87432;
  assign n87434 = P2_P1_INSTADDRPOINTER_REG_22_ & n87357;
  assign n87435 = ~P2_P1_INSTADDRPOINTER_REG_23_ & n87434;
  assign n87436 = P2_P1_INSTADDRPOINTER_REG_23_ & ~n87434;
  assign n87437 = ~n87435 & ~n87436;
  assign n87438 = n85370 & ~n87437;
  assign n87439 = n85374 & ~n87437;
  assign n87440 = n77102 & ~n87437;
  assign n87441 = ~n87438 & ~n87439;
  assign n87442 = ~n87440 & n87441;
  assign n87443 = P2_P1_INSTADDRPOINTER_REG_22_ & n87311;
  assign n87444 = ~P2_P1_INSTADDRPOINTER_REG_23_ & ~n87443;
  assign n87445 = P2_P1_INSTADDRPOINTER_REG_22_ & P2_P1_INSTADDRPOINTER_REG_23_;
  assign n87446 = n87311 & n87445;
  assign n87447 = ~n87444 & ~n87446;
  assign n87448 = n77059 & n87447;
  assign n87449 = n85381 & ~n87437;
  assign n87450 = ~n87448 & ~n87449;
  assign n87451 = n87424 & n87433;
  assign n87452 = n87442 & n87451;
  assign n87453 = n87450 & n87452;
  assign n87454 = ~P2_P1_INSTADDRPOINTER_REG_22_ & n86192;
  assign n87455 = n87377 & ~n87454;
  assign n87456 = ~n87083 & n87455;
  assign n87457 = P2_P1_INSTADDRPOINTER_REG_22_ & ~n86192;
  assign n87458 = n87382 & ~n87457;
  assign n87459 = ~n87456 & n87458;
  assign n87460 = ~P2_P1_INSTADDRPOINTER_REG_23_ & ~n86192;
  assign n87461 = P2_P1_INSTADDRPOINTER_REG_23_ & n86192;
  assign n87462 = ~n87460 & ~n87461;
  assign n87463 = n87459 & ~n87462;
  assign n87464 = ~n87459 & n87462;
  assign n87465 = ~n87463 & ~n87464;
  assign n87466 = n85362 & ~n87465;
  assign n87467 = ~n77145 & ~n87437;
  assign n87468 = n77255 & ~n87437;
  assign n87469 = n77098 & ~n87437;
  assign n87470 = ~n87468 & ~n87469;
  assign n87471 = n77216 & ~n87428;
  assign n87472 = n77217 & ~n87428;
  assign n87473 = n85265 & ~n87437;
  assign n87474 = n77032 & ~n87428;
  assign n87475 = n85268 & ~n87437;
  assign n87476 = ~n87474 & ~n87475;
  assign n87477 = ~n87471 & ~n87472;
  assign n87478 = ~n87473 & n87477;
  assign n87479 = n87476 & n87478;
  assign n87480 = P2_P1_INSTADDRPOINTER_REG_22_ & n87286;
  assign n87481 = ~P2_P1_INSTADDRPOINTER_REG_23_ & ~n87480;
  assign n87482 = n87286 & n87445;
  assign n87483 = ~n87481 & ~n87482;
  assign n87484 = n85364 & n87483;
  assign n87485 = ~n87466 & ~n87467;
  assign n87486 = n87470 & n87485;
  assign n87487 = n87479 & n87486;
  assign n87488 = ~n87484 & n87487;
  assign n87489 = n87453 & n87488;
  assign n87490 = n85257 & ~n87489;
  assign n15646 = ~n87417 | n87490;
  assign n87492 = P2_P1_INSTADDRPOINTER_REG_24_ & n85256;
  assign n87493 = P2_P1_REIP_REG_24_ & n85401;
  assign n87494 = ~n87492 & ~n87493;
  assign n87495 = P2_P1_INSTADDRPOINTER_REG_23_ & n87418;
  assign n87496 = ~P2_P1_INSTADDRPOINTER_REG_24_ & n87495;
  assign n87497 = P2_P1_INSTADDRPOINTER_REG_24_ & ~n87495;
  assign n87498 = ~n87496 & ~n87497;
  assign n87499 = n77056 & ~n87498;
  assign n87500 = n77048 & ~n87498;
  assign n87501 = ~n87499 & ~n87500;
  assign n87502 = P2_P1_INSTADDRPOINTER_REG_23_ & n87425;
  assign n87503 = ~P2_P1_INSTADDRPOINTER_REG_24_ & n87502;
  assign n87504 = P2_P1_INSTADDRPOINTER_REG_24_ & ~n87502;
  assign n87505 = ~n87503 & ~n87504;
  assign n87506 = n76958 & ~n87505;
  assign n87507 = n77036 & ~n87505;
  assign n87508 = n77040 & ~n87505;
  assign n87509 = ~n87506 & ~n87507;
  assign n87510 = ~n87508 & n87509;
  assign n87511 = ~P2_P1_INSTADDRPOINTER_REG_24_ & n87446;
  assign n87512 = P2_P1_INSTADDRPOINTER_REG_24_ & ~n87446;
  assign n87513 = ~n87511 & ~n87512;
  assign n87514 = n77059 & ~n87513;
  assign n87515 = P2_P1_INSTADDRPOINTER_REG_23_ & n87434;
  assign n87516 = ~P2_P1_INSTADDRPOINTER_REG_24_ & n87515;
  assign n87517 = P2_P1_INSTADDRPOINTER_REG_24_ & ~n87515;
  assign n87518 = ~n87516 & ~n87517;
  assign n87519 = n85381 & ~n87518;
  assign n87520 = ~n87514 & ~n87519;
  assign n87521 = n85370 & ~n87518;
  assign n87522 = n85374 & ~n87518;
  assign n87523 = n77102 & ~n87518;
  assign n87524 = ~n87521 & ~n87522;
  assign n87525 = ~n87523 & n87524;
  assign n87526 = n87501 & n87510;
  assign n87527 = n87520 & n87526;
  assign n87528 = n87525 & n87527;
  assign n87529 = P2_P1_INSTADDRPOINTER_REG_23_ & ~n86192;
  assign n87530 = n87458 & ~n87529;
  assign n87531 = ~P2_P1_INSTADDRPOINTER_REG_23_ & n86192;
  assign n87532 = n87455 & ~n87531;
  assign n87533 = ~n87083 & n87532;
  assign n87534 = n87530 & ~n87533;
  assign n87535 = ~P2_P1_INSTADDRPOINTER_REG_24_ & ~n86192;
  assign n87536 = P2_P1_INSTADDRPOINTER_REG_24_ & n86192;
  assign n87537 = ~n87535 & ~n87536;
  assign n87538 = n87534 & ~n87537;
  assign n87539 = ~n87534 & n87537;
  assign n87540 = ~n87538 & ~n87539;
  assign n87541 = n85362 & ~n87540;
  assign n87542 = ~n77145 & ~n87518;
  assign n87543 = n77255 & ~n87518;
  assign n87544 = n77098 & ~n87518;
  assign n87545 = ~n87543 & ~n87544;
  assign n87546 = ~P2_P1_INSTADDRPOINTER_REG_24_ & n87482;
  assign n87547 = P2_P1_INSTADDRPOINTER_REG_24_ & ~n87482;
  assign n87548 = ~n87546 & ~n87547;
  assign n87549 = n85364 & ~n87548;
  assign n87550 = n77216 & ~n87505;
  assign n87551 = n77217 & ~n87505;
  assign n87552 = n85265 & ~n87518;
  assign n87553 = n77032 & ~n87505;
  assign n87554 = n85268 & ~n87518;
  assign n87555 = ~n87553 & ~n87554;
  assign n87556 = ~n87550 & ~n87551;
  assign n87557 = ~n87552 & n87556;
  assign n87558 = n87555 & n87557;
  assign n87559 = ~n87541 & ~n87542;
  assign n87560 = n87545 & n87559;
  assign n87561 = ~n87549 & n87560;
  assign n87562 = n87558 & n87561;
  assign n87563 = n87528 & n87562;
  assign n87564 = n85257 & ~n87563;
  assign n15651 = ~n87494 | n87564;
  assign n87566 = P2_P1_INSTADDRPOINTER_REG_25_ & n85256;
  assign n87567 = P2_P1_REIP_REG_25_ & n85401;
  assign n87568 = ~n87566 & ~n87567;
  assign n87569 = P2_P1_INSTADDRPOINTER_REG_24_ & n87495;
  assign n87570 = ~P2_P1_INSTADDRPOINTER_REG_25_ & n87569;
  assign n87571 = P2_P1_INSTADDRPOINTER_REG_25_ & ~n87569;
  assign n87572 = ~n87570 & ~n87571;
  assign n87573 = n77056 & ~n87572;
  assign n87574 = n77048 & ~n87572;
  assign n87575 = ~n87573 & ~n87574;
  assign n87576 = P2_P1_INSTADDRPOINTER_REG_24_ & n87502;
  assign n87577 = ~P2_P1_INSTADDRPOINTER_REG_25_ & n87576;
  assign n87578 = P2_P1_INSTADDRPOINTER_REG_25_ & ~n87576;
  assign n87579 = ~n87577 & ~n87578;
  assign n87580 = n76958 & ~n87579;
  assign n87581 = n77036 & ~n87579;
  assign n87582 = n77040 & ~n87579;
  assign n87583 = ~n87580 & ~n87581;
  assign n87584 = ~n87582 & n87583;
  assign n87585 = P2_P1_INSTADDRPOINTER_REG_24_ & n87446;
  assign n87586 = ~P2_P1_INSTADDRPOINTER_REG_25_ & ~n87585;
  assign n87587 = P2_P1_INSTADDRPOINTER_REG_24_ & P2_P1_INSTADDRPOINTER_REG_25_;
  assign n87588 = n87446 & n87587;
  assign n87589 = ~n87586 & ~n87588;
  assign n87590 = n77059 & n87589;
  assign n87591 = P2_P1_INSTADDRPOINTER_REG_24_ & n87515;
  assign n87592 = ~P2_P1_INSTADDRPOINTER_REG_25_ & n87591;
  assign n87593 = P2_P1_INSTADDRPOINTER_REG_25_ & ~n87591;
  assign n87594 = ~n87592 & ~n87593;
  assign n87595 = n85381 & ~n87594;
  assign n87596 = ~n87590 & ~n87595;
  assign n87597 = n85370 & ~n87594;
  assign n87598 = n85374 & ~n87594;
  assign n87599 = n77102 & ~n87594;
  assign n87600 = ~n87597 & ~n87598;
  assign n87601 = ~n87599 & n87600;
  assign n87602 = n87575 & n87584;
  assign n87603 = n87596 & n87602;
  assign n87604 = n87601 & n87603;
  assign n87605 = ~P2_P1_INSTADDRPOINTER_REG_25_ & ~n86192;
  assign n87606 = P2_P1_INSTADDRPOINTER_REG_25_ & n86192;
  assign n87607 = ~n87605 & ~n87606;
  assign n87608 = P2_P1_INSTADDRPOINTER_REG_24_ & ~n86192;
  assign n87609 = ~P2_P1_INSTADDRPOINTER_REG_24_ & n86192;
  assign n87610 = ~n87534 & ~n87609;
  assign n87611 = ~n87608 & ~n87610;
  assign n87612 = ~n87607 & n87611;
  assign n87613 = ~P2_P1_INSTADDRPOINTER_REG_25_ & n86192;
  assign n87614 = P2_P1_INSTADDRPOINTER_REG_25_ & ~n86192;
  assign n87615 = ~n87613 & ~n87614;
  assign n87616 = ~n87611 & ~n87615;
  assign n87617 = ~n87612 & ~n87616;
  assign n87618 = n85362 & ~n87617;
  assign n87619 = ~n77145 & ~n87594;
  assign n87620 = P2_P1_INSTADDRPOINTER_REG_24_ & n87482;
  assign n87621 = ~P2_P1_INSTADDRPOINTER_REG_25_ & ~n87620;
  assign n87622 = n87482 & n87587;
  assign n87623 = ~n87621 & ~n87622;
  assign n87624 = n85364 & n87623;
  assign n87625 = n77255 & ~n87594;
  assign n87626 = n77098 & ~n87594;
  assign n87627 = ~n87625 & ~n87626;
  assign n87628 = n77216 & ~n87579;
  assign n87629 = n77217 & ~n87579;
  assign n87630 = n85265 & ~n87594;
  assign n87631 = n77032 & ~n87579;
  assign n87632 = n85268 & ~n87594;
  assign n87633 = ~n87631 & ~n87632;
  assign n87634 = ~n87628 & ~n87629;
  assign n87635 = ~n87630 & n87634;
  assign n87636 = n87633 & n87635;
  assign n87637 = ~n87618 & ~n87619;
  assign n87638 = ~n87624 & n87637;
  assign n87639 = n87627 & n87638;
  assign n87640 = n87636 & n87639;
  assign n87641 = n87604 & n87640;
  assign n87642 = n85257 & ~n87641;
  assign n15656 = ~n87568 | n87642;
  assign n87644 = P2_P1_INSTADDRPOINTER_REG_26_ & n85256;
  assign n87645 = P2_P1_REIP_REG_26_ & n85401;
  assign n87646 = P2_P1_INSTADDRPOINTER_REG_26_ & ~n86192;
  assign n87647 = P2_P1_INSTADDRPOINTER_REG_25_ & P2_P1_INSTADDRPOINTER_REG_26_;
  assign n87648 = n86192 & ~n87647;
  assign n87649 = ~n87646 & ~n87648;
  assign n87650 = n87611 & ~n87614;
  assign n87651 = n87649 & ~n87650;
  assign n87652 = ~P2_P1_INSTADDRPOINTER_REG_26_ & ~n86192;
  assign n87653 = P2_P1_INSTADDRPOINTER_REG_26_ & n86192;
  assign n87654 = ~n87652 & ~n87653;
  assign n87655 = ~n87614 & n87654;
  assign n87656 = ~n87611 & ~n87613;
  assign n87657 = n87655 & ~n87656;
  assign n87658 = ~n87651 & ~n87657;
  assign n87659 = n85362 & n87658;
  assign n87660 = ~P2_P1_INSTADDRPOINTER_REG_26_ & ~n87622;
  assign n87661 = P2_P1_INSTADDRPOINTER_REG_26_ & n87622;
  assign n87662 = ~n87660 & ~n87661;
  assign n87663 = n85364 & n87662;
  assign n87664 = ~n87659 & ~n87663;
  assign n87665 = P2_P1_INSTADDRPOINTER_REG_25_ & n87591;
  assign n87666 = ~P2_P1_INSTADDRPOINTER_REG_26_ & n87665;
  assign n87667 = P2_P1_INSTADDRPOINTER_REG_26_ & ~n87665;
  assign n87668 = ~n87666 & ~n87667;
  assign n87669 = ~n77145 & ~n87668;
  assign n87670 = n77255 & ~n87668;
  assign n87671 = n77098 & ~n87668;
  assign n87672 = ~n87670 & ~n87671;
  assign n87673 = P2_P1_INSTADDRPOINTER_REG_25_ & n87576;
  assign n87674 = ~P2_P1_INSTADDRPOINTER_REG_26_ & n87673;
  assign n87675 = P2_P1_INSTADDRPOINTER_REG_26_ & ~n87673;
  assign n87676 = ~n87674 & ~n87675;
  assign n87677 = n77216 & ~n87676;
  assign n87678 = n77217 & ~n87676;
  assign n87679 = n85265 & ~n87668;
  assign n87680 = n77032 & ~n87676;
  assign n87681 = n85268 & ~n87668;
  assign n87682 = ~n87680 & ~n87681;
  assign n87683 = ~n87677 & ~n87678;
  assign n87684 = ~n87679 & n87683;
  assign n87685 = n87682 & n87684;
  assign n87686 = P2_P1_INSTADDRPOINTER_REG_25_ & n87569;
  assign n87687 = ~P2_P1_INSTADDRPOINTER_REG_26_ & n87686;
  assign n87688 = P2_P1_INSTADDRPOINTER_REG_26_ & ~n87686;
  assign n87689 = ~n87687 & ~n87688;
  assign n87690 = n77056 & ~n87689;
  assign n87691 = n77048 & ~n87689;
  assign n87692 = ~n87690 & ~n87691;
  assign n87693 = n76958 & ~n87676;
  assign n87694 = n77036 & ~n87676;
  assign n87695 = n77040 & ~n87676;
  assign n87696 = ~n87693 & ~n87694;
  assign n87697 = ~n87695 & n87696;
  assign n87698 = ~P2_P1_INSTADDRPOINTER_REG_26_ & ~n87588;
  assign n87699 = P2_P1_INSTADDRPOINTER_REG_26_ & n87588;
  assign n87700 = ~n87698 & ~n87699;
  assign n87701 = n77059 & n87700;
  assign n87702 = n85381 & ~n87668;
  assign n87703 = ~n87701 & ~n87702;
  assign n87704 = n85370 & ~n87668;
  assign n87705 = n85374 & ~n87668;
  assign n87706 = n77102 & ~n87668;
  assign n87707 = ~n87704 & ~n87705;
  assign n87708 = ~n87706 & n87707;
  assign n87709 = n87692 & n87697;
  assign n87710 = n87703 & n87709;
  assign n87711 = n87708 & n87710;
  assign n87712 = n87664 & ~n87669;
  assign n87713 = n87672 & n87712;
  assign n87714 = n87685 & n87713;
  assign n87715 = n87711 & n87714;
  assign n87716 = n85257 & ~n87715;
  assign n87717 = ~n87644 & ~n87645;
  assign n15661 = n87716 | ~n87717;
  assign n87719 = P2_P1_INSTADDRPOINTER_REG_27_ & n85256;
  assign n87720 = P2_P1_REIP_REG_27_ & n85401;
  assign n87721 = ~n87614 & ~n87646;
  assign n87722 = ~n87611 & ~n87648;
  assign n87723 = n87721 & ~n87722;
  assign n87724 = ~P2_P1_INSTADDRPOINTER_REG_27_ & ~n86192;
  assign n87725 = P2_P1_INSTADDRPOINTER_REG_27_ & n86192;
  assign n87726 = ~n87724 & ~n87725;
  assign n87727 = n87723 & ~n87726;
  assign n87728 = ~n87723 & n87726;
  assign n87729 = ~n87727 & ~n87728;
  assign n87730 = n85362 & ~n87729;
  assign n87731 = ~P2_P1_INSTADDRPOINTER_REG_27_ & n87661;
  assign n87732 = P2_P1_INSTADDRPOINTER_REG_27_ & ~n87661;
  assign n87733 = ~n87731 & ~n87732;
  assign n87734 = n85364 & ~n87733;
  assign n87735 = ~n87730 & ~n87734;
  assign n87736 = P2_P1_INSTADDRPOINTER_REG_26_ & n87665;
  assign n87737 = ~P2_P1_INSTADDRPOINTER_REG_27_ & n87736;
  assign n87738 = P2_P1_INSTADDRPOINTER_REG_27_ & ~n87736;
  assign n87739 = ~n87737 & ~n87738;
  assign n87740 = ~n77145 & ~n87739;
  assign n87741 = n77255 & ~n87739;
  assign n87742 = n77098 & ~n87739;
  assign n87743 = ~n87741 & ~n87742;
  assign n87744 = P2_P1_INSTADDRPOINTER_REG_26_ & n87673;
  assign n87745 = ~P2_P1_INSTADDRPOINTER_REG_27_ & n87744;
  assign n87746 = P2_P1_INSTADDRPOINTER_REG_27_ & ~n87744;
  assign n87747 = ~n87745 & ~n87746;
  assign n87748 = n77216 & ~n87747;
  assign n87749 = n77217 & ~n87747;
  assign n87750 = n85265 & ~n87739;
  assign n87751 = n77032 & ~n87747;
  assign n87752 = n85268 & ~n87739;
  assign n87753 = ~n87751 & ~n87752;
  assign n87754 = ~n87748 & ~n87749;
  assign n87755 = ~n87750 & n87754;
  assign n87756 = n87753 & n87755;
  assign n87757 = P2_P1_INSTADDRPOINTER_REG_26_ & n87686;
  assign n87758 = ~P2_P1_INSTADDRPOINTER_REG_27_ & n87757;
  assign n87759 = P2_P1_INSTADDRPOINTER_REG_27_ & ~n87757;
  assign n87760 = ~n87758 & ~n87759;
  assign n87761 = n77056 & ~n87760;
  assign n87762 = n77048 & ~n87760;
  assign n87763 = ~n87761 & ~n87762;
  assign n87764 = n76958 & ~n87747;
  assign n87765 = n77036 & ~n87747;
  assign n87766 = n77040 & ~n87747;
  assign n87767 = ~n87764 & ~n87765;
  assign n87768 = ~n87766 & n87767;
  assign n87769 = ~P2_P1_INSTADDRPOINTER_REG_27_ & n87699;
  assign n87770 = P2_P1_INSTADDRPOINTER_REG_27_ & ~n87699;
  assign n87771 = ~n87769 & ~n87770;
  assign n87772 = n77059 & ~n87771;
  assign n87773 = n85381 & ~n87739;
  assign n87774 = ~n87772 & ~n87773;
  assign n87775 = n85370 & ~n87739;
  assign n87776 = n85374 & ~n87739;
  assign n87777 = n77102 & ~n87739;
  assign n87778 = ~n87775 & ~n87776;
  assign n87779 = ~n87777 & n87778;
  assign n87780 = n87763 & n87768;
  assign n87781 = n87774 & n87780;
  assign n87782 = n87779 & n87781;
  assign n87783 = n87735 & ~n87740;
  assign n87784 = n87743 & n87783;
  assign n87785 = n87756 & n87784;
  assign n87786 = n87782 & n87785;
  assign n87787 = n85257 & ~n87786;
  assign n87788 = ~n87719 & ~n87720;
  assign n15666 = n87787 | ~n87788;
  assign n87790 = P2_P1_INSTADDRPOINTER_REG_28_ & n85256;
  assign n87791 = P2_P1_REIP_REG_28_ & n85401;
  assign n87792 = P2_P1_INSTADDRPOINTER_REG_27_ & P2_P1_INSTADDRPOINTER_REG_28_;
  assign n87793 = ~n87723 & n87792;
  assign n87794 = n86192 & ~n87793;
  assign n87795 = P2_P1_INSTADDRPOINTER_REG_28_ & ~n86192;
  assign n87796 = ~P2_P1_INSTADDRPOINTER_REG_27_ & ~n87614;
  assign n87797 = ~n87646 & n87796;
  assign n87798 = ~n87722 & n87797;
  assign n87799 = ~n87794 & ~n87795;
  assign n87800 = ~n87798 & n87799;
  assign n87801 = P2_P1_INSTADDRPOINTER_REG_28_ & n87798;
  assign n87802 = ~n86192 & ~n87801;
  assign n87803 = P2_P1_INSTADDRPOINTER_REG_28_ & n86192;
  assign n87804 = P2_P1_INSTADDRPOINTER_REG_27_ & ~n87723;
  assign n87805 = ~n87802 & ~n87803;
  assign n87806 = ~n87804 & n87805;
  assign n87807 = ~n87800 & ~n87806;
  assign n87808 = n85362 & n87807;
  assign n87809 = P2_P1_INSTADDRPOINTER_REG_27_ & n87661;
  assign n87810 = ~P2_P1_INSTADDRPOINTER_REG_28_ & ~n87809;
  assign n87811 = n87661 & n87792;
  assign n87812 = ~n87810 & ~n87811;
  assign n87813 = n85364 & n87812;
  assign n87814 = ~n87808 & ~n87813;
  assign n87815 = P2_P1_INSTADDRPOINTER_REG_27_ & n87736;
  assign n87816 = ~P2_P1_INSTADDRPOINTER_REG_28_ & n87815;
  assign n87817 = P2_P1_INSTADDRPOINTER_REG_28_ & ~n87815;
  assign n87818 = ~n87816 & ~n87817;
  assign n87819 = ~n77145 & ~n87818;
  assign n87820 = n77255 & ~n87818;
  assign n87821 = n77098 & ~n87818;
  assign n87822 = ~n87820 & ~n87821;
  assign n87823 = P2_P1_INSTADDRPOINTER_REG_27_ & n87744;
  assign n87824 = ~P2_P1_INSTADDRPOINTER_REG_28_ & n87823;
  assign n87825 = P2_P1_INSTADDRPOINTER_REG_28_ & ~n87823;
  assign n87826 = ~n87824 & ~n87825;
  assign n87827 = n77216 & ~n87826;
  assign n87828 = n77217 & ~n87826;
  assign n87829 = n85265 & ~n87818;
  assign n87830 = n77032 & ~n87826;
  assign n87831 = n85268 & ~n87818;
  assign n87832 = ~n87830 & ~n87831;
  assign n87833 = ~n87827 & ~n87828;
  assign n87834 = ~n87829 & n87833;
  assign n87835 = n87832 & n87834;
  assign n87836 = P2_P1_INSTADDRPOINTER_REG_27_ & n87757;
  assign n87837 = ~P2_P1_INSTADDRPOINTER_REG_28_ & n87836;
  assign n87838 = P2_P1_INSTADDRPOINTER_REG_28_ & ~n87836;
  assign n87839 = ~n87837 & ~n87838;
  assign n87840 = n77056 & ~n87839;
  assign n87841 = n77048 & ~n87839;
  assign n87842 = ~n87840 & ~n87841;
  assign n87843 = n76958 & ~n87826;
  assign n87844 = n77036 & ~n87826;
  assign n87845 = n77040 & ~n87826;
  assign n87846 = ~n87843 & ~n87844;
  assign n87847 = ~n87845 & n87846;
  assign n87848 = P2_P1_INSTADDRPOINTER_REG_27_ & n87699;
  assign n87849 = ~P2_P1_INSTADDRPOINTER_REG_28_ & ~n87848;
  assign n87850 = n87699 & n87792;
  assign n87851 = ~n87849 & ~n87850;
  assign n87852 = n77059 & n87851;
  assign n87853 = n85381 & ~n87818;
  assign n87854 = ~n87852 & ~n87853;
  assign n87855 = n85370 & ~n87818;
  assign n87856 = n85374 & ~n87818;
  assign n87857 = n77102 & ~n87818;
  assign n87858 = ~n87855 & ~n87856;
  assign n87859 = ~n87857 & n87858;
  assign n87860 = n87842 & n87847;
  assign n87861 = n87854 & n87860;
  assign n87862 = n87859 & n87861;
  assign n87863 = n87814 & ~n87819;
  assign n87864 = n87822 & n87863;
  assign n87865 = n87835 & n87864;
  assign n87866 = n87862 & n87865;
  assign n87867 = n85257 & ~n87866;
  assign n87868 = ~n87790 & ~n87791;
  assign n15671 = n87867 | ~n87868;
  assign n87870 = P2_P1_INSTADDRPOINTER_REG_29_ & n85256;
  assign n87871 = P2_P1_REIP_REG_29_ & n85401;
  assign n87872 = ~n86192 & ~n87798;
  assign n87873 = ~n87795 & ~n87872;
  assign n87874 = ~n87793 & n87873;
  assign n87875 = ~P2_P1_INSTADDRPOINTER_REG_29_ & ~n86192;
  assign n87876 = P2_P1_INSTADDRPOINTER_REG_29_ & n86192;
  assign n87877 = ~n87875 & ~n87876;
  assign n87878 = n87874 & ~n87877;
  assign n87879 = ~n87874 & n87877;
  assign n87880 = ~n87878 & ~n87879;
  assign n87881 = n85362 & ~n87880;
  assign n87882 = ~P2_P1_INSTADDRPOINTER_REG_29_ & ~n87811;
  assign n87883 = P2_P1_INSTADDRPOINTER_REG_29_ & n87811;
  assign n87884 = ~n87882 & ~n87883;
  assign n87885 = n85364 & n87884;
  assign n87886 = ~n87881 & ~n87885;
  assign n87887 = P2_P1_INSTADDRPOINTER_REG_28_ & n87815;
  assign n87888 = ~P2_P1_INSTADDRPOINTER_REG_29_ & n87887;
  assign n87889 = P2_P1_INSTADDRPOINTER_REG_29_ & ~n87887;
  assign n87890 = ~n87888 & ~n87889;
  assign n87891 = ~n77145 & ~n87890;
  assign n87892 = n77255 & ~n87890;
  assign n87893 = n77098 & ~n87890;
  assign n87894 = ~n87892 & ~n87893;
  assign n87895 = P2_P1_INSTADDRPOINTER_REG_28_ & n87823;
  assign n87896 = ~P2_P1_INSTADDRPOINTER_REG_29_ & n87895;
  assign n87897 = P2_P1_INSTADDRPOINTER_REG_29_ & ~n87895;
  assign n87898 = ~n87896 & ~n87897;
  assign n87899 = n77216 & ~n87898;
  assign n87900 = n77217 & ~n87898;
  assign n87901 = n85265 & ~n87890;
  assign n87902 = n77032 & ~n87898;
  assign n87903 = n85268 & ~n87890;
  assign n87904 = ~n87902 & ~n87903;
  assign n87905 = ~n87899 & ~n87900;
  assign n87906 = ~n87901 & n87905;
  assign n87907 = n87904 & n87906;
  assign n87908 = P2_P1_INSTADDRPOINTER_REG_28_ & n87836;
  assign n87909 = ~P2_P1_INSTADDRPOINTER_REG_29_ & n87908;
  assign n87910 = P2_P1_INSTADDRPOINTER_REG_29_ & ~n87908;
  assign n87911 = ~n87909 & ~n87910;
  assign n87912 = n77056 & ~n87911;
  assign n87913 = n77048 & ~n87911;
  assign n87914 = ~n87912 & ~n87913;
  assign n87915 = n76958 & ~n87898;
  assign n87916 = n77036 & ~n87898;
  assign n87917 = n77040 & ~n87898;
  assign n87918 = ~n87915 & ~n87916;
  assign n87919 = ~n87917 & n87918;
  assign n87920 = ~P2_P1_INSTADDRPOINTER_REG_29_ & ~n87850;
  assign n87921 = P2_P1_INSTADDRPOINTER_REG_29_ & n87850;
  assign n87922 = ~n87920 & ~n87921;
  assign n87923 = n77059 & n87922;
  assign n87924 = n85381 & ~n87890;
  assign n87925 = ~n87923 & ~n87924;
  assign n87926 = n85370 & ~n87890;
  assign n87927 = n85374 & ~n87890;
  assign n87928 = n77102 & ~n87890;
  assign n87929 = ~n87926 & ~n87927;
  assign n87930 = ~n87928 & n87929;
  assign n87931 = n87914 & n87919;
  assign n87932 = n87925 & n87931;
  assign n87933 = n87930 & n87932;
  assign n87934 = n87886 & ~n87891;
  assign n87935 = n87894 & n87934;
  assign n87936 = n87907 & n87935;
  assign n87937 = n87933 & n87936;
  assign n87938 = n85257 & ~n87937;
  assign n87939 = ~n87870 & ~n87871;
  assign n15676 = n87938 | ~n87939;
  assign n87941 = P2_P1_INSTADDRPOINTER_REG_30_ & n85256;
  assign n87942 = P2_P1_REIP_REG_30_ & n85401;
  assign n87943 = ~P2_P1_INSTADDRPOINTER_REG_30_ & ~n86192;
  assign n87944 = P2_P1_INSTADDRPOINTER_REG_30_ & n86192;
  assign n87945 = ~n87943 & ~n87944;
  assign n87946 = P2_P1_INSTADDRPOINTER_REG_29_ & ~n86192;
  assign n87947 = ~P2_P1_INSTADDRPOINTER_REG_29_ & n86192;
  assign n87948 = ~n87874 & ~n87947;
  assign n87949 = ~n87946 & ~n87948;
  assign n87950 = ~n87945 & n87949;
  assign n87951 = n87945 & ~n87949;
  assign n87952 = ~n87950 & ~n87951;
  assign n87953 = n85362 & ~n87952;
  assign n87954 = ~P2_P1_INSTADDRPOINTER_REG_30_ & n87883;
  assign n87955 = P2_P1_INSTADDRPOINTER_REG_30_ & ~n87883;
  assign n87956 = ~n87954 & ~n87955;
  assign n87957 = n85364 & ~n87956;
  assign n87958 = ~n87953 & ~n87957;
  assign n87959 = P2_P1_INSTADDRPOINTER_REG_29_ & n87887;
  assign n87960 = ~P2_P1_INSTADDRPOINTER_REG_30_ & n87959;
  assign n87961 = P2_P1_INSTADDRPOINTER_REG_30_ & ~n87959;
  assign n87962 = ~n87960 & ~n87961;
  assign n87963 = ~n77145 & ~n87962;
  assign n87964 = n77255 & ~n87962;
  assign n87965 = n77098 & ~n87962;
  assign n87966 = ~n87964 & ~n87965;
  assign n87967 = P2_P1_INSTADDRPOINTER_REG_29_ & n87895;
  assign n87968 = ~P2_P1_INSTADDRPOINTER_REG_30_ & n87967;
  assign n87969 = P2_P1_INSTADDRPOINTER_REG_30_ & ~n87967;
  assign n87970 = ~n87968 & ~n87969;
  assign n87971 = n77216 & ~n87970;
  assign n87972 = n77217 & ~n87970;
  assign n87973 = n85265 & ~n87962;
  assign n87974 = n77032 & ~n87970;
  assign n87975 = n85268 & ~n87962;
  assign n87976 = ~n87974 & ~n87975;
  assign n87977 = ~n87971 & ~n87972;
  assign n87978 = ~n87973 & n87977;
  assign n87979 = n87976 & n87978;
  assign n87980 = P2_P1_INSTADDRPOINTER_REG_29_ & n87908;
  assign n87981 = ~P2_P1_INSTADDRPOINTER_REG_30_ & n87980;
  assign n87982 = P2_P1_INSTADDRPOINTER_REG_30_ & ~n87980;
  assign n87983 = ~n87981 & ~n87982;
  assign n87984 = n77056 & ~n87983;
  assign n87985 = n77048 & ~n87983;
  assign n87986 = ~n87984 & ~n87985;
  assign n87987 = n76958 & ~n87970;
  assign n87988 = n77036 & ~n87970;
  assign n87989 = n77040 & ~n87970;
  assign n87990 = ~n87987 & ~n87988;
  assign n87991 = ~n87989 & n87990;
  assign n87992 = ~P2_P1_INSTADDRPOINTER_REG_30_ & n87921;
  assign n87993 = P2_P1_INSTADDRPOINTER_REG_30_ & ~n87921;
  assign n87994 = ~n87992 & ~n87993;
  assign n87995 = n77059 & ~n87994;
  assign n87996 = n85381 & ~n87962;
  assign n87997 = ~n87995 & ~n87996;
  assign n87998 = n85370 & ~n87962;
  assign n87999 = n85374 & ~n87962;
  assign n88000 = n77102 & ~n87962;
  assign n88001 = ~n87998 & ~n87999;
  assign n88002 = ~n88000 & n88001;
  assign n88003 = n87986 & n87991;
  assign n88004 = n87997 & n88003;
  assign n88005 = n88002 & n88004;
  assign n88006 = n87958 & ~n87963;
  assign n88007 = n87966 & n88006;
  assign n88008 = n87979 & n88007;
  assign n88009 = n88005 & n88008;
  assign n88010 = n85257 & ~n88009;
  assign n88011 = ~n87941 & ~n87942;
  assign n15681 = n88010 | ~n88011;
  assign n88013 = P2_P1_INSTADDRPOINTER_REG_31_ & n85256;
  assign n88014 = P2_P1_REIP_REG_31_ & n85401;
  assign n88015 = P2_P1_INSTADDRPOINTER_REG_30_ & P2_P1_INSTADDRPOINTER_REG_31_;
  assign n88016 = ~n87949 & n88015;
  assign n88017 = n86192 & ~n88016;
  assign n88018 = P2_P1_INSTADDRPOINTER_REG_31_ & ~n86192;
  assign n88019 = ~P2_P1_INSTADDRPOINTER_REG_30_ & n87949;
  assign n88020 = ~n88017 & ~n88018;
  assign n88021 = ~n88019 & n88020;
  assign n88022 = ~P2_P1_INSTADDRPOINTER_REG_30_ & P2_P1_INSTADDRPOINTER_REG_31_;
  assign n88023 = ~n87946 & n88022;
  assign n88024 = ~n87948 & n88023;
  assign n88025 = ~n86192 & ~n88024;
  assign n88026 = P2_P1_INSTADDRPOINTER_REG_31_ & n86192;
  assign n88027 = P2_P1_INSTADDRPOINTER_REG_30_ & ~n87949;
  assign n88028 = ~n88025 & ~n88026;
  assign n88029 = ~n88027 & n88028;
  assign n88030 = ~n88021 & ~n88029;
  assign n88031 = n85362 & n88030;
  assign n88032 = P2_P1_INSTADDRPOINTER_REG_30_ & n87883;
  assign n88033 = ~P2_P1_INSTADDRPOINTER_REG_31_ & n88032;
  assign n88034 = P2_P1_INSTADDRPOINTER_REG_31_ & ~n88032;
  assign n88035 = ~n88033 & ~n88034;
  assign n88036 = n85364 & ~n88035;
  assign n88037 = ~n88031 & ~n88036;
  assign n88038 = P2_P1_INSTADDRPOINTER_REG_30_ & n87959;
  assign n88039 = ~P2_P1_INSTADDRPOINTER_REG_31_ & n88038;
  assign n88040 = P2_P1_INSTADDRPOINTER_REG_31_ & ~n88038;
  assign n88041 = ~n88039 & ~n88040;
  assign n88042 = ~n77145 & ~n88041;
  assign n88043 = n77255 & ~n88041;
  assign n88044 = n77098 & ~n88041;
  assign n88045 = ~n88043 & ~n88044;
  assign n88046 = P2_P1_INSTADDRPOINTER_REG_30_ & n87967;
  assign n88047 = ~P2_P1_INSTADDRPOINTER_REG_31_ & n88046;
  assign n88048 = P2_P1_INSTADDRPOINTER_REG_31_ & ~n88046;
  assign n88049 = ~n88047 & ~n88048;
  assign n88050 = n77216 & ~n88049;
  assign n88051 = n77217 & ~n88049;
  assign n88052 = n85265 & ~n88041;
  assign n88053 = n77032 & ~n88049;
  assign n88054 = n85268 & ~n88041;
  assign n88055 = ~n88053 & ~n88054;
  assign n88056 = ~n88050 & ~n88051;
  assign n88057 = ~n88052 & n88056;
  assign n88058 = n88055 & n88057;
  assign n88059 = P2_P1_INSTADDRPOINTER_REG_30_ & n87980;
  assign n88060 = ~P2_P1_INSTADDRPOINTER_REG_31_ & n88059;
  assign n88061 = P2_P1_INSTADDRPOINTER_REG_31_ & ~n88059;
  assign n88062 = ~n88060 & ~n88061;
  assign n88063 = n77056 & ~n88062;
  assign n88064 = n77048 & ~n88062;
  assign n88065 = ~n88063 & ~n88064;
  assign n88066 = n76958 & ~n88049;
  assign n88067 = n77036 & ~n88049;
  assign n88068 = n77040 & ~n88049;
  assign n88069 = ~n88066 & ~n88067;
  assign n88070 = ~n88068 & n88069;
  assign n88071 = P2_P1_INSTADDRPOINTER_REG_30_ & n87921;
  assign n88072 = ~P2_P1_INSTADDRPOINTER_REG_31_ & n88071;
  assign n88073 = P2_P1_INSTADDRPOINTER_REG_31_ & ~n88071;
  assign n88074 = ~n88072 & ~n88073;
  assign n88075 = n77059 & ~n88074;
  assign n88076 = n85381 & ~n88041;
  assign n88077 = ~n88075 & ~n88076;
  assign n88078 = n85370 & ~n88041;
  assign n88079 = n85374 & ~n88041;
  assign n88080 = n77102 & ~n88041;
  assign n88081 = ~n88078 & ~n88079;
  assign n88082 = ~n88080 & n88081;
  assign n88083 = n88065 & n88070;
  assign n88084 = n88077 & n88083;
  assign n88085 = n88082 & n88084;
  assign n88086 = n88037 & ~n88042;
  assign n88087 = n88045 & n88086;
  assign n88088 = n88058 & n88087;
  assign n88089 = n88085 & n88088;
  assign n88090 = n85257 & ~n88089;
  assign n88091 = ~n88013 & ~n88014;
  assign n15686 = n88090 | ~n88091;
  assign n88093 = P2_P1_STATE2_REG_0_ & ~n76925;
  assign n88094 = ~P2_P1_STATE2_REG_0_ & ~n85224;
  assign n88095 = n77059 & n77062;
  assign n88096 = n77064 & n77068;
  assign n88097 = ~n88095 & ~n88096;
  assign n88098 = n77311 & ~n88097;
  assign n88099 = ~n88094 & ~n88098;
  assign n88100 = n88093 & ~n88099;
  assign n88101 = ~n85361 & n88100;
  assign n88102 = ~n85330 & n88101;
  assign n88103 = n85361 & n88100;
  assign n88104 = ~n85330 & n88103;
  assign n88105 = P2_P1_STATE2_REG_1_ & ~n88099;
  assign n88106 = P2_P1_STATEBS16_REG & n88105;
  assign n88107 = P2_P1_PHYADDRPOINTER_REG_0_ & n88106;
  assign n88108 = ~P2_P1_STATEBS16_REG & n88105;
  assign n88109 = P2_P1_PHYADDRPOINTER_REG_0_ & n88108;
  assign n88110 = P2_P1_PHYADDRPOINTER_REG_0_ & n88099;
  assign n88111 = P2_P1_STATE2_REG_0_ & n76925;
  assign n88112 = ~n88099 & n88111;
  assign n88113 = ~n85378 & n88112;
  assign n88114 = P2_P1_STATE2_REG_2_ & ~P2_P1_STATE2_REG_0_;
  assign n88115 = ~n88099 & n88114;
  assign n88116 = P2_P1_PHYADDRPOINTER_REG_0_ & n88115;
  assign n88117 = n77327 & ~n88099;
  assign n88118 = P2_P1_REIP_REG_0_ & n88117;
  assign n88119 = ~n88110 & ~n88113;
  assign n88120 = ~n88116 & n88119;
  assign n88121 = ~n88118 & n88120;
  assign n88122 = ~n88102 & ~n88104;
  assign n88123 = ~n88107 & n88122;
  assign n88124 = ~n88109 & n88123;
  assign n15691 = ~n88121 | ~n88124;
  assign n88126 = ~n85502 & n88101;
  assign n88127 = ~n85452 & n88103;
  assign n88128 = P2_P1_PHYADDRPOINTER_REG_1_ & n88106;
  assign n88129 = ~P2_P1_PHYADDRPOINTER_REG_1_ & n88108;
  assign n88130 = P2_P1_PHYADDRPOINTER_REG_1_ & n88099;
  assign n88131 = ~n85482 & n88112;
  assign n88132 = ~P2_P1_PHYADDRPOINTER_REG_1_ & n88115;
  assign n88133 = P2_P1_REIP_REG_1_ & n88117;
  assign n88134 = ~n88130 & ~n88131;
  assign n88135 = ~n88132 & n88134;
  assign n88136 = ~n88133 & n88135;
  assign n88137 = ~n88126 & ~n88127;
  assign n88138 = ~n88128 & n88137;
  assign n88139 = ~n88129 & n88138;
  assign n15696 = ~n88136 | ~n88139;
  assign n88141 = ~n85587 & n88101;
  assign n88142 = ~n85574 & n88103;
  assign n88143 = ~P2_P1_PHYADDRPOINTER_REG_2_ & n88106;
  assign n88144 = P2_P1_PHYADDRPOINTER_REG_1_ & ~P2_P1_PHYADDRPOINTER_REG_2_;
  assign n88145 = ~P2_P1_PHYADDRPOINTER_REG_1_ & P2_P1_PHYADDRPOINTER_REG_2_;
  assign n88146 = ~n88144 & ~n88145;
  assign n88147 = n88108 & ~n88146;
  assign n88148 = n88115 & ~n88146;
  assign n88149 = P2_P1_REIP_REG_2_ & n88117;
  assign n88150 = P2_P1_PHYADDRPOINTER_REG_2_ & n88099;
  assign n88151 = ~n85624 & n88112;
  assign n88152 = ~n88148 & ~n88149;
  assign n88153 = ~n88150 & n88152;
  assign n88154 = ~n88151 & n88153;
  assign n88155 = ~n88141 & ~n88142;
  assign n88156 = ~n88143 & n88155;
  assign n88157 = ~n88147 & n88156;
  assign n15701 = ~n88154 | ~n88157;
  assign n88159 = ~n85702 & n88101;
  assign n88160 = n85717 & n88103;
  assign n88161 = P2_P1_PHYADDRPOINTER_REG_2_ & ~P2_P1_PHYADDRPOINTER_REG_3_;
  assign n88162 = ~P2_P1_PHYADDRPOINTER_REG_2_ & P2_P1_PHYADDRPOINTER_REG_3_;
  assign n88163 = ~n88161 & ~n88162;
  assign n88164 = n88106 & ~n88163;
  assign n88165 = P2_P1_PHYADDRPOINTER_REG_1_ & P2_P1_PHYADDRPOINTER_REG_2_;
  assign n88166 = ~P2_P1_PHYADDRPOINTER_REG_3_ & n88165;
  assign n88167 = P2_P1_PHYADDRPOINTER_REG_3_ & ~n88165;
  assign n88168 = ~n88166 & ~n88167;
  assign n88169 = n88108 & ~n88168;
  assign n88170 = n88115 & ~n88168;
  assign n88171 = P2_P1_REIP_REG_3_ & n88117;
  assign n88172 = P2_P1_PHYADDRPOINTER_REG_3_ & n88099;
  assign n88173 = n85755 & n88112;
  assign n88174 = ~n88170 & ~n88171;
  assign n88175 = ~n88172 & n88174;
  assign n88176 = ~n88173 & n88175;
  assign n88177 = ~n88159 & ~n88160;
  assign n88178 = ~n88164 & n88177;
  assign n88179 = ~n88169 & n88178;
  assign n15706 = ~n88176 | ~n88179;
  assign n88181 = P2_P1_PHYADDRPOINTER_REG_2_ & P2_P1_PHYADDRPOINTER_REG_3_;
  assign n88182 = ~P2_P1_PHYADDRPOINTER_REG_4_ & n88181;
  assign n88183 = P2_P1_PHYADDRPOINTER_REG_4_ & ~n88181;
  assign n88184 = ~n88182 & ~n88183;
  assign n88185 = n88106 & ~n88184;
  assign n88186 = P2_P1_PHYADDRPOINTER_REG_3_ & n88165;
  assign n88187 = ~P2_P1_PHYADDRPOINTER_REG_4_ & n88186;
  assign n88188 = P2_P1_PHYADDRPOINTER_REG_4_ & ~n88186;
  assign n88189 = ~n88187 & ~n88188;
  assign n88190 = n88108 & ~n88189;
  assign n88191 = n85830 & n88103;
  assign n88192 = ~n85852 & n88101;
  assign n88193 = n88115 & ~n88189;
  assign n88194 = P2_P1_REIP_REG_4_ & n88117;
  assign n88195 = P2_P1_PHYADDRPOINTER_REG_4_ & n88099;
  assign n88196 = ~n85891 & n88112;
  assign n88197 = ~n88193 & ~n88194;
  assign n88198 = ~n88195 & n88197;
  assign n88199 = ~n88196 & n88198;
  assign n88200 = ~n88185 & ~n88190;
  assign n88201 = ~n88191 & n88200;
  assign n88202 = ~n88192 & n88201;
  assign n15711 = ~n88199 | ~n88202;
  assign n88204 = P2_P1_PHYADDRPOINTER_REG_4_ & n88181;
  assign n88205 = ~P2_P1_PHYADDRPOINTER_REG_5_ & n88204;
  assign n88206 = P2_P1_PHYADDRPOINTER_REG_5_ & ~n88204;
  assign n88207 = ~n88205 & ~n88206;
  assign n88208 = n88106 & ~n88207;
  assign n88209 = P2_P1_PHYADDRPOINTER_REG_4_ & n88186;
  assign n88210 = ~P2_P1_PHYADDRPOINTER_REG_5_ & n88209;
  assign n88211 = P2_P1_PHYADDRPOINTER_REG_5_ & ~n88209;
  assign n88212 = ~n88210 & ~n88211;
  assign n88213 = n88108 & ~n88212;
  assign n88214 = ~n85967 & n88101;
  assign n88215 = ~n85985 & n88103;
  assign n88216 = n88115 & ~n88212;
  assign n88217 = P2_P1_REIP_REG_5_ & n88117;
  assign n88218 = P2_P1_PHYADDRPOINTER_REG_5_ & n88099;
  assign n88219 = n86024 & n88112;
  assign n88220 = ~n88216 & ~n88217;
  assign n88221 = ~n88218 & n88220;
  assign n88222 = ~n88219 & n88221;
  assign n88223 = ~n88208 & ~n88213;
  assign n88224 = ~n88214 & n88223;
  assign n88225 = ~n88215 & n88224;
  assign n15716 = ~n88222 | ~n88225;
  assign n88227 = P2_P1_PHYADDRPOINTER_REG_5_ & n88204;
  assign n88228 = ~P2_P1_PHYADDRPOINTER_REG_6_ & n88227;
  assign n88229 = P2_P1_PHYADDRPOINTER_REG_6_ & ~n88227;
  assign n88230 = ~n88228 & ~n88229;
  assign n88231 = n88106 & ~n88230;
  assign n88232 = P2_P1_PHYADDRPOINTER_REG_5_ & n88209;
  assign n88233 = ~P2_P1_PHYADDRPOINTER_REG_6_ & n88232;
  assign n88234 = P2_P1_PHYADDRPOINTER_REG_6_ & ~n88232;
  assign n88235 = ~n88233 & ~n88234;
  assign n88236 = n88108 & ~n88235;
  assign n88237 = ~n86098 & n88101;
  assign n88238 = ~n86117 & n88103;
  assign n88239 = n88115 & ~n88235;
  assign n88240 = P2_P1_REIP_REG_6_ & n88117;
  assign n88241 = P2_P1_PHYADDRPOINTER_REG_6_ & n88099;
  assign n88242 = ~n86155 & n88112;
  assign n88243 = ~n88239 & ~n88240;
  assign n88244 = ~n88241 & n88243;
  assign n88245 = ~n88242 & n88244;
  assign n88246 = ~n88231 & ~n88236;
  assign n88247 = ~n88237 & n88246;
  assign n88248 = ~n88238 & n88247;
  assign n15721 = ~n88245 | ~n88248;
  assign n88250 = P2_P1_PHYADDRPOINTER_REG_6_ & n88227;
  assign n88251 = ~P2_P1_PHYADDRPOINTER_REG_7_ & n88250;
  assign n88252 = P2_P1_PHYADDRPOINTER_REG_7_ & ~n88250;
  assign n88253 = ~n88251 & ~n88252;
  assign n88254 = n88106 & ~n88253;
  assign n88255 = P2_P1_PHYADDRPOINTER_REG_6_ & n88232;
  assign n88256 = ~P2_P1_PHYADDRPOINTER_REG_7_ & n88255;
  assign n88257 = P2_P1_PHYADDRPOINTER_REG_7_ & ~n88255;
  assign n88258 = ~n88256 & ~n88257;
  assign n88259 = n88108 & ~n88258;
  assign n88260 = ~n86199 & n88101;
  assign n88261 = ~n86217 & n88103;
  assign n88262 = n88115 & ~n88258;
  assign n88263 = P2_P1_REIP_REG_7_ & n88117;
  assign n88264 = P2_P1_PHYADDRPOINTER_REG_7_ & n88099;
  assign n88265 = ~n86253 & n88112;
  assign n88266 = ~n88262 & ~n88263;
  assign n88267 = ~n88264 & n88266;
  assign n88268 = ~n88265 & n88267;
  assign n88269 = ~n88254 & ~n88259;
  assign n88270 = ~n88260 & n88269;
  assign n88271 = ~n88261 & n88270;
  assign n15726 = ~n88268 | ~n88271;
  assign n88273 = P2_P1_PHYADDRPOINTER_REG_7_ & n88250;
  assign n88274 = ~P2_P1_PHYADDRPOINTER_REG_8_ & n88273;
  assign n88275 = P2_P1_PHYADDRPOINTER_REG_8_ & ~n88273;
  assign n88276 = ~n88274 & ~n88275;
  assign n88277 = n88106 & ~n88276;
  assign n88278 = P2_P1_PHYADDRPOINTER_REG_7_ & n88255;
  assign n88279 = ~P2_P1_PHYADDRPOINTER_REG_8_ & n88278;
  assign n88280 = P2_P1_PHYADDRPOINTER_REG_8_ & ~n88278;
  assign n88281 = ~n88279 & ~n88280;
  assign n88282 = n88108 & ~n88281;
  assign n88283 = ~n86293 & n88101;
  assign n88284 = ~n86309 & n88103;
  assign n88285 = n88115 & ~n88281;
  assign n88286 = P2_P1_REIP_REG_8_ & n88117;
  assign n88287 = P2_P1_PHYADDRPOINTER_REG_8_ & n88099;
  assign n88288 = ~n86343 & n88112;
  assign n88289 = ~n88285 & ~n88286;
  assign n88290 = ~n88287 & n88289;
  assign n88291 = ~n88288 & n88290;
  assign n88292 = ~n88277 & ~n88282;
  assign n88293 = ~n88283 & n88292;
  assign n88294 = ~n88284 & n88293;
  assign n15731 = ~n88291 | ~n88294;
  assign n88296 = P2_P1_PHYADDRPOINTER_REG_8_ & n88273;
  assign n88297 = ~P2_P1_PHYADDRPOINTER_REG_9_ & n88296;
  assign n88298 = P2_P1_PHYADDRPOINTER_REG_9_ & ~n88296;
  assign n88299 = ~n88297 & ~n88298;
  assign n88300 = n88106 & ~n88299;
  assign n88301 = P2_P1_PHYADDRPOINTER_REG_8_ & n88278;
  assign n88302 = ~P2_P1_PHYADDRPOINTER_REG_9_ & n88301;
  assign n88303 = P2_P1_PHYADDRPOINTER_REG_9_ & ~n88301;
  assign n88304 = ~n88302 & ~n88303;
  assign n88305 = n88108 & ~n88304;
  assign n88306 = ~n86386 & n88101;
  assign n88307 = n86397 & n88103;
  assign n88308 = n88115 & ~n88304;
  assign n88309 = P2_P1_REIP_REG_9_ & n88117;
  assign n88310 = P2_P1_PHYADDRPOINTER_REG_9_ & n88099;
  assign n88311 = n86426 & n88112;
  assign n88312 = ~n88308 & ~n88309;
  assign n88313 = ~n88310 & n88312;
  assign n88314 = ~n88311 & n88313;
  assign n88315 = ~n88300 & ~n88305;
  assign n88316 = ~n88306 & n88315;
  assign n88317 = ~n88307 & n88316;
  assign n15736 = ~n88314 | ~n88317;
  assign n88319 = P2_P1_PHYADDRPOINTER_REG_9_ & n88296;
  assign n88320 = ~P2_P1_PHYADDRPOINTER_REG_10_ & n88319;
  assign n88321 = P2_P1_PHYADDRPOINTER_REG_10_ & ~n88319;
  assign n88322 = ~n88320 & ~n88321;
  assign n88323 = n88106 & ~n88322;
  assign n88324 = P2_P1_PHYADDRPOINTER_REG_9_ & n88301;
  assign n88325 = ~P2_P1_PHYADDRPOINTER_REG_10_ & n88324;
  assign n88326 = P2_P1_PHYADDRPOINTER_REG_10_ & ~n88324;
  assign n88327 = ~n88325 & ~n88326;
  assign n88328 = n88108 & ~n88327;
  assign n88329 = ~n86469 & n88101;
  assign n88330 = n86477 & n88103;
  assign n88331 = n88115 & ~n88327;
  assign n88332 = P2_P1_REIP_REG_10_ & n88117;
  assign n88333 = P2_P1_PHYADDRPOINTER_REG_10_ & n88099;
  assign n88334 = n86502 & n88112;
  assign n88335 = ~n88331 & ~n88332;
  assign n88336 = ~n88333 & n88335;
  assign n88337 = ~n88334 & n88336;
  assign n88338 = ~n88323 & ~n88328;
  assign n88339 = ~n88329 & n88338;
  assign n88340 = ~n88330 & n88339;
  assign n15741 = ~n88337 | ~n88340;
  assign n88342 = P2_P1_PHYADDRPOINTER_REG_10_ & n88319;
  assign n88343 = ~P2_P1_PHYADDRPOINTER_REG_11_ & n88342;
  assign n88344 = P2_P1_PHYADDRPOINTER_REG_11_ & ~n88342;
  assign n88345 = ~n88343 & ~n88344;
  assign n88346 = n88106 & ~n88345;
  assign n88347 = P2_P1_PHYADDRPOINTER_REG_10_ & n88324;
  assign n88348 = ~P2_P1_PHYADDRPOINTER_REG_11_ & n88347;
  assign n88349 = P2_P1_PHYADDRPOINTER_REG_11_ & ~n88347;
  assign n88350 = ~n88348 & ~n88349;
  assign n88351 = n88108 & ~n88350;
  assign n88352 = ~n86563 & n88101;
  assign n88353 = ~n86576 & n88103;
  assign n88354 = n88115 & ~n88350;
  assign n88355 = P2_P1_REIP_REG_11_ & n88117;
  assign n88356 = P2_P1_PHYADDRPOINTER_REG_11_ & n88099;
  assign n88357 = ~n86546 & n88112;
  assign n88358 = ~n88354 & ~n88355;
  assign n88359 = ~n88356 & n88358;
  assign n88360 = ~n88357 & n88359;
  assign n88361 = ~n88346 & ~n88351;
  assign n88362 = ~n88352 & n88361;
  assign n88363 = ~n88353 & n88362;
  assign n15746 = ~n88360 | ~n88363;
  assign n88365 = P2_P1_PHYADDRPOINTER_REG_11_ & n88342;
  assign n88366 = ~P2_P1_PHYADDRPOINTER_REG_12_ & n88365;
  assign n88367 = P2_P1_PHYADDRPOINTER_REG_12_ & ~n88365;
  assign n88368 = ~n88366 & ~n88367;
  assign n88369 = n88106 & ~n88368;
  assign n88370 = P2_P1_PHYADDRPOINTER_REG_11_ & n88347;
  assign n88371 = ~P2_P1_PHYADDRPOINTER_REG_12_ & n88370;
  assign n88372 = P2_P1_PHYADDRPOINTER_REG_12_ & ~n88370;
  assign n88373 = ~n88371 & ~n88372;
  assign n88374 = n88108 & ~n88373;
  assign n88375 = ~n86617 & n88101;
  assign n88376 = n86626 & n88103;
  assign n88377 = P2_P1_PHYADDRPOINTER_REG_12_ & n88099;
  assign n88378 = P2_P1_REIP_REG_12_ & n88117;
  assign n88379 = n88115 & ~n88373;
  assign n88380 = n86652 & n88112;
  assign n88381 = ~n88377 & ~n88378;
  assign n88382 = ~n88379 & n88381;
  assign n88383 = ~n88380 & n88382;
  assign n88384 = ~n88369 & ~n88374;
  assign n88385 = ~n88375 & n88384;
  assign n88386 = ~n88376 & n88385;
  assign n15751 = ~n88383 | ~n88386;
  assign n88388 = P2_P1_PHYADDRPOINTER_REG_12_ & n88365;
  assign n88389 = ~P2_P1_PHYADDRPOINTER_REG_13_ & n88388;
  assign n88390 = P2_P1_PHYADDRPOINTER_REG_13_ & ~n88388;
  assign n88391 = ~n88389 & ~n88390;
  assign n88392 = n88106 & ~n88391;
  assign n88393 = P2_P1_PHYADDRPOINTER_REG_12_ & n88370;
  assign n88394 = ~P2_P1_PHYADDRPOINTER_REG_13_ & n88393;
  assign n88395 = P2_P1_PHYADDRPOINTER_REG_13_ & ~n88393;
  assign n88396 = ~n88394 & ~n88395;
  assign n88397 = n88108 & ~n88396;
  assign n88398 = n86695 & n88101;
  assign n88399 = n86702 & n88103;
  assign n88400 = P2_P1_PHYADDRPOINTER_REG_13_ & n88099;
  assign n88401 = P2_P1_REIP_REG_13_ & n88117;
  assign n88402 = n88115 & ~n88396;
  assign n88403 = n86727 & n88112;
  assign n88404 = ~n88400 & ~n88401;
  assign n88405 = ~n88402 & n88404;
  assign n88406 = ~n88403 & n88405;
  assign n88407 = ~n88392 & ~n88397;
  assign n88408 = ~n88398 & n88407;
  assign n88409 = ~n88399 & n88408;
  assign n15756 = ~n88406 | ~n88409;
  assign n88411 = P2_P1_PHYADDRPOINTER_REG_13_ & n88388;
  assign n88412 = ~P2_P1_PHYADDRPOINTER_REG_14_ & n88411;
  assign n88413 = P2_P1_PHYADDRPOINTER_REG_14_ & ~n88411;
  assign n88414 = ~n88412 & ~n88413;
  assign n88415 = n88106 & ~n88414;
  assign n88416 = P2_P1_PHYADDRPOINTER_REG_13_ & n88393;
  assign n88417 = ~P2_P1_PHYADDRPOINTER_REG_14_ & n88416;
  assign n88418 = P2_P1_PHYADDRPOINTER_REG_14_ & ~n88416;
  assign n88419 = ~n88417 & ~n88418;
  assign n88420 = n88108 & ~n88419;
  assign n88421 = ~n86798 & n88101;
  assign n88422 = ~n86802 & n88103;
  assign n88423 = P2_P1_PHYADDRPOINTER_REG_14_ & n88099;
  assign n88424 = P2_P1_REIP_REG_14_ & n88117;
  assign n88425 = n88115 & ~n88419;
  assign n88426 = ~n86771 & n88112;
  assign n88427 = ~n88423 & ~n88424;
  assign n88428 = ~n88425 & n88427;
  assign n88429 = ~n88426 & n88428;
  assign n88430 = ~n88415 & ~n88420;
  assign n88431 = ~n88421 & n88430;
  assign n88432 = ~n88422 & n88431;
  assign n15761 = ~n88429 | ~n88432;
  assign n88434 = P2_P1_PHYADDRPOINTER_REG_14_ & n88411;
  assign n88435 = ~P2_P1_PHYADDRPOINTER_REG_15_ & n88434;
  assign n88436 = P2_P1_PHYADDRPOINTER_REG_15_ & ~n88434;
  assign n88437 = ~n88435 & ~n88436;
  assign n88438 = n88106 & ~n88437;
  assign n88439 = P2_P1_PHYADDRPOINTER_REG_14_ & n88416;
  assign n88440 = ~P2_P1_PHYADDRPOINTER_REG_15_ & n88439;
  assign n88441 = P2_P1_PHYADDRPOINTER_REG_15_ & ~n88439;
  assign n88442 = ~n88440 & ~n88441;
  assign n88443 = n88108 & ~n88442;
  assign n88444 = ~n86875 & n88101;
  assign n88445 = n86880 & n88103;
  assign n88446 = P2_P1_PHYADDRPOINTER_REG_15_ & n88099;
  assign n88447 = P2_P1_REIP_REG_15_ & n88117;
  assign n88448 = n88115 & ~n88442;
  assign n88449 = n86847 & n88112;
  assign n88450 = ~n88446 & ~n88447;
  assign n88451 = ~n88448 & n88450;
  assign n88452 = ~n88449 & n88451;
  assign n88453 = ~n88438 & ~n88443;
  assign n88454 = ~n88444 & n88453;
  assign n88455 = ~n88445 & n88454;
  assign n15766 = ~n88452 | ~n88455;
  assign n88457 = P2_P1_PHYADDRPOINTER_REG_15_ & n88434;
  assign n88458 = ~P2_P1_PHYADDRPOINTER_REG_16_ & n88457;
  assign n88459 = P2_P1_PHYADDRPOINTER_REG_16_ & ~n88457;
  assign n88460 = ~n88458 & ~n88459;
  assign n88461 = n88106 & ~n88460;
  assign n88462 = P2_P1_PHYADDRPOINTER_REG_15_ & n88439;
  assign n88463 = ~P2_P1_PHYADDRPOINTER_REG_16_ & n88462;
  assign n88464 = P2_P1_PHYADDRPOINTER_REG_16_ & ~n88462;
  assign n88465 = ~n88463 & ~n88464;
  assign n88466 = n88108 & ~n88465;
  assign n88467 = ~n86939 & n88101;
  assign n88468 = ~n86952 & n88103;
  assign n88469 = P2_P1_PHYADDRPOINTER_REG_16_ & n88099;
  assign n88470 = P2_P1_REIP_REG_16_ & n88117;
  assign n88471 = n88115 & ~n88465;
  assign n88472 = ~n86922 & n88112;
  assign n88473 = ~n88469 & ~n88470;
  assign n88474 = ~n88471 & n88473;
  assign n88475 = ~n88472 & n88474;
  assign n88476 = ~n88461 & ~n88466;
  assign n88477 = ~n88467 & n88476;
  assign n88478 = ~n88468 & n88477;
  assign n15771 = ~n88475 | ~n88478;
  assign n88480 = P2_P1_PHYADDRPOINTER_REG_16_ & n88457;
  assign n88481 = ~P2_P1_PHYADDRPOINTER_REG_17_ & n88480;
  assign n88482 = P2_P1_PHYADDRPOINTER_REG_17_ & ~n88480;
  assign n88483 = ~n88481 & ~n88482;
  assign n88484 = n88106 & ~n88483;
  assign n88485 = P2_P1_PHYADDRPOINTER_REG_16_ & n88462;
  assign n88486 = ~P2_P1_PHYADDRPOINTER_REG_17_ & n88485;
  assign n88487 = P2_P1_PHYADDRPOINTER_REG_17_ & ~n88485;
  assign n88488 = ~n88486 & ~n88487;
  assign n88489 = n88108 & ~n88488;
  assign n88490 = n86995 & n88101;
  assign n88491 = n87003 & n88103;
  assign n88492 = P2_P1_PHYADDRPOINTER_REG_17_ & n88099;
  assign n88493 = P2_P1_REIP_REG_17_ & n88117;
  assign n88494 = n88115 & ~n88488;
  assign n88495 = n87029 & n88112;
  assign n88496 = ~n88492 & ~n88493;
  assign n88497 = ~n88494 & n88496;
  assign n88498 = ~n88495 & n88497;
  assign n88499 = ~n88484 & ~n88489;
  assign n88500 = ~n88490 & n88499;
  assign n88501 = ~n88491 & n88500;
  assign n15776 = ~n88498 | ~n88501;
  assign n88503 = P2_P1_PHYADDRPOINTER_REG_17_ & n88480;
  assign n88504 = ~P2_P1_PHYADDRPOINTER_REG_18_ & n88503;
  assign n88505 = P2_P1_PHYADDRPOINTER_REG_18_ & ~n88503;
  assign n88506 = ~n88504 & ~n88505;
  assign n88507 = n88106 & ~n88506;
  assign n88508 = P2_P1_PHYADDRPOINTER_REG_17_ & n88485;
  assign n88509 = ~P2_P1_PHYADDRPOINTER_REG_18_ & n88508;
  assign n88510 = P2_P1_PHYADDRPOINTER_REG_18_ & ~n88508;
  assign n88511 = ~n88509 & ~n88510;
  assign n88512 = n88108 & ~n88511;
  assign n88513 = ~n87089 & n88101;
  assign n88514 = ~n87102 & n88103;
  assign n88515 = P2_P1_PHYADDRPOINTER_REG_18_ & n88099;
  assign n88516 = P2_P1_REIP_REG_18_ & n88117;
  assign n88517 = n88115 & ~n88511;
  assign n88518 = ~n87073 & n88112;
  assign n88519 = ~n88515 & ~n88516;
  assign n88520 = ~n88517 & n88519;
  assign n88521 = ~n88518 & n88520;
  assign n88522 = ~n88507 & ~n88512;
  assign n88523 = ~n88513 & n88522;
  assign n88524 = ~n88514 & n88523;
  assign n15781 = ~n88521 | ~n88524;
  assign n88526 = P2_P1_PHYADDRPOINTER_REG_18_ & n88503;
  assign n88527 = ~P2_P1_PHYADDRPOINTER_REG_19_ & n88526;
  assign n88528 = P2_P1_PHYADDRPOINTER_REG_19_ & ~n88526;
  assign n88529 = ~n88527 & ~n88528;
  assign n88530 = n88106 & ~n88529;
  assign n88531 = P2_P1_PHYADDRPOINTER_REG_18_ & n88508;
  assign n88532 = ~P2_P1_PHYADDRPOINTER_REG_19_ & n88531;
  assign n88533 = P2_P1_PHYADDRPOINTER_REG_19_ & ~n88531;
  assign n88534 = ~n88532 & ~n88533;
  assign n88535 = n88108 & ~n88534;
  assign n88536 = ~n87143 & n88101;
  assign n88537 = n87152 & n88103;
  assign n88538 = P2_P1_PHYADDRPOINTER_REG_19_ & n88099;
  assign n88539 = P2_P1_REIP_REG_19_ & n88117;
  assign n88540 = n88115 & ~n88534;
  assign n88541 = n87178 & n88112;
  assign n88542 = ~n88538 & ~n88539;
  assign n88543 = ~n88540 & n88542;
  assign n88544 = ~n88541 & n88543;
  assign n88545 = ~n88530 & ~n88535;
  assign n88546 = ~n88536 & n88545;
  assign n88547 = ~n88537 & n88546;
  assign n15786 = ~n88544 | ~n88547;
  assign n88549 = P2_P1_PHYADDRPOINTER_REG_19_ & n88526;
  assign n88550 = ~P2_P1_PHYADDRPOINTER_REG_20_ & n88549;
  assign n88551 = P2_P1_PHYADDRPOINTER_REG_20_ & ~n88549;
  assign n88552 = ~n88550 & ~n88551;
  assign n88553 = n88106 & ~n88552;
  assign n88554 = P2_P1_PHYADDRPOINTER_REG_19_ & n88531;
  assign n88555 = ~P2_P1_PHYADDRPOINTER_REG_20_ & n88554;
  assign n88556 = P2_P1_PHYADDRPOINTER_REG_20_ & ~n88554;
  assign n88557 = ~n88555 & ~n88556;
  assign n88558 = n88108 & ~n88557;
  assign n88559 = n87230 & n88103;
  assign n88560 = P2_P1_PHYADDRPOINTER_REG_20_ & n88099;
  assign n88561 = P2_P1_REIP_REG_20_ & n88117;
  assign n88562 = n88115 & ~n88557;
  assign n88563 = n87254 & n88112;
  assign n88564 = ~n88560 & ~n88561;
  assign n88565 = ~n88562 & n88564;
  assign n88566 = ~n88563 & n88565;
  assign n88567 = n87205 & n88101;
  assign n88568 = ~n88553 & ~n88558;
  assign n88569 = ~n88559 & n88568;
  assign n88570 = n88566 & n88569;
  assign n15791 = n88567 | ~n88570;
  assign n88572 = P2_P1_PHYADDRPOINTER_REG_20_ & n88549;
  assign n88573 = ~P2_P1_PHYADDRPOINTER_REG_21_ & n88572;
  assign n88574 = P2_P1_PHYADDRPOINTER_REG_21_ & ~n88572;
  assign n88575 = ~n88573 & ~n88574;
  assign n88576 = n88106 & ~n88575;
  assign n88577 = P2_P1_PHYADDRPOINTER_REG_20_ & n88554;
  assign n88578 = ~P2_P1_PHYADDRPOINTER_REG_21_ & n88577;
  assign n88579 = P2_P1_PHYADDRPOINTER_REG_21_ & ~n88577;
  assign n88580 = ~n88578 & ~n88579;
  assign n88581 = n88108 & ~n88580;
  assign n88582 = n87287 & n88103;
  assign n88583 = P2_P1_PHYADDRPOINTER_REG_21_ & n88099;
  assign n88584 = P2_P1_REIP_REG_21_ & n88117;
  assign n88585 = n88115 & ~n88580;
  assign n88586 = n87312 & n88112;
  assign n88587 = ~n88583 & ~n88584;
  assign n88588 = ~n88585 & n88587;
  assign n88589 = ~n88586 & n88588;
  assign n88590 = ~n87328 & n88101;
  assign n88591 = ~n88576 & ~n88581;
  assign n88592 = ~n88582 & n88591;
  assign n88593 = n88589 & n88592;
  assign n15796 = n88590 | ~n88593;
  assign n88595 = P2_P1_PHYADDRPOINTER_REG_21_ & n88572;
  assign n88596 = ~P2_P1_PHYADDRPOINTER_REG_22_ & n88595;
  assign n88597 = P2_P1_PHYADDRPOINTER_REG_22_ & ~n88595;
  assign n88598 = ~n88596 & ~n88597;
  assign n88599 = n88106 & ~n88598;
  assign n88600 = ~n87389 & n88101;
  assign n88601 = P2_P1_PHYADDRPOINTER_REG_21_ & n88577;
  assign n88602 = ~P2_P1_PHYADDRPOINTER_REG_22_ & n88601;
  assign n88603 = P2_P1_PHYADDRPOINTER_REG_22_ & ~n88601;
  assign n88604 = ~n88602 & ~n88603;
  assign n88605 = n88108 & ~n88604;
  assign n88606 = ~n87406 & n88103;
  assign n88607 = P2_P1_PHYADDRPOINTER_REG_22_ & n88099;
  assign n88608 = P2_P1_REIP_REG_22_ & n88117;
  assign n88609 = n88115 & ~n88604;
  assign n88610 = ~n87368 & n88112;
  assign n88611 = ~n88607 & ~n88608;
  assign n88612 = ~n88609 & n88611;
  assign n88613 = ~n88610 & n88612;
  assign n88614 = ~n88599 & ~n88600;
  assign n88615 = ~n88605 & n88614;
  assign n88616 = ~n88606 & n88615;
  assign n15801 = ~n88613 | ~n88616;
  assign n88618 = P2_P1_PHYADDRPOINTER_REG_22_ & n88595;
  assign n88619 = ~P2_P1_PHYADDRPOINTER_REG_23_ & n88618;
  assign n88620 = P2_P1_PHYADDRPOINTER_REG_23_ & ~n88618;
  assign n88621 = ~n88619 & ~n88620;
  assign n88622 = n88106 & ~n88621;
  assign n88623 = ~n87465 & n88101;
  assign n88624 = P2_P1_PHYADDRPOINTER_REG_22_ & n88601;
  assign n88625 = ~P2_P1_PHYADDRPOINTER_REG_23_ & n88624;
  assign n88626 = P2_P1_PHYADDRPOINTER_REG_23_ & ~n88624;
  assign n88627 = ~n88625 & ~n88626;
  assign n88628 = n88108 & ~n88627;
  assign n88629 = n87483 & n88103;
  assign n88630 = P2_P1_PHYADDRPOINTER_REG_23_ & n88099;
  assign n88631 = P2_P1_REIP_REG_23_ & n88117;
  assign n88632 = n88115 & ~n88627;
  assign n88633 = n87447 & n88112;
  assign n88634 = ~n88630 & ~n88631;
  assign n88635 = ~n88632 & n88634;
  assign n88636 = ~n88633 & n88635;
  assign n88637 = ~n88622 & ~n88623;
  assign n88638 = ~n88628 & n88637;
  assign n88639 = ~n88629 & n88638;
  assign n15806 = ~n88636 | ~n88639;
  assign n88641 = P2_P1_PHYADDRPOINTER_REG_23_ & n88618;
  assign n88642 = ~P2_P1_PHYADDRPOINTER_REG_24_ & n88641;
  assign n88643 = P2_P1_PHYADDRPOINTER_REG_24_ & ~n88641;
  assign n88644 = ~n88642 & ~n88643;
  assign n88645 = n88106 & ~n88644;
  assign n88646 = ~n87540 & n88101;
  assign n88647 = P2_P1_PHYADDRPOINTER_REG_23_ & n88624;
  assign n88648 = ~P2_P1_PHYADDRPOINTER_REG_24_ & n88647;
  assign n88649 = P2_P1_PHYADDRPOINTER_REG_24_ & ~n88647;
  assign n88650 = ~n88648 & ~n88649;
  assign n88651 = n88108 & ~n88650;
  assign n88652 = ~n87548 & n88103;
  assign n88653 = P2_P1_PHYADDRPOINTER_REG_24_ & n88099;
  assign n88654 = P2_P1_REIP_REG_24_ & n88117;
  assign n88655 = n88115 & ~n88650;
  assign n88656 = ~n87513 & n88112;
  assign n88657 = ~n88653 & ~n88654;
  assign n88658 = ~n88655 & n88657;
  assign n88659 = ~n88656 & n88658;
  assign n88660 = ~n88645 & ~n88646;
  assign n88661 = ~n88651 & n88660;
  assign n88662 = ~n88652 & n88661;
  assign n15811 = ~n88659 | ~n88662;
  assign n88664 = P2_P1_PHYADDRPOINTER_REG_24_ & n88641;
  assign n88665 = ~P2_P1_PHYADDRPOINTER_REG_25_ & n88664;
  assign n88666 = P2_P1_PHYADDRPOINTER_REG_25_ & ~n88664;
  assign n88667 = ~n88665 & ~n88666;
  assign n88668 = n88106 & ~n88667;
  assign n88669 = ~n87617 & n88101;
  assign n88670 = P2_P1_PHYADDRPOINTER_REG_24_ & n88647;
  assign n88671 = ~P2_P1_PHYADDRPOINTER_REG_25_ & n88670;
  assign n88672 = P2_P1_PHYADDRPOINTER_REG_25_ & ~n88670;
  assign n88673 = ~n88671 & ~n88672;
  assign n88674 = n88108 & ~n88673;
  assign n88675 = n87623 & n88103;
  assign n88676 = P2_P1_PHYADDRPOINTER_REG_25_ & n88099;
  assign n88677 = P2_P1_REIP_REG_25_ & n88117;
  assign n88678 = n88115 & ~n88673;
  assign n88679 = n87589 & n88112;
  assign n88680 = ~n88676 & ~n88677;
  assign n88681 = ~n88678 & n88680;
  assign n88682 = ~n88679 & n88681;
  assign n88683 = ~n88668 & ~n88669;
  assign n88684 = ~n88674 & n88683;
  assign n88685 = ~n88675 & n88684;
  assign n15816 = ~n88682 | ~n88685;
  assign n88687 = P2_P1_PHYADDRPOINTER_REG_25_ & n88664;
  assign n88688 = ~P2_P1_PHYADDRPOINTER_REG_26_ & n88687;
  assign n88689 = P2_P1_PHYADDRPOINTER_REG_26_ & ~n88687;
  assign n88690 = ~n88688 & ~n88689;
  assign n88691 = n88106 & ~n88690;
  assign n88692 = n87658 & n88101;
  assign n88693 = P2_P1_PHYADDRPOINTER_REG_25_ & n88670;
  assign n88694 = ~P2_P1_PHYADDRPOINTER_REG_26_ & n88693;
  assign n88695 = P2_P1_PHYADDRPOINTER_REG_26_ & ~n88693;
  assign n88696 = ~n88694 & ~n88695;
  assign n88697 = n88108 & ~n88696;
  assign n88698 = n87662 & n88103;
  assign n88699 = P2_P1_PHYADDRPOINTER_REG_26_ & n88099;
  assign n88700 = n87700 & n88112;
  assign n88701 = n88115 & ~n88696;
  assign n88702 = P2_P1_REIP_REG_26_ & n88117;
  assign n88703 = ~n88699 & ~n88700;
  assign n88704 = ~n88701 & n88703;
  assign n88705 = ~n88702 & n88704;
  assign n88706 = ~n88691 & ~n88692;
  assign n88707 = ~n88697 & n88706;
  assign n88708 = ~n88698 & n88707;
  assign n15821 = ~n88705 | ~n88708;
  assign n88710 = P2_P1_PHYADDRPOINTER_REG_26_ & n88687;
  assign n88711 = ~P2_P1_PHYADDRPOINTER_REG_27_ & n88710;
  assign n88712 = P2_P1_PHYADDRPOINTER_REG_27_ & ~n88710;
  assign n88713 = ~n88711 & ~n88712;
  assign n88714 = n88106 & ~n88713;
  assign n88715 = ~n87729 & n88101;
  assign n88716 = P2_P1_PHYADDRPOINTER_REG_26_ & n88693;
  assign n88717 = ~P2_P1_PHYADDRPOINTER_REG_27_ & n88716;
  assign n88718 = P2_P1_PHYADDRPOINTER_REG_27_ & ~n88716;
  assign n88719 = ~n88717 & ~n88718;
  assign n88720 = n88108 & ~n88719;
  assign n88721 = ~n87733 & n88103;
  assign n88722 = P2_P1_PHYADDRPOINTER_REG_27_ & n88099;
  assign n88723 = ~n87771 & n88112;
  assign n88724 = n88115 & ~n88719;
  assign n88725 = P2_P1_REIP_REG_27_ & n88117;
  assign n88726 = ~n88722 & ~n88723;
  assign n88727 = ~n88724 & n88726;
  assign n88728 = ~n88725 & n88727;
  assign n88729 = ~n88714 & ~n88715;
  assign n88730 = ~n88720 & n88729;
  assign n88731 = ~n88721 & n88730;
  assign n15826 = ~n88728 | ~n88731;
  assign n88733 = n87807 & n88101;
  assign n88734 = n87812 & n88103;
  assign n88735 = P2_P1_PHYADDRPOINTER_REG_27_ & n88710;
  assign n88736 = ~P2_P1_PHYADDRPOINTER_REG_28_ & n88735;
  assign n88737 = P2_P1_PHYADDRPOINTER_REG_28_ & ~n88735;
  assign n88738 = ~n88736 & ~n88737;
  assign n88739 = n88106 & ~n88738;
  assign n88740 = P2_P1_PHYADDRPOINTER_REG_27_ & n88716;
  assign n88741 = ~P2_P1_PHYADDRPOINTER_REG_28_ & n88740;
  assign n88742 = P2_P1_PHYADDRPOINTER_REG_28_ & ~n88740;
  assign n88743 = ~n88741 & ~n88742;
  assign n88744 = n88108 & ~n88743;
  assign n88745 = P2_P1_PHYADDRPOINTER_REG_28_ & n88099;
  assign n88746 = n87851 & n88112;
  assign n88747 = n88115 & ~n88743;
  assign n88748 = P2_P1_REIP_REG_28_ & n88117;
  assign n88749 = ~n88745 & ~n88746;
  assign n88750 = ~n88747 & n88749;
  assign n88751 = ~n88748 & n88750;
  assign n88752 = ~n88733 & ~n88734;
  assign n88753 = ~n88739 & n88752;
  assign n88754 = ~n88744 & n88753;
  assign n15831 = ~n88751 | ~n88754;
  assign n88756 = ~n87880 & n88101;
  assign n88757 = n87884 & n88103;
  assign n88758 = P2_P1_PHYADDRPOINTER_REG_28_ & n88735;
  assign n88759 = ~P2_P1_PHYADDRPOINTER_REG_29_ & n88758;
  assign n88760 = P2_P1_PHYADDRPOINTER_REG_29_ & ~n88758;
  assign n88761 = ~n88759 & ~n88760;
  assign n88762 = n88106 & ~n88761;
  assign n88763 = P2_P1_PHYADDRPOINTER_REG_28_ & n88740;
  assign n88764 = ~P2_P1_PHYADDRPOINTER_REG_29_ & n88763;
  assign n88765 = P2_P1_PHYADDRPOINTER_REG_29_ & ~n88763;
  assign n88766 = ~n88764 & ~n88765;
  assign n88767 = n88108 & ~n88766;
  assign n88768 = P2_P1_PHYADDRPOINTER_REG_29_ & n88099;
  assign n88769 = P2_P1_REIP_REG_29_ & n88117;
  assign n88770 = n87922 & n88112;
  assign n88771 = n88115 & ~n88766;
  assign n88772 = ~n88768 & ~n88769;
  assign n88773 = ~n88770 & n88772;
  assign n88774 = ~n88771 & n88773;
  assign n88775 = ~n88756 & ~n88757;
  assign n88776 = ~n88762 & n88775;
  assign n88777 = ~n88767 & n88776;
  assign n15836 = ~n88774 | ~n88777;
  assign n88779 = ~n87952 & n88101;
  assign n88780 = ~n87956 & n88103;
  assign n88781 = P2_P1_PHYADDRPOINTER_REG_29_ & n88758;
  assign n88782 = ~P2_P1_PHYADDRPOINTER_REG_30_ & n88781;
  assign n88783 = P2_P1_PHYADDRPOINTER_REG_30_ & ~n88781;
  assign n88784 = ~n88782 & ~n88783;
  assign n88785 = n88106 & ~n88784;
  assign n88786 = P2_P1_PHYADDRPOINTER_REG_29_ & n88763;
  assign n88787 = ~P2_P1_PHYADDRPOINTER_REG_30_ & n88786;
  assign n88788 = P2_P1_PHYADDRPOINTER_REG_30_ & ~n88786;
  assign n88789 = ~n88787 & ~n88788;
  assign n88790 = n88108 & ~n88789;
  assign n88791 = P2_P1_PHYADDRPOINTER_REG_30_ & n88099;
  assign n88792 = P2_P1_REIP_REG_30_ & n88117;
  assign n88793 = ~n87994 & n88112;
  assign n88794 = n88115 & ~n88789;
  assign n88795 = ~n88791 & ~n88792;
  assign n88796 = ~n88793 & n88795;
  assign n88797 = ~n88794 & n88796;
  assign n88798 = ~n88779 & ~n88780;
  assign n88799 = ~n88785 & n88798;
  assign n88800 = ~n88790 & n88799;
  assign n15841 = ~n88797 | ~n88800;
  assign n88802 = n88030 & n88101;
  assign n88803 = P2_P1_PHYADDRPOINTER_REG_30_ & n88781;
  assign n88804 = ~P2_P1_PHYADDRPOINTER_REG_31_ & n88803;
  assign n88805 = P2_P1_PHYADDRPOINTER_REG_31_ & ~n88803;
  assign n88806 = ~n88804 & ~n88805;
  assign n88807 = n88106 & ~n88806;
  assign n88808 = ~n88035 & n88103;
  assign n88809 = P2_P1_PHYADDRPOINTER_REG_30_ & n88786;
  assign n88810 = ~P2_P1_PHYADDRPOINTER_REG_31_ & n88809;
  assign n88811 = P2_P1_PHYADDRPOINTER_REG_31_ & ~n88809;
  assign n88812 = ~n88810 & ~n88811;
  assign n88813 = n88108 & ~n88812;
  assign n88814 = P2_P1_PHYADDRPOINTER_REG_31_ & n88099;
  assign n88815 = P2_P1_REIP_REG_31_ & n88117;
  assign n88816 = ~n88074 & n88112;
  assign n88817 = n88115 & ~n88812;
  assign n88818 = ~n88814 & ~n88815;
  assign n88819 = ~n88816 & n88818;
  assign n88820 = ~n88817 & n88819;
  assign n88821 = ~n88802 & ~n88807;
  assign n88822 = ~n88808 & n88821;
  assign n88823 = ~n88813 & n88822;
  assign n15846 = ~n88820 | ~n88823;
  assign n88825 = ~n76584 & n77040;
  assign n88826 = n77009 & n88825;
  assign n88827 = ~n77196 & ~n88826;
  assign n88828 = n77311 & ~n88827;
  assign n88829 = P2_P1_LWORD_REG_15_ & ~n88828;
  assign n88830 = n76925 & n88828;
  assign n88831 = P2_P1_EAX_REG_15_ & n88830;
  assign n88832 = P2_BUF1_REG_15_ & n12802;
  assign n88833 = ~n80442 & ~n80446;
  assign n88834 = n80442 & n80446;
  assign n88835 = ~n88833 & ~n88834;
  assign n88836 = n80532 & ~n88835;
  assign n88837 = ~n80447 & ~n80448;
  assign n88838 = ~n80532 & ~n88837;
  assign n88839 = ~n88836 & ~n88838;
  assign n88840 = ~n12802 & ~n88839;
  assign n88841 = ~n88832 & ~n88840;
  assign n88842 = ~n76925 & n88828;
  assign n88843 = ~n88841 & n88842;
  assign n88844 = ~n88829 & ~n88831;
  assign n15851 = n88843 | ~n88844;
  assign n88846 = P2_P1_LWORD_REG_14_ & ~n88828;
  assign n88847 = P2_P1_EAX_REG_14_ & n88830;
  assign n88848 = P2_BUF1_REG_14_ & n12802;
  assign n88849 = n80457 & ~n80530;
  assign n88850 = ~n80457 & n80530;
  assign n88851 = ~n88849 & ~n88850;
  assign n88852 = ~n80456 & n88851;
  assign n88853 = n80456 & n88850;
  assign n88854 = n80458 & ~n80530;
  assign n88855 = ~n88852 & ~n88853;
  assign n88856 = ~n88854 & n88855;
  assign n88857 = ~n12802 & ~n88856;
  assign n88858 = ~n88848 & ~n88857;
  assign n88859 = n88842 & ~n88858;
  assign n88860 = ~n88846 & ~n88847;
  assign n15856 = n88859 | ~n88860;
  assign n88862 = P2_P1_LWORD_REG_13_ & ~n88828;
  assign n88863 = P2_P1_EAX_REG_13_ & n88830;
  assign n88864 = P2_BUF1_REG_13_ & n12802;
  assign n88865 = ~n80460 & ~n80467;
  assign n88866 = n80460 & n80467;
  assign n88867 = ~n88865 & ~n88866;
  assign n88868 = n80528 & ~n88867;
  assign n88869 = ~n80528 & n88867;
  assign n88870 = ~n88868 & ~n88869;
  assign n88871 = ~n12802 & ~n88870;
  assign n88872 = ~n88864 & ~n88871;
  assign n88873 = n88842 & ~n88872;
  assign n88874 = ~n88862 & ~n88863;
  assign n15861 = n88873 | ~n88874;
  assign n88876 = P2_P1_LWORD_REG_12_ & ~n88828;
  assign n88877 = P2_P1_EAX_REG_12_ & n88830;
  assign n88878 = P2_BUF1_REG_12_ & n12802;
  assign n88879 = ~n80470 & n80526;
  assign n88880 = n80476 & n88879;
  assign n88881 = n80470 & ~n80526;
  assign n88882 = ~n88879 & ~n88881;
  assign n88883 = ~n80476 & n88882;
  assign n88884 = n80477 & ~n80526;
  assign n88885 = ~n88880 & ~n88883;
  assign n88886 = ~n88884 & n88885;
  assign n88887 = ~n12802 & ~n88886;
  assign n88888 = ~n88878 & ~n88887;
  assign n88889 = n88842 & ~n88888;
  assign n88890 = ~n88876 & ~n88877;
  assign n15866 = n88889 | ~n88890;
  assign n88892 = P2_P1_LWORD_REG_11_ & ~n88828;
  assign n88893 = P2_P1_EAX_REG_11_ & n88830;
  assign n88894 = P2_BUF1_REG_11_ & n12802;
  assign n88895 = ~n80479 & ~n80483;
  assign n88896 = n80479 & n80483;
  assign n88897 = ~n88895 & ~n88896;
  assign n88898 = n80524 & ~n88897;
  assign n88899 = ~n80484 & ~n80485;
  assign n88900 = ~n80524 & ~n88899;
  assign n88901 = ~n88898 & ~n88900;
  assign n88902 = ~n12802 & ~n88901;
  assign n88903 = ~n88894 & ~n88902;
  assign n88904 = n88842 & ~n88903;
  assign n88905 = ~n88892 & ~n88893;
  assign n15871 = n88904 | ~n88905;
  assign n88907 = P2_P1_LWORD_REG_10_ & ~n88828;
  assign n88908 = P2_P1_EAX_REG_10_ & n88830;
  assign n88909 = P2_BUF1_REG_10_ & n12802;
  assign n88910 = n80494 & ~n80522;
  assign n88911 = ~n80494 & n80522;
  assign n88912 = ~n88910 & ~n88911;
  assign n88913 = ~n80493 & n88912;
  assign n88914 = n80493 & n88911;
  assign n88915 = ~n88913 & ~n88914;
  assign n88916 = n80495 & ~n80522;
  assign n88917 = n88915 & ~n88916;
  assign n88918 = ~n12802 & ~n88917;
  assign n88919 = ~n88909 & ~n88918;
  assign n88920 = n88842 & ~n88919;
  assign n88921 = ~n88907 & ~n88908;
  assign n15876 = n88920 | ~n88921;
  assign n88923 = P2_P1_LWORD_REG_9_ & ~n88828;
  assign n88924 = P2_P1_EAX_REG_9_ & n88830;
  assign n88925 = P2_BUF1_REG_9_ & n12802;
  assign n88926 = ~n80506 & ~n80507;
  assign n88927 = n80520 & n88926;
  assign n88928 = ~n80520 & ~n88926;
  assign n88929 = ~n88927 & ~n88928;
  assign n88930 = ~n12802 & ~n88929;
  assign n88931 = ~n88925 & ~n88930;
  assign n88932 = n88842 & ~n88931;
  assign n88933 = ~n88923 & ~n88924;
  assign n15881 = n88932 | ~n88933;
  assign n88935 = P2_P1_LWORD_REG_8_ & ~n88828;
  assign n88936 = P2_P1_EAX_REG_8_ & n88830;
  assign n88937 = P2_BUF1_REG_8_ & n12802;
  assign n88938 = ~n80508 & ~n80517;
  assign n88939 = n80508 & n80517;
  assign n88940 = ~n88938 & ~n88939;
  assign n88941 = n80510 & ~n88940;
  assign n88942 = ~n80508 & n80517;
  assign n88943 = ~n80510 & n88942;
  assign n88944 = n80511 & ~n80517;
  assign n88945 = ~n88941 & ~n88943;
  assign n88946 = ~n88944 & n88945;
  assign n88947 = ~n12802 & ~n88946;
  assign n88948 = ~n88937 & ~n88947;
  assign n88949 = n88842 & ~n88948;
  assign n88950 = ~n88935 & ~n88936;
  assign n15886 = n88949 | ~n88950;
  assign n88952 = P2_P1_LWORD_REG_7_ & ~n88828;
  assign n88953 = P2_P1_EAX_REG_7_ & n88830;
  assign n88954 = ~n77700 & n88842;
  assign n88955 = ~n88952 & ~n88953;
  assign n15891 = n88954 | ~n88955;
  assign n88957 = P2_P1_LWORD_REG_6_ & ~n88828;
  assign n88958 = P2_P1_EAX_REG_6_ & n88830;
  assign n88959 = ~n83535 & n88842;
  assign n88960 = ~n88957 & ~n88958;
  assign n15896 = n88959 | ~n88960;
  assign n88962 = P2_P1_LWORD_REG_5_ & ~n88828;
  assign n88963 = P2_P1_EAX_REG_5_ & n88830;
  assign n88964 = ~n83582 & n88842;
  assign n88965 = ~n88962 & ~n88963;
  assign n15901 = n88964 | ~n88965;
  assign n88967 = ~n83626 & n88842;
  assign n88968 = P2_P1_EAX_REG_4_ & n88830;
  assign n88969 = P2_P1_LWORD_REG_4_ & ~n88828;
  assign n88970 = ~n88967 & ~n88968;
  assign n15906 = n88969 | ~n88970;
  assign n88972 = ~n83670 & n88842;
  assign n88973 = P2_P1_EAX_REG_3_ & n88830;
  assign n88974 = P2_P1_LWORD_REG_3_ & ~n88828;
  assign n88975 = ~n88972 & ~n88973;
  assign n15911 = n88974 | ~n88975;
  assign n88977 = ~n83712 & n88842;
  assign n88978 = P2_P1_EAX_REG_2_ & n88830;
  assign n88979 = P2_P1_LWORD_REG_2_ & ~n88828;
  assign n88980 = ~n88977 & ~n88978;
  assign n15916 = n88979 | ~n88980;
  assign n88982 = ~n83757 & n88842;
  assign n88983 = P2_P1_EAX_REG_1_ & n88830;
  assign n88984 = P2_P1_LWORD_REG_1_ & ~n88828;
  assign n88985 = ~n88982 & ~n88983;
  assign n15921 = n88984 | ~n88985;
  assign n88987 = ~n83790 & n88842;
  assign n88988 = P2_P1_EAX_REG_0_ & n88830;
  assign n88989 = P2_P1_LWORD_REG_0_ & ~n88828;
  assign n88990 = ~n88987 & ~n88988;
  assign n15926 = n88989 | ~n88990;
  assign n88992 = P2_P1_UWORD_REG_14_ & ~n88828;
  assign n88993 = P2_P1_EAX_REG_30_ & n88830;
  assign n88994 = ~n88992 & ~n88993;
  assign n15931 = n88859 | ~n88994;
  assign n88996 = P2_P1_UWORD_REG_13_ & ~n88828;
  assign n88997 = P2_P1_EAX_REG_29_ & n88830;
  assign n88998 = ~n88996 & ~n88997;
  assign n15936 = n88873 | ~n88998;
  assign n89000 = P2_P1_UWORD_REG_12_ & ~n88828;
  assign n89001 = P2_P1_EAX_REG_28_ & n88830;
  assign n89002 = ~n89000 & ~n89001;
  assign n15941 = n88889 | ~n89002;
  assign n89004 = P2_P1_UWORD_REG_11_ & ~n88828;
  assign n89005 = P2_P1_EAX_REG_27_ & n88830;
  assign n89006 = ~n89004 & ~n89005;
  assign n15946 = n88904 | ~n89006;
  assign n89008 = P2_P1_UWORD_REG_10_ & ~n88828;
  assign n89009 = P2_P1_EAX_REG_26_ & n88830;
  assign n89010 = ~n89008 & ~n89009;
  assign n15951 = n88920 | ~n89010;
  assign n89012 = P2_P1_UWORD_REG_9_ & ~n88828;
  assign n89013 = P2_P1_EAX_REG_25_ & n88830;
  assign n89014 = ~n89012 & ~n89013;
  assign n15956 = n88932 | ~n89014;
  assign n89016 = P2_P1_UWORD_REG_8_ & ~n88828;
  assign n89017 = P2_P1_EAX_REG_24_ & n88830;
  assign n89018 = ~n89016 & ~n89017;
  assign n15961 = n88949 | ~n89018;
  assign n89020 = P2_P1_UWORD_REG_7_ & ~n88828;
  assign n89021 = P2_P1_EAX_REG_23_ & n88830;
  assign n89022 = ~n89020 & ~n89021;
  assign n15966 = n88954 | ~n89022;
  assign n89024 = P2_P1_UWORD_REG_6_ & ~n88828;
  assign n89025 = P2_P1_EAX_REG_22_ & n88830;
  assign n89026 = ~n89024 & ~n89025;
  assign n15971 = n88959 | ~n89026;
  assign n89028 = P2_P1_UWORD_REG_5_ & ~n88828;
  assign n89029 = P2_P1_EAX_REG_21_ & n88830;
  assign n89030 = ~n89028 & ~n89029;
  assign n15976 = n88964 | ~n89030;
  assign n89032 = P2_P1_EAX_REG_20_ & n88830;
  assign n89033 = P2_P1_UWORD_REG_4_ & ~n88828;
  assign n89034 = ~n88967 & ~n89032;
  assign n15981 = n89033 | ~n89034;
  assign n89036 = P2_P1_EAX_REG_19_ & n88830;
  assign n89037 = P2_P1_UWORD_REG_3_ & ~n88828;
  assign n89038 = ~n88972 & ~n89036;
  assign n15986 = n89037 | ~n89038;
  assign n89040 = P2_P1_EAX_REG_18_ & n88830;
  assign n89041 = P2_P1_UWORD_REG_2_ & ~n88828;
  assign n89042 = ~n88977 & ~n89040;
  assign n15991 = n89041 | ~n89042;
  assign n89044 = P2_P1_EAX_REG_17_ & n88830;
  assign n89045 = P2_P1_UWORD_REG_1_ & ~n88828;
  assign n89046 = ~n88982 & ~n89044;
  assign n15996 = n89045 | ~n89046;
  assign n89048 = P2_P1_EAX_REG_16_ & n88830;
  assign n89049 = P2_P1_UWORD_REG_0_ & ~n88828;
  assign n89050 = ~n88987 & ~n89048;
  assign n16001 = n89049 | ~n89050;
  assign n89052 = ~P2_P1_STATE2_REG_0_ & n76669;
  assign n89053 = n76675 & n77311;
  assign n89054 = ~n77197 & n89053;
  assign n89055 = ~n89052 & ~n89054;
  assign n89056 = P2_P1_STATE2_REG_0_ & ~n89055;
  assign n89057 = P2_P1_EAX_REG_0_ & n89056;
  assign n89058 = ~P2_P1_STATE2_REG_0_ & ~n89055;
  assign n89059 = P2_P1_LWORD_REG_0_ & n89058;
  assign n89060 = P2_P1_DATAO_REG_0_ & n89055;
  assign n89061 = ~n89057 & ~n89059;
  assign n16006 = n89060 | ~n89061;
  assign n89063 = P2_P1_EAX_REG_1_ & n89056;
  assign n89064 = P2_P1_LWORD_REG_1_ & n89058;
  assign n89065 = P2_P1_DATAO_REG_1_ & n89055;
  assign n89066 = ~n89063 & ~n89064;
  assign n16011 = n89065 | ~n89066;
  assign n89068 = P2_P1_EAX_REG_2_ & n89056;
  assign n89069 = P2_P1_LWORD_REG_2_ & n89058;
  assign n89070 = P2_P1_DATAO_REG_2_ & n89055;
  assign n89071 = ~n89068 & ~n89069;
  assign n16016 = n89070 | ~n89071;
  assign n89073 = P2_P1_EAX_REG_3_ & n89056;
  assign n89074 = P2_P1_LWORD_REG_3_ & n89058;
  assign n89075 = P2_P1_DATAO_REG_3_ & n89055;
  assign n89076 = ~n89073 & ~n89074;
  assign n16021 = n89075 | ~n89076;
  assign n89078 = P2_P1_EAX_REG_4_ & n89056;
  assign n89079 = P2_P1_LWORD_REG_4_ & n89058;
  assign n89080 = P2_P1_DATAO_REG_4_ & n89055;
  assign n89081 = ~n89078 & ~n89079;
  assign n16026 = n89080 | ~n89081;
  assign n89083 = P2_P1_EAX_REG_5_ & n89056;
  assign n89084 = P2_P1_LWORD_REG_5_ & n89058;
  assign n89085 = P2_P1_DATAO_REG_5_ & n89055;
  assign n89086 = ~n89083 & ~n89084;
  assign n16031 = n89085 | ~n89086;
  assign n89088 = P2_P1_EAX_REG_6_ & n89056;
  assign n89089 = P2_P1_LWORD_REG_6_ & n89058;
  assign n89090 = P2_P1_DATAO_REG_6_ & n89055;
  assign n89091 = ~n89088 & ~n89089;
  assign n16036 = n89090 | ~n89091;
  assign n89093 = P2_P1_EAX_REG_7_ & n89056;
  assign n89094 = P2_P1_LWORD_REG_7_ & n89058;
  assign n89095 = P2_P1_DATAO_REG_7_ & n89055;
  assign n89096 = ~n89093 & ~n89094;
  assign n16041 = n89095 | ~n89096;
  assign n89098 = P2_P1_EAX_REG_8_ & n89056;
  assign n89099 = P2_P1_LWORD_REG_8_ & n89058;
  assign n89100 = P2_P1_DATAO_REG_8_ & n89055;
  assign n89101 = ~n89098 & ~n89099;
  assign n16046 = n89100 | ~n89101;
  assign n89103 = P2_P1_EAX_REG_9_ & n89056;
  assign n89104 = P2_P1_LWORD_REG_9_ & n89058;
  assign n89105 = P2_P1_DATAO_REG_9_ & n89055;
  assign n89106 = ~n89103 & ~n89104;
  assign n16051 = n89105 | ~n89106;
  assign n89108 = P2_P1_EAX_REG_10_ & n89056;
  assign n89109 = P2_P1_LWORD_REG_10_ & n89058;
  assign n89110 = P2_P1_DATAO_REG_10_ & n89055;
  assign n89111 = ~n89108 & ~n89109;
  assign n16056 = n89110 | ~n89111;
  assign n89113 = P2_P1_EAX_REG_11_ & n89056;
  assign n89114 = P2_P1_LWORD_REG_11_ & n89058;
  assign n89115 = P2_P1_DATAO_REG_11_ & n89055;
  assign n89116 = ~n89113 & ~n89114;
  assign n16061 = n89115 | ~n89116;
  assign n89118 = P2_P1_EAX_REG_12_ & n89056;
  assign n89119 = P2_P1_LWORD_REG_12_ & n89058;
  assign n89120 = P2_P1_DATAO_REG_12_ & n89055;
  assign n89121 = ~n89118 & ~n89119;
  assign n16066 = n89120 | ~n89121;
  assign n89123 = P2_P1_EAX_REG_13_ & n89056;
  assign n89124 = P2_P1_LWORD_REG_13_ & n89058;
  assign n89125 = P2_P1_DATAO_REG_13_ & n89055;
  assign n89126 = ~n89123 & ~n89124;
  assign n16071 = n89125 | ~n89126;
  assign n89128 = P2_P1_EAX_REG_14_ & n89056;
  assign n89129 = P2_P1_LWORD_REG_14_ & n89058;
  assign n89130 = P2_P1_DATAO_REG_14_ & n89055;
  assign n89131 = ~n89128 & ~n89129;
  assign n16076 = n89130 | ~n89131;
  assign n89133 = P2_P1_EAX_REG_15_ & n89056;
  assign n89134 = P2_P1_LWORD_REG_15_ & n89058;
  assign n89135 = P2_P1_DATAO_REG_15_ & n89055;
  assign n89136 = ~n89133 & ~n89134;
  assign n16081 = n89135 | ~n89136;
  assign n89138 = P2_P1_UWORD_REG_0_ & n89058;
  assign n89139 = P2_P1_DATAO_REG_16_ & n89055;
  assign n89140 = ~n89138 & ~n89139;
  assign n89141 = ~n76956 & n89056;
  assign n89142 = P2_P1_EAX_REG_16_ & n89141;
  assign n16086 = ~n89140 | n89142;
  assign n89144 = P2_P1_UWORD_REG_1_ & n89058;
  assign n89145 = P2_P1_DATAO_REG_17_ & n89055;
  assign n89146 = ~n89144 & ~n89145;
  assign n89147 = P2_P1_EAX_REG_17_ & n89141;
  assign n16091 = ~n89146 | n89147;
  assign n89149 = P2_P1_UWORD_REG_2_ & n89058;
  assign n89150 = P2_P1_DATAO_REG_18_ & n89055;
  assign n89151 = ~n89149 & ~n89150;
  assign n89152 = P2_P1_EAX_REG_18_ & n89141;
  assign n16096 = ~n89151 | n89152;
  assign n89154 = P2_P1_UWORD_REG_3_ & n89058;
  assign n89155 = P2_P1_DATAO_REG_19_ & n89055;
  assign n89156 = ~n89154 & ~n89155;
  assign n89157 = P2_P1_EAX_REG_19_ & n89141;
  assign n16101 = ~n89156 | n89157;
  assign n89159 = P2_P1_UWORD_REG_4_ & n89058;
  assign n89160 = P2_P1_DATAO_REG_20_ & n89055;
  assign n89161 = ~n89159 & ~n89160;
  assign n89162 = P2_P1_EAX_REG_20_ & n89141;
  assign n16106 = ~n89161 | n89162;
  assign n89164 = P2_P1_UWORD_REG_5_ & n89058;
  assign n89165 = P2_P1_DATAO_REG_21_ & n89055;
  assign n89166 = ~n89164 & ~n89165;
  assign n89167 = P2_P1_EAX_REG_21_ & n89141;
  assign n16111 = ~n89166 | n89167;
  assign n89169 = P2_P1_UWORD_REG_6_ & n89058;
  assign n89170 = P2_P1_DATAO_REG_22_ & n89055;
  assign n89171 = ~n89169 & ~n89170;
  assign n89172 = P2_P1_EAX_REG_22_ & n89141;
  assign n16116 = ~n89171 | n89172;
  assign n89174 = P2_P1_UWORD_REG_7_ & n89058;
  assign n89175 = P2_P1_DATAO_REG_23_ & n89055;
  assign n89176 = ~n89174 & ~n89175;
  assign n89177 = P2_P1_EAX_REG_23_ & n89141;
  assign n16121 = ~n89176 | n89177;
  assign n89179 = P2_P1_UWORD_REG_8_ & n89058;
  assign n89180 = P2_P1_DATAO_REG_24_ & n89055;
  assign n89181 = ~n89179 & ~n89180;
  assign n89182 = P2_P1_EAX_REG_24_ & n89141;
  assign n16126 = ~n89181 | n89182;
  assign n89184 = P2_P1_UWORD_REG_9_ & n89058;
  assign n89185 = P2_P1_DATAO_REG_25_ & n89055;
  assign n89186 = ~n89184 & ~n89185;
  assign n89187 = P2_P1_EAX_REG_25_ & n89141;
  assign n16131 = ~n89186 | n89187;
  assign n89189 = P2_P1_UWORD_REG_10_ & n89058;
  assign n89190 = P2_P1_DATAO_REG_26_ & n89055;
  assign n89191 = ~n89189 & ~n89190;
  assign n89192 = P2_P1_EAX_REG_26_ & n89141;
  assign n16136 = ~n89191 | n89192;
  assign n89194 = P2_P1_UWORD_REG_11_ & n89058;
  assign n89195 = P2_P1_DATAO_REG_27_ & n89055;
  assign n89196 = ~n89194 & ~n89195;
  assign n89197 = P2_P1_EAX_REG_27_ & n89141;
  assign n16141 = ~n89196 | n89197;
  assign n89199 = P2_P1_UWORD_REG_12_ & n89058;
  assign n89200 = P2_P1_DATAO_REG_28_ & n89055;
  assign n89201 = ~n89199 & ~n89200;
  assign n89202 = P2_P1_EAX_REG_28_ & n89141;
  assign n16146 = ~n89201 | n89202;
  assign n89204 = P2_P1_UWORD_REG_13_ & n89058;
  assign n89205 = P2_P1_DATAO_REG_29_ & n89055;
  assign n89206 = ~n89204 & ~n89205;
  assign n89207 = P2_P1_EAX_REG_29_ & n89141;
  assign n16151 = ~n89206 | n89207;
  assign n89209 = P2_P1_UWORD_REG_14_ & n89058;
  assign n89210 = P2_P1_DATAO_REG_30_ & n89055;
  assign n89211 = ~n89209 & ~n89210;
  assign n89212 = P2_P1_EAX_REG_30_ & n89141;
  assign n16156 = ~n89211 | n89212;
  assign n16161 = P2_P1_DATAO_REG_31_ & n89055;
  assign n89215 = n77191 & ~n77255;
  assign n89216 = n77311 & ~n89215;
  assign n89217 = n77045 & n89216;
  assign n89218 = ~n85327 & n89217;
  assign n89219 = ~n76828 & n89216;
  assign n89220 = ~n77045 & n89219;
  assign n89221 = ~n83790 & n89220;
  assign n89222 = P2_P1_EAX_REG_0_ & ~n89216;
  assign n89223 = n76828 & n89216;
  assign n89224 = ~P2_P1_EAX_REG_0_ & n89223;
  assign n89225 = ~n89222 & ~n89224;
  assign n89226 = ~n89218 & ~n89221;
  assign n16166 = ~n89225 | ~n89226;
  assign n89228 = ~n85445 & n89217;
  assign n89229 = ~n83757 & n89220;
  assign n89230 = P2_P1_EAX_REG_1_ & ~n89216;
  assign n89231 = P2_P1_EAX_REG_0_ & ~P2_P1_EAX_REG_1_;
  assign n89232 = ~P2_P1_EAX_REG_0_ & P2_P1_EAX_REG_1_;
  assign n89233 = ~n89231 & ~n89232;
  assign n89234 = n89223 & ~n89233;
  assign n89235 = ~n89230 & ~n89234;
  assign n89236 = ~n89228 & ~n89229;
  assign n16171 = ~n89235 | ~n89236;
  assign n89238 = ~n85565 & n89217;
  assign n89239 = ~n83712 & n89220;
  assign n89240 = P2_P1_EAX_REG_2_ & ~n89216;
  assign n89241 = P2_P1_EAX_REG_0_ & P2_P1_EAX_REG_1_;
  assign n89242 = ~P2_P1_EAX_REG_2_ & n89241;
  assign n89243 = P2_P1_EAX_REG_2_ & ~n89241;
  assign n89244 = ~n89242 & ~n89243;
  assign n89245 = n89223 & ~n89244;
  assign n89246 = ~n89240 & ~n89245;
  assign n89247 = ~n89238 & ~n89239;
  assign n16176 = ~n89246 | ~n89247;
  assign n89249 = ~n85689 & n89217;
  assign n89250 = ~n83670 & n89220;
  assign n89251 = P2_P1_EAX_REG_3_ & ~n89216;
  assign n89252 = P2_P1_EAX_REG_2_ & n89241;
  assign n89253 = ~P2_P1_EAX_REG_3_ & n89252;
  assign n89254 = P2_P1_EAX_REG_3_ & ~n89252;
  assign n89255 = ~n89253 & ~n89254;
  assign n89256 = n89223 & ~n89255;
  assign n89257 = ~n89251 & ~n89256;
  assign n89258 = ~n89249 & ~n89250;
  assign n16181 = ~n89257 | ~n89258;
  assign n89260 = ~n85816 & n89217;
  assign n89261 = ~n83626 & n89220;
  assign n89262 = P2_P1_EAX_REG_4_ & ~n89216;
  assign n89263 = P2_P1_EAX_REG_3_ & n89252;
  assign n89264 = ~P2_P1_EAX_REG_4_ & n89263;
  assign n89265 = P2_P1_EAX_REG_4_ & ~n89263;
  assign n89266 = ~n89264 & ~n89265;
  assign n89267 = n89223 & ~n89266;
  assign n89268 = ~n89262 & ~n89267;
  assign n89269 = ~n89260 & ~n89261;
  assign n16186 = ~n89268 | ~n89269;
  assign n89271 = ~n85957 & n89217;
  assign n89272 = ~n83582 & n89220;
  assign n89273 = P2_P1_EAX_REG_5_ & ~n89216;
  assign n89274 = P2_P1_EAX_REG_4_ & n89263;
  assign n89275 = ~P2_P1_EAX_REG_5_ & n89274;
  assign n89276 = P2_P1_EAX_REG_5_ & ~n89274;
  assign n89277 = ~n89275 & ~n89276;
  assign n89278 = n89223 & ~n89277;
  assign n89279 = ~n89273 & ~n89278;
  assign n89280 = ~n89271 & ~n89272;
  assign n16191 = ~n89279 | ~n89280;
  assign n89282 = ~n83535 & n89220;
  assign n89283 = P2_P1_EAX_REG_6_ & ~n89216;
  assign n89284 = P2_P1_EAX_REG_5_ & n89274;
  assign n89285 = ~P2_P1_EAX_REG_6_ & n89284;
  assign n89286 = P2_P1_EAX_REG_6_ & ~n89284;
  assign n89287 = ~n89285 & ~n89286;
  assign n89288 = n89223 & ~n89287;
  assign n89289 = ~n86089 & n89217;
  assign n89290 = ~n89283 & ~n89288;
  assign n89291 = ~n89289 & n89290;
  assign n16196 = n89282 | ~n89291;
  assign n89293 = ~n77700 & n89220;
  assign n89294 = P2_P1_EAX_REG_7_ & ~n89216;
  assign n89295 = P2_P1_EAX_REG_6_ & n89284;
  assign n89296 = ~P2_P1_EAX_REG_7_ & n89295;
  assign n89297 = P2_P1_EAX_REG_7_ & ~n89295;
  assign n89298 = ~n89296 & ~n89297;
  assign n89299 = n89223 & ~n89298;
  assign n89300 = ~n85361 & n89217;
  assign n89301 = ~n89294 & ~n89299;
  assign n89302 = ~n89300 & n89301;
  assign n16201 = n89293 | ~n89302;
  assign n89304 = ~n88948 & n89220;
  assign n89305 = P2_P1_EAX_REG_8_ & ~n89216;
  assign n89306 = P2_P1_EAX_REG_7_ & n89295;
  assign n89307 = ~P2_P1_EAX_REG_8_ & n89306;
  assign n89308 = P2_P1_EAX_REG_8_ & ~n89306;
  assign n89309 = ~n89307 & ~n89308;
  assign n89310 = n89223 & ~n89309;
  assign n89311 = ~n77205 & ~n77212;
  assign n89312 = ~n77156 & ~n89311;
  assign n89313 = n76686 & n89312;
  assign n89314 = P2_P1_INSTQUEUE_REG_15__0_ & n89313;
  assign n89315 = n76690 & n89312;
  assign n89316 = P2_P1_INSTQUEUE_REG_14__0_ & n89315;
  assign n89317 = n76677 & n89312;
  assign n89318 = P2_P1_INSTQUEUE_REG_13__0_ & n89317;
  assign n89319 = n76681 & n89312;
  assign n89320 = P2_P1_INSTQUEUE_REG_12__0_ & n89319;
  assign n89321 = ~n89314 & ~n89316;
  assign n89322 = ~n89318 & n89321;
  assign n89323 = ~n89320 & n89322;
  assign n89324 = n77156 & ~n89311;
  assign n89325 = n76686 & n89324;
  assign n89326 = P2_P1_INSTQUEUE_REG_11__0_ & n89325;
  assign n89327 = n76690 & n89324;
  assign n89328 = P2_P1_INSTQUEUE_REG_10__0_ & n89327;
  assign n89329 = n76677 & n89324;
  assign n89330 = P2_P1_INSTQUEUE_REG_9__0_ & n89329;
  assign n89331 = n76681 & n89324;
  assign n89332 = P2_P1_INSTQUEUE_REG_8__0_ & n89331;
  assign n89333 = ~n89326 & ~n89328;
  assign n89334 = ~n89330 & n89333;
  assign n89335 = ~n89332 & n89334;
  assign n89336 = ~n77156 & n89311;
  assign n89337 = n76686 & n89336;
  assign n89338 = P2_P1_INSTQUEUE_REG_7__0_ & n89337;
  assign n89339 = n76690 & n89336;
  assign n89340 = P2_P1_INSTQUEUE_REG_6__0_ & n89339;
  assign n89341 = n76677 & n89336;
  assign n89342 = P2_P1_INSTQUEUE_REG_5__0_ & n89341;
  assign n89343 = n76681 & n89336;
  assign n89344 = P2_P1_INSTQUEUE_REG_4__0_ & n89343;
  assign n89345 = ~n89338 & ~n89340;
  assign n89346 = ~n89342 & n89345;
  assign n89347 = ~n89344 & n89346;
  assign n89348 = n77156 & n89311;
  assign n89349 = n76686 & n89348;
  assign n89350 = P2_P1_INSTQUEUE_REG_3__0_ & n89349;
  assign n89351 = n76690 & n89348;
  assign n89352 = P2_P1_INSTQUEUE_REG_2__0_ & n89351;
  assign n89353 = n76677 & n89348;
  assign n89354 = P2_P1_INSTQUEUE_REG_1__0_ & n89353;
  assign n89355 = n76681 & n89348;
  assign n89356 = P2_P1_INSTQUEUE_REG_0__0_ & n89355;
  assign n89357 = ~n89350 & ~n89352;
  assign n89358 = ~n89354 & n89357;
  assign n89359 = ~n89356 & n89358;
  assign n89360 = n89323 & n89335;
  assign n89361 = n89347 & n89360;
  assign n89362 = n89359 & n89361;
  assign n89363 = n89217 & ~n89362;
  assign n89364 = ~n89305 & ~n89310;
  assign n89365 = ~n89363 & n89364;
  assign n16206 = n89304 | ~n89365;
  assign n89367 = ~n88931 & n89220;
  assign n89368 = P2_P1_EAX_REG_9_ & ~n89216;
  assign n89369 = P2_P1_EAX_REG_8_ & n89306;
  assign n89370 = ~P2_P1_EAX_REG_9_ & n89369;
  assign n89371 = P2_P1_EAX_REG_9_ & ~n89369;
  assign n89372 = ~n89370 & ~n89371;
  assign n89373 = n89223 & ~n89372;
  assign n89374 = P2_P1_INSTQUEUE_REG_15__1_ & n89313;
  assign n89375 = P2_P1_INSTQUEUE_REG_14__1_ & n89315;
  assign n89376 = P2_P1_INSTQUEUE_REG_13__1_ & n89317;
  assign n89377 = P2_P1_INSTQUEUE_REG_12__1_ & n89319;
  assign n89378 = ~n89374 & ~n89375;
  assign n89379 = ~n89376 & n89378;
  assign n89380 = ~n89377 & n89379;
  assign n89381 = P2_P1_INSTQUEUE_REG_11__1_ & n89325;
  assign n89382 = P2_P1_INSTQUEUE_REG_10__1_ & n89327;
  assign n89383 = P2_P1_INSTQUEUE_REG_9__1_ & n89329;
  assign n89384 = P2_P1_INSTQUEUE_REG_8__1_ & n89331;
  assign n89385 = ~n89381 & ~n89382;
  assign n89386 = ~n89383 & n89385;
  assign n89387 = ~n89384 & n89386;
  assign n89388 = P2_P1_INSTQUEUE_REG_7__1_ & n89337;
  assign n89389 = P2_P1_INSTQUEUE_REG_6__1_ & n89339;
  assign n89390 = P2_P1_INSTQUEUE_REG_5__1_ & n89341;
  assign n89391 = P2_P1_INSTQUEUE_REG_4__1_ & n89343;
  assign n89392 = ~n89388 & ~n89389;
  assign n89393 = ~n89390 & n89392;
  assign n89394 = ~n89391 & n89393;
  assign n89395 = P2_P1_INSTQUEUE_REG_3__1_ & n89349;
  assign n89396 = P2_P1_INSTQUEUE_REG_2__1_ & n89351;
  assign n89397 = P2_P1_INSTQUEUE_REG_1__1_ & n89353;
  assign n89398 = P2_P1_INSTQUEUE_REG_0__1_ & n89355;
  assign n89399 = ~n89395 & ~n89396;
  assign n89400 = ~n89397 & n89399;
  assign n89401 = ~n89398 & n89400;
  assign n89402 = n89380 & n89387;
  assign n89403 = n89394 & n89402;
  assign n89404 = n89401 & n89403;
  assign n89405 = n89217 & ~n89404;
  assign n89406 = ~n89368 & ~n89373;
  assign n89407 = ~n89405 & n89406;
  assign n16211 = n89367 | ~n89407;
  assign n89409 = ~n88919 & n89220;
  assign n89410 = P2_P1_EAX_REG_10_ & ~n89216;
  assign n89411 = P2_P1_EAX_REG_9_ & n89369;
  assign n89412 = ~P2_P1_EAX_REG_10_ & n89411;
  assign n89413 = P2_P1_EAX_REG_10_ & ~n89411;
  assign n89414 = ~n89412 & ~n89413;
  assign n89415 = n89223 & ~n89414;
  assign n89416 = P2_P1_INSTQUEUE_REG_15__2_ & n89313;
  assign n89417 = P2_P1_INSTQUEUE_REG_14__2_ & n89315;
  assign n89418 = P2_P1_INSTQUEUE_REG_13__2_ & n89317;
  assign n89419 = P2_P1_INSTQUEUE_REG_12__2_ & n89319;
  assign n89420 = ~n89416 & ~n89417;
  assign n89421 = ~n89418 & n89420;
  assign n89422 = ~n89419 & n89421;
  assign n89423 = P2_P1_INSTQUEUE_REG_11__2_ & n89325;
  assign n89424 = P2_P1_INSTQUEUE_REG_10__2_ & n89327;
  assign n89425 = P2_P1_INSTQUEUE_REG_9__2_ & n89329;
  assign n89426 = P2_P1_INSTQUEUE_REG_8__2_ & n89331;
  assign n89427 = ~n89423 & ~n89424;
  assign n89428 = ~n89425 & n89427;
  assign n89429 = ~n89426 & n89428;
  assign n89430 = P2_P1_INSTQUEUE_REG_7__2_ & n89337;
  assign n89431 = P2_P1_INSTQUEUE_REG_6__2_ & n89339;
  assign n89432 = P2_P1_INSTQUEUE_REG_5__2_ & n89341;
  assign n89433 = P2_P1_INSTQUEUE_REG_4__2_ & n89343;
  assign n89434 = ~n89430 & ~n89431;
  assign n89435 = ~n89432 & n89434;
  assign n89436 = ~n89433 & n89435;
  assign n89437 = P2_P1_INSTQUEUE_REG_3__2_ & n89349;
  assign n89438 = P2_P1_INSTQUEUE_REG_2__2_ & n89351;
  assign n89439 = P2_P1_INSTQUEUE_REG_1__2_ & n89353;
  assign n89440 = P2_P1_INSTQUEUE_REG_0__2_ & n89355;
  assign n89441 = ~n89437 & ~n89438;
  assign n89442 = ~n89439 & n89441;
  assign n89443 = ~n89440 & n89442;
  assign n89444 = n89422 & n89429;
  assign n89445 = n89436 & n89444;
  assign n89446 = n89443 & n89445;
  assign n89447 = n89217 & ~n89446;
  assign n89448 = ~n89410 & ~n89415;
  assign n89449 = ~n89447 & n89448;
  assign n16216 = n89409 | ~n89449;
  assign n89451 = ~n88903 & n89220;
  assign n89452 = P2_P1_EAX_REG_11_ & ~n89216;
  assign n89453 = P2_P1_EAX_REG_10_ & n89411;
  assign n89454 = ~P2_P1_EAX_REG_11_ & n89453;
  assign n89455 = P2_P1_EAX_REG_11_ & ~n89453;
  assign n89456 = ~n89454 & ~n89455;
  assign n89457 = n89223 & ~n89456;
  assign n89458 = P2_P1_INSTQUEUE_REG_15__3_ & n89313;
  assign n89459 = P2_P1_INSTQUEUE_REG_14__3_ & n89315;
  assign n89460 = P2_P1_INSTQUEUE_REG_13__3_ & n89317;
  assign n89461 = P2_P1_INSTQUEUE_REG_12__3_ & n89319;
  assign n89462 = ~n89458 & ~n89459;
  assign n89463 = ~n89460 & n89462;
  assign n89464 = ~n89461 & n89463;
  assign n89465 = P2_P1_INSTQUEUE_REG_11__3_ & n89325;
  assign n89466 = P2_P1_INSTQUEUE_REG_10__3_ & n89327;
  assign n89467 = P2_P1_INSTQUEUE_REG_9__3_ & n89329;
  assign n89468 = P2_P1_INSTQUEUE_REG_8__3_ & n89331;
  assign n89469 = ~n89465 & ~n89466;
  assign n89470 = ~n89467 & n89469;
  assign n89471 = ~n89468 & n89470;
  assign n89472 = P2_P1_INSTQUEUE_REG_7__3_ & n89337;
  assign n89473 = P2_P1_INSTQUEUE_REG_6__3_ & n89339;
  assign n89474 = P2_P1_INSTQUEUE_REG_5__3_ & n89341;
  assign n89475 = P2_P1_INSTQUEUE_REG_4__3_ & n89343;
  assign n89476 = ~n89472 & ~n89473;
  assign n89477 = ~n89474 & n89476;
  assign n89478 = ~n89475 & n89477;
  assign n89479 = P2_P1_INSTQUEUE_REG_3__3_ & n89349;
  assign n89480 = P2_P1_INSTQUEUE_REG_2__3_ & n89351;
  assign n89481 = P2_P1_INSTQUEUE_REG_1__3_ & n89353;
  assign n89482 = P2_P1_INSTQUEUE_REG_0__3_ & n89355;
  assign n89483 = ~n89479 & ~n89480;
  assign n89484 = ~n89481 & n89483;
  assign n89485 = ~n89482 & n89484;
  assign n89486 = n89464 & n89471;
  assign n89487 = n89478 & n89486;
  assign n89488 = n89485 & n89487;
  assign n89489 = n89217 & ~n89488;
  assign n89490 = ~n89452 & ~n89457;
  assign n89491 = ~n89489 & n89490;
  assign n16221 = n89451 | ~n89491;
  assign n89493 = ~n88888 & n89220;
  assign n89494 = P2_P1_EAX_REG_12_ & ~n89216;
  assign n89495 = P2_P1_INSTQUEUE_REG_15__4_ & n89313;
  assign n89496 = P2_P1_INSTQUEUE_REG_14__4_ & n89315;
  assign n89497 = P2_P1_INSTQUEUE_REG_13__4_ & n89317;
  assign n89498 = P2_P1_INSTQUEUE_REG_12__4_ & n89319;
  assign n89499 = ~n89495 & ~n89496;
  assign n89500 = ~n89497 & n89499;
  assign n89501 = ~n89498 & n89500;
  assign n89502 = P2_P1_INSTQUEUE_REG_11__4_ & n89325;
  assign n89503 = P2_P1_INSTQUEUE_REG_10__4_ & n89327;
  assign n89504 = P2_P1_INSTQUEUE_REG_9__4_ & n89329;
  assign n89505 = P2_P1_INSTQUEUE_REG_8__4_ & n89331;
  assign n89506 = ~n89502 & ~n89503;
  assign n89507 = ~n89504 & n89506;
  assign n89508 = ~n89505 & n89507;
  assign n89509 = P2_P1_INSTQUEUE_REG_7__4_ & n89337;
  assign n89510 = P2_P1_INSTQUEUE_REG_6__4_ & n89339;
  assign n89511 = P2_P1_INSTQUEUE_REG_5__4_ & n89341;
  assign n89512 = P2_P1_INSTQUEUE_REG_4__4_ & n89343;
  assign n89513 = ~n89509 & ~n89510;
  assign n89514 = ~n89511 & n89513;
  assign n89515 = ~n89512 & n89514;
  assign n89516 = P2_P1_INSTQUEUE_REG_3__4_ & n89349;
  assign n89517 = P2_P1_INSTQUEUE_REG_2__4_ & n89351;
  assign n89518 = P2_P1_INSTQUEUE_REG_1__4_ & n89353;
  assign n89519 = P2_P1_INSTQUEUE_REG_0__4_ & n89355;
  assign n89520 = ~n89516 & ~n89517;
  assign n89521 = ~n89518 & n89520;
  assign n89522 = ~n89519 & n89521;
  assign n89523 = n89501 & n89508;
  assign n89524 = n89515 & n89523;
  assign n89525 = n89522 & n89524;
  assign n89526 = n89217 & ~n89525;
  assign n89527 = P2_P1_EAX_REG_11_ & n89453;
  assign n89528 = ~P2_P1_EAX_REG_12_ & n89527;
  assign n89529 = P2_P1_EAX_REG_12_ & ~n89527;
  assign n89530 = ~n89528 & ~n89529;
  assign n89531 = n89223 & ~n89530;
  assign n89532 = ~n89494 & ~n89526;
  assign n89533 = ~n89531 & n89532;
  assign n16226 = n89493 | ~n89533;
  assign n89535 = ~n88872 & n89220;
  assign n89536 = P2_P1_EAX_REG_13_ & ~n89216;
  assign n89537 = P2_P1_INSTQUEUE_REG_15__5_ & n89313;
  assign n89538 = P2_P1_INSTQUEUE_REG_14__5_ & n89315;
  assign n89539 = P2_P1_INSTQUEUE_REG_13__5_ & n89317;
  assign n89540 = P2_P1_INSTQUEUE_REG_12__5_ & n89319;
  assign n89541 = ~n89537 & ~n89538;
  assign n89542 = ~n89539 & n89541;
  assign n89543 = ~n89540 & n89542;
  assign n89544 = P2_P1_INSTQUEUE_REG_11__5_ & n89325;
  assign n89545 = P2_P1_INSTQUEUE_REG_10__5_ & n89327;
  assign n89546 = P2_P1_INSTQUEUE_REG_9__5_ & n89329;
  assign n89547 = P2_P1_INSTQUEUE_REG_8__5_ & n89331;
  assign n89548 = ~n89544 & ~n89545;
  assign n89549 = ~n89546 & n89548;
  assign n89550 = ~n89547 & n89549;
  assign n89551 = P2_P1_INSTQUEUE_REG_7__5_ & n89337;
  assign n89552 = P2_P1_INSTQUEUE_REG_6__5_ & n89339;
  assign n89553 = P2_P1_INSTQUEUE_REG_5__5_ & n89341;
  assign n89554 = P2_P1_INSTQUEUE_REG_4__5_ & n89343;
  assign n89555 = ~n89551 & ~n89552;
  assign n89556 = ~n89553 & n89555;
  assign n89557 = ~n89554 & n89556;
  assign n89558 = P2_P1_INSTQUEUE_REG_3__5_ & n89349;
  assign n89559 = P2_P1_INSTQUEUE_REG_2__5_ & n89351;
  assign n89560 = P2_P1_INSTQUEUE_REG_1__5_ & n89353;
  assign n89561 = P2_P1_INSTQUEUE_REG_0__5_ & n89355;
  assign n89562 = ~n89558 & ~n89559;
  assign n89563 = ~n89560 & n89562;
  assign n89564 = ~n89561 & n89563;
  assign n89565 = n89543 & n89550;
  assign n89566 = n89557 & n89565;
  assign n89567 = n89564 & n89566;
  assign n89568 = n89217 & ~n89567;
  assign n89569 = P2_P1_EAX_REG_12_ & n89527;
  assign n89570 = ~P2_P1_EAX_REG_13_ & n89569;
  assign n89571 = P2_P1_EAX_REG_13_ & ~n89569;
  assign n89572 = ~n89570 & ~n89571;
  assign n89573 = n89223 & ~n89572;
  assign n89574 = ~n89536 & ~n89568;
  assign n89575 = ~n89573 & n89574;
  assign n16231 = n89535 | ~n89575;
  assign n89577 = ~n88858 & n89220;
  assign n89578 = P2_P1_EAX_REG_14_ & ~n89216;
  assign n89579 = P2_P1_INSTQUEUE_REG_15__6_ & n89313;
  assign n89580 = P2_P1_INSTQUEUE_REG_14__6_ & n89315;
  assign n89581 = P2_P1_INSTQUEUE_REG_13__6_ & n89317;
  assign n89582 = P2_P1_INSTQUEUE_REG_12__6_ & n89319;
  assign n89583 = ~n89579 & ~n89580;
  assign n89584 = ~n89581 & n89583;
  assign n89585 = ~n89582 & n89584;
  assign n89586 = P2_P1_INSTQUEUE_REG_11__6_ & n89325;
  assign n89587 = P2_P1_INSTQUEUE_REG_10__6_ & n89327;
  assign n89588 = P2_P1_INSTQUEUE_REG_9__6_ & n89329;
  assign n89589 = P2_P1_INSTQUEUE_REG_8__6_ & n89331;
  assign n89590 = ~n89586 & ~n89587;
  assign n89591 = ~n89588 & n89590;
  assign n89592 = ~n89589 & n89591;
  assign n89593 = P2_P1_INSTQUEUE_REG_7__6_ & n89337;
  assign n89594 = P2_P1_INSTQUEUE_REG_6__6_ & n89339;
  assign n89595 = P2_P1_INSTQUEUE_REG_5__6_ & n89341;
  assign n89596 = P2_P1_INSTQUEUE_REG_4__6_ & n89343;
  assign n89597 = ~n89593 & ~n89594;
  assign n89598 = ~n89595 & n89597;
  assign n89599 = ~n89596 & n89598;
  assign n89600 = P2_P1_INSTQUEUE_REG_3__6_ & n89349;
  assign n89601 = P2_P1_INSTQUEUE_REG_2__6_ & n89351;
  assign n89602 = P2_P1_INSTQUEUE_REG_1__6_ & n89353;
  assign n89603 = P2_P1_INSTQUEUE_REG_0__6_ & n89355;
  assign n89604 = ~n89600 & ~n89601;
  assign n89605 = ~n89602 & n89604;
  assign n89606 = ~n89603 & n89605;
  assign n89607 = n89585 & n89592;
  assign n89608 = n89599 & n89607;
  assign n89609 = n89606 & n89608;
  assign n89610 = n89217 & ~n89609;
  assign n89611 = P2_P1_EAX_REG_13_ & n89569;
  assign n89612 = ~P2_P1_EAX_REG_14_ & n89611;
  assign n89613 = P2_P1_EAX_REG_14_ & ~n89611;
  assign n89614 = ~n89612 & ~n89613;
  assign n89615 = n89223 & ~n89614;
  assign n89616 = ~n89578 & ~n89610;
  assign n89617 = ~n89615 & n89616;
  assign n16236 = n89577 | ~n89617;
  assign n89619 = ~n88841 & n89220;
  assign n89620 = P2_P1_EAX_REG_15_ & ~n89216;
  assign n89621 = P2_P1_INSTQUEUE_REG_15__7_ & n89313;
  assign n89622 = P2_P1_INSTQUEUE_REG_14__7_ & n89315;
  assign n89623 = P2_P1_INSTQUEUE_REG_13__7_ & n89317;
  assign n89624 = P2_P1_INSTQUEUE_REG_12__7_ & n89319;
  assign n89625 = ~n89621 & ~n89622;
  assign n89626 = ~n89623 & n89625;
  assign n89627 = ~n89624 & n89626;
  assign n89628 = P2_P1_INSTQUEUE_REG_11__7_ & n89325;
  assign n89629 = P2_P1_INSTQUEUE_REG_10__7_ & n89327;
  assign n89630 = P2_P1_INSTQUEUE_REG_9__7_ & n89329;
  assign n89631 = P2_P1_INSTQUEUE_REG_8__7_ & n89331;
  assign n89632 = ~n89628 & ~n89629;
  assign n89633 = ~n89630 & n89632;
  assign n89634 = ~n89631 & n89633;
  assign n89635 = P2_P1_INSTQUEUE_REG_7__7_ & n89337;
  assign n89636 = P2_P1_INSTQUEUE_REG_6__7_ & n89339;
  assign n89637 = P2_P1_INSTQUEUE_REG_5__7_ & n89341;
  assign n89638 = P2_P1_INSTQUEUE_REG_4__7_ & n89343;
  assign n89639 = ~n89635 & ~n89636;
  assign n89640 = ~n89637 & n89639;
  assign n89641 = ~n89638 & n89640;
  assign n89642 = P2_P1_INSTQUEUE_REG_3__7_ & n89349;
  assign n89643 = P2_P1_INSTQUEUE_REG_2__7_ & n89351;
  assign n89644 = P2_P1_INSTQUEUE_REG_1__7_ & n89353;
  assign n89645 = P2_P1_INSTQUEUE_REG_0__7_ & n89355;
  assign n89646 = ~n89642 & ~n89643;
  assign n89647 = ~n89644 & n89646;
  assign n89648 = ~n89645 & n89647;
  assign n89649 = n89627 & n89634;
  assign n89650 = n89641 & n89649;
  assign n89651 = n89648 & n89650;
  assign n89652 = n89217 & ~n89651;
  assign n89653 = P2_P1_EAX_REG_14_ & n89611;
  assign n89654 = ~P2_P1_EAX_REG_15_ & n89653;
  assign n89655 = P2_P1_EAX_REG_15_ & ~n89653;
  assign n89656 = ~n89654 & ~n89655;
  assign n89657 = n89223 & ~n89656;
  assign n89658 = ~n89620 & ~n89652;
  assign n89659 = ~n89657 & n89658;
  assign n16241 = n89619 | ~n89659;
  assign n89661 = P2_P1_INSTQUEUERD_ADDR_REG_2_ & ~n76690;
  assign n89662 = ~P2_P1_INSTQUEUERD_ADDR_REG_3_ & n89661;
  assign n89663 = P2_P1_INSTQUEUERD_ADDR_REG_3_ & ~n89661;
  assign n89664 = ~n89662 & ~n89663;
  assign n89665 = ~n76691 & ~n89661;
  assign n89666 = n89664 & n89665;
  assign n89667 = n85277 & n89666;
  assign n89668 = P2_P1_INSTQUEUE_REG_7__0_ & n89667;
  assign n89669 = n85274 & n89666;
  assign n89670 = P2_P1_INSTQUEUE_REG_6__0_ & n89669;
  assign n89671 = n85283 & n89666;
  assign n89672 = P2_P1_INSTQUEUE_REG_5__0_ & n89671;
  assign n89673 = n85280 & n89666;
  assign n89674 = P2_P1_INSTQUEUE_REG_4__0_ & n89673;
  assign n89675 = ~n89668 & ~n89670;
  assign n89676 = ~n89672 & n89675;
  assign n89677 = ~n89674 & n89676;
  assign n89678 = n89664 & ~n89665;
  assign n89679 = n85277 & n89678;
  assign n89680 = P2_P1_INSTQUEUE_REG_3__0_ & n89679;
  assign n89681 = n85274 & n89678;
  assign n89682 = P2_P1_INSTQUEUE_REG_2__0_ & n89681;
  assign n89683 = n85283 & n89678;
  assign n89684 = P2_P1_INSTQUEUE_REG_1__0_ & n89683;
  assign n89685 = n85280 & n89678;
  assign n89686 = P2_P1_INSTQUEUE_REG_0__0_ & n89685;
  assign n89687 = ~n89680 & ~n89682;
  assign n89688 = ~n89684 & n89687;
  assign n89689 = ~n89686 & n89688;
  assign n89690 = ~n89664 & n89665;
  assign n89691 = n85277 & n89690;
  assign n89692 = P2_P1_INSTQUEUE_REG_15__0_ & n89691;
  assign n89693 = n85274 & n89690;
  assign n89694 = P2_P1_INSTQUEUE_REG_14__0_ & n89693;
  assign n89695 = n85283 & n89690;
  assign n89696 = P2_P1_INSTQUEUE_REG_13__0_ & n89695;
  assign n89697 = n85280 & n89690;
  assign n89698 = P2_P1_INSTQUEUE_REG_12__0_ & n89697;
  assign n89699 = ~n89692 & ~n89694;
  assign n89700 = ~n89696 & n89699;
  assign n89701 = ~n89698 & n89700;
  assign n89702 = ~n89664 & ~n89665;
  assign n89703 = n85277 & n89702;
  assign n89704 = P2_P1_INSTQUEUE_REG_11__0_ & n89703;
  assign n89705 = n85274 & n89702;
  assign n89706 = P2_P1_INSTQUEUE_REG_10__0_ & n89705;
  assign n89707 = n85283 & n89702;
  assign n89708 = P2_P1_INSTQUEUE_REG_9__0_ & n89707;
  assign n89709 = n85280 & n89702;
  assign n89710 = P2_P1_INSTQUEUE_REG_8__0_ & n89709;
  assign n89711 = ~n89704 & ~n89706;
  assign n89712 = ~n89708 & n89711;
  assign n89713 = ~n89710 & n89712;
  assign n89714 = n89677 & n89689;
  assign n89715 = n89701 & n89714;
  assign n89716 = n89713 & n89715;
  assign n89717 = n89217 & ~n89716;
  assign n89718 = n76734 & n89219;
  assign n89719 = ~n83790 & n89718;
  assign n89720 = P2_P1_EAX_REG_16_ & ~n89216;
  assign n89721 = P2_P1_EAX_REG_15_ & n89653;
  assign n89722 = ~P2_P1_EAX_REG_16_ & n89721;
  assign n89723 = P2_P1_EAX_REG_16_ & ~n89721;
  assign n89724 = ~n89722 & ~n89723;
  assign n89725 = n89223 & ~n89724;
  assign n89726 = ~n76765 & n89219;
  assign n89727 = ~n83805 & n89726;
  assign n89728 = ~n89717 & ~n89719;
  assign n89729 = ~n89720 & n89728;
  assign n89730 = ~n89725 & n89729;
  assign n16246 = n89727 | ~n89730;
  assign n89732 = P2_P1_INSTQUEUE_REG_7__1_ & n89667;
  assign n89733 = P2_P1_INSTQUEUE_REG_6__1_ & n89669;
  assign n89734 = P2_P1_INSTQUEUE_REG_5__1_ & n89671;
  assign n89735 = P2_P1_INSTQUEUE_REG_4__1_ & n89673;
  assign n89736 = ~n89732 & ~n89733;
  assign n89737 = ~n89734 & n89736;
  assign n89738 = ~n89735 & n89737;
  assign n89739 = P2_P1_INSTQUEUE_REG_3__1_ & n89679;
  assign n89740 = P2_P1_INSTQUEUE_REG_2__1_ & n89681;
  assign n89741 = P2_P1_INSTQUEUE_REG_1__1_ & n89683;
  assign n89742 = P2_P1_INSTQUEUE_REG_0__1_ & n89685;
  assign n89743 = ~n89739 & ~n89740;
  assign n89744 = ~n89741 & n89743;
  assign n89745 = ~n89742 & n89744;
  assign n89746 = P2_P1_INSTQUEUE_REG_15__1_ & n89691;
  assign n89747 = P2_P1_INSTQUEUE_REG_14__1_ & n89693;
  assign n89748 = P2_P1_INSTQUEUE_REG_13__1_ & n89695;
  assign n89749 = P2_P1_INSTQUEUE_REG_12__1_ & n89697;
  assign n89750 = ~n89746 & ~n89747;
  assign n89751 = ~n89748 & n89750;
  assign n89752 = ~n89749 & n89751;
  assign n89753 = P2_P1_INSTQUEUE_REG_11__1_ & n89703;
  assign n89754 = P2_P1_INSTQUEUE_REG_10__1_ & n89705;
  assign n89755 = P2_P1_INSTQUEUE_REG_9__1_ & n89707;
  assign n89756 = P2_P1_INSTQUEUE_REG_8__1_ & n89709;
  assign n89757 = ~n89753 & ~n89754;
  assign n89758 = ~n89755 & n89757;
  assign n89759 = ~n89756 & n89758;
  assign n89760 = n89738 & n89745;
  assign n89761 = n89752 & n89760;
  assign n89762 = n89759 & n89761;
  assign n89763 = n89217 & ~n89762;
  assign n89764 = ~n83757 & n89718;
  assign n89765 = P2_P1_EAX_REG_17_ & ~n89216;
  assign n89766 = P2_P1_EAX_REG_16_ & n89721;
  assign n89767 = ~P2_P1_EAX_REG_17_ & n89766;
  assign n89768 = P2_P1_EAX_REG_17_ & ~n89766;
  assign n89769 = ~n89767 & ~n89768;
  assign n89770 = n89223 & ~n89769;
  assign n89771 = ~n83768 & n89726;
  assign n89772 = ~n89763 & ~n89764;
  assign n89773 = ~n89765 & n89772;
  assign n89774 = ~n89770 & n89773;
  assign n16251 = n89771 | ~n89774;
  assign n89776 = P2_P1_INSTQUEUE_REG_7__2_ & n89667;
  assign n89777 = P2_P1_INSTQUEUE_REG_6__2_ & n89669;
  assign n89778 = P2_P1_INSTQUEUE_REG_5__2_ & n89671;
  assign n89779 = P2_P1_INSTQUEUE_REG_4__2_ & n89673;
  assign n89780 = ~n89776 & ~n89777;
  assign n89781 = ~n89778 & n89780;
  assign n89782 = ~n89779 & n89781;
  assign n89783 = P2_P1_INSTQUEUE_REG_3__2_ & n89679;
  assign n89784 = P2_P1_INSTQUEUE_REG_2__2_ & n89681;
  assign n89785 = P2_P1_INSTQUEUE_REG_1__2_ & n89683;
  assign n89786 = P2_P1_INSTQUEUE_REG_0__2_ & n89685;
  assign n89787 = ~n89783 & ~n89784;
  assign n89788 = ~n89785 & n89787;
  assign n89789 = ~n89786 & n89788;
  assign n89790 = P2_P1_INSTQUEUE_REG_15__2_ & n89691;
  assign n89791 = P2_P1_INSTQUEUE_REG_14__2_ & n89693;
  assign n89792 = P2_P1_INSTQUEUE_REG_13__2_ & n89695;
  assign n89793 = P2_P1_INSTQUEUE_REG_12__2_ & n89697;
  assign n89794 = ~n89790 & ~n89791;
  assign n89795 = ~n89792 & n89794;
  assign n89796 = ~n89793 & n89795;
  assign n89797 = P2_P1_INSTQUEUE_REG_11__2_ & n89703;
  assign n89798 = P2_P1_INSTQUEUE_REG_10__2_ & n89705;
  assign n89799 = P2_P1_INSTQUEUE_REG_9__2_ & n89707;
  assign n89800 = P2_P1_INSTQUEUE_REG_8__2_ & n89709;
  assign n89801 = ~n89797 & ~n89798;
  assign n89802 = ~n89799 & n89801;
  assign n89803 = ~n89800 & n89802;
  assign n89804 = n89782 & n89789;
  assign n89805 = n89796 & n89804;
  assign n89806 = n89803 & n89805;
  assign n89807 = n89217 & ~n89806;
  assign n89808 = ~n83712 & n89718;
  assign n89809 = P2_P1_EAX_REG_18_ & ~n89216;
  assign n89810 = P2_P1_EAX_REG_17_ & n89766;
  assign n89811 = ~P2_P1_EAX_REG_18_ & n89810;
  assign n89812 = P2_P1_EAX_REG_18_ & ~n89810;
  assign n89813 = ~n89811 & ~n89812;
  assign n89814 = n89223 & ~n89813;
  assign n89815 = ~n83728 & n89726;
  assign n89816 = ~n89807 & ~n89808;
  assign n89817 = ~n89809 & n89816;
  assign n89818 = ~n89814 & n89817;
  assign n16256 = n89815 | ~n89818;
  assign n89820 = P2_P1_INSTQUEUE_REG_7__3_ & n89667;
  assign n89821 = P2_P1_INSTQUEUE_REG_6__3_ & n89669;
  assign n89822 = P2_P1_INSTQUEUE_REG_5__3_ & n89671;
  assign n89823 = P2_P1_INSTQUEUE_REG_4__3_ & n89673;
  assign n89824 = ~n89820 & ~n89821;
  assign n89825 = ~n89822 & n89824;
  assign n89826 = ~n89823 & n89825;
  assign n89827 = P2_P1_INSTQUEUE_REG_3__3_ & n89679;
  assign n89828 = P2_P1_INSTQUEUE_REG_2__3_ & n89681;
  assign n89829 = P2_P1_INSTQUEUE_REG_1__3_ & n89683;
  assign n89830 = P2_P1_INSTQUEUE_REG_0__3_ & n89685;
  assign n89831 = ~n89827 & ~n89828;
  assign n89832 = ~n89829 & n89831;
  assign n89833 = ~n89830 & n89832;
  assign n89834 = P2_P1_INSTQUEUE_REG_15__3_ & n89691;
  assign n89835 = P2_P1_INSTQUEUE_REG_14__3_ & n89693;
  assign n89836 = P2_P1_INSTQUEUE_REG_13__3_ & n89695;
  assign n89837 = P2_P1_INSTQUEUE_REG_12__3_ & n89697;
  assign n89838 = ~n89834 & ~n89835;
  assign n89839 = ~n89836 & n89838;
  assign n89840 = ~n89837 & n89839;
  assign n89841 = P2_P1_INSTQUEUE_REG_11__3_ & n89703;
  assign n89842 = P2_P1_INSTQUEUE_REG_10__3_ & n89705;
  assign n89843 = P2_P1_INSTQUEUE_REG_9__3_ & n89707;
  assign n89844 = P2_P1_INSTQUEUE_REG_8__3_ & n89709;
  assign n89845 = ~n89841 & ~n89842;
  assign n89846 = ~n89843 & n89845;
  assign n89847 = ~n89844 & n89846;
  assign n89848 = n89826 & n89833;
  assign n89849 = n89840 & n89848;
  assign n89850 = n89847 & n89849;
  assign n89851 = n89217 & ~n89850;
  assign n89852 = ~n83670 & n89718;
  assign n89853 = P2_P1_EAX_REG_19_ & ~n89216;
  assign n89854 = P2_P1_EAX_REG_18_ & n89810;
  assign n89855 = ~P2_P1_EAX_REG_19_ & n89854;
  assign n89856 = P2_P1_EAX_REG_19_ & ~n89854;
  assign n89857 = ~n89855 & ~n89856;
  assign n89858 = n89223 & ~n89857;
  assign n89859 = ~n83684 & n89726;
  assign n89860 = ~n89851 & ~n89852;
  assign n89861 = ~n89853 & n89860;
  assign n89862 = ~n89858 & n89861;
  assign n16261 = n89859 | ~n89862;
  assign n89864 = P2_P1_INSTQUEUE_REG_7__4_ & n89667;
  assign n89865 = P2_P1_INSTQUEUE_REG_6__4_ & n89669;
  assign n89866 = P2_P1_INSTQUEUE_REG_5__4_ & n89671;
  assign n89867 = P2_P1_INSTQUEUE_REG_4__4_ & n89673;
  assign n89868 = ~n89864 & ~n89865;
  assign n89869 = ~n89866 & n89868;
  assign n89870 = ~n89867 & n89869;
  assign n89871 = P2_P1_INSTQUEUE_REG_3__4_ & n89679;
  assign n89872 = P2_P1_INSTQUEUE_REG_2__4_ & n89681;
  assign n89873 = P2_P1_INSTQUEUE_REG_1__4_ & n89683;
  assign n89874 = P2_P1_INSTQUEUE_REG_0__4_ & n89685;
  assign n89875 = ~n89871 & ~n89872;
  assign n89876 = ~n89873 & n89875;
  assign n89877 = ~n89874 & n89876;
  assign n89878 = P2_P1_INSTQUEUE_REG_15__4_ & n89691;
  assign n89879 = P2_P1_INSTQUEUE_REG_14__4_ & n89693;
  assign n89880 = P2_P1_INSTQUEUE_REG_13__4_ & n89695;
  assign n89881 = P2_P1_INSTQUEUE_REG_12__4_ & n89697;
  assign n89882 = ~n89878 & ~n89879;
  assign n89883 = ~n89880 & n89882;
  assign n89884 = ~n89881 & n89883;
  assign n89885 = P2_P1_INSTQUEUE_REG_11__4_ & n89703;
  assign n89886 = P2_P1_INSTQUEUE_REG_10__4_ & n89705;
  assign n89887 = P2_P1_INSTQUEUE_REG_9__4_ & n89707;
  assign n89888 = P2_P1_INSTQUEUE_REG_8__4_ & n89709;
  assign n89889 = ~n89885 & ~n89886;
  assign n89890 = ~n89887 & n89889;
  assign n89891 = ~n89888 & n89890;
  assign n89892 = n89870 & n89877;
  assign n89893 = n89884 & n89892;
  assign n89894 = n89891 & n89893;
  assign n89895 = n89217 & ~n89894;
  assign n89896 = ~n83626 & n89718;
  assign n89897 = P2_P1_EAX_REG_20_ & ~n89216;
  assign n89898 = P2_P1_EAX_REG_19_ & n89854;
  assign n89899 = ~P2_P1_EAX_REG_20_ & n89898;
  assign n89900 = P2_P1_EAX_REG_20_ & ~n89898;
  assign n89901 = ~n89899 & ~n89900;
  assign n89902 = n89223 & ~n89901;
  assign n89903 = ~n83641 & n89726;
  assign n89904 = ~n89895 & ~n89896;
  assign n89905 = ~n89897 & n89904;
  assign n89906 = ~n89902 & n89905;
  assign n16266 = n89903 | ~n89906;
  assign n89908 = P2_P1_INSTQUEUE_REG_7__5_ & n89667;
  assign n89909 = P2_P1_INSTQUEUE_REG_6__5_ & n89669;
  assign n89910 = P2_P1_INSTQUEUE_REG_5__5_ & n89671;
  assign n89911 = P2_P1_INSTQUEUE_REG_4__5_ & n89673;
  assign n89912 = ~n89908 & ~n89909;
  assign n89913 = ~n89910 & n89912;
  assign n89914 = ~n89911 & n89913;
  assign n89915 = P2_P1_INSTQUEUE_REG_3__5_ & n89679;
  assign n89916 = P2_P1_INSTQUEUE_REG_2__5_ & n89681;
  assign n89917 = P2_P1_INSTQUEUE_REG_1__5_ & n89683;
  assign n89918 = P2_P1_INSTQUEUE_REG_0__5_ & n89685;
  assign n89919 = ~n89915 & ~n89916;
  assign n89920 = ~n89917 & n89919;
  assign n89921 = ~n89918 & n89920;
  assign n89922 = P2_P1_INSTQUEUE_REG_15__5_ & n89691;
  assign n89923 = P2_P1_INSTQUEUE_REG_14__5_ & n89693;
  assign n89924 = P2_P1_INSTQUEUE_REG_13__5_ & n89695;
  assign n89925 = P2_P1_INSTQUEUE_REG_12__5_ & n89697;
  assign n89926 = ~n89922 & ~n89923;
  assign n89927 = ~n89924 & n89926;
  assign n89928 = ~n89925 & n89927;
  assign n89929 = P2_P1_INSTQUEUE_REG_11__5_ & n89703;
  assign n89930 = P2_P1_INSTQUEUE_REG_10__5_ & n89705;
  assign n89931 = P2_P1_INSTQUEUE_REG_9__5_ & n89707;
  assign n89932 = P2_P1_INSTQUEUE_REG_8__5_ & n89709;
  assign n89933 = ~n89929 & ~n89930;
  assign n89934 = ~n89931 & n89933;
  assign n89935 = ~n89932 & n89934;
  assign n89936 = n89914 & n89921;
  assign n89937 = n89928 & n89936;
  assign n89938 = n89935 & n89937;
  assign n89939 = n89217 & ~n89938;
  assign n89940 = ~n83582 & n89718;
  assign n89941 = P2_P1_EAX_REG_21_ & ~n89216;
  assign n89942 = P2_P1_EAX_REG_20_ & n89898;
  assign n89943 = ~P2_P1_EAX_REG_21_ & n89942;
  assign n89944 = P2_P1_EAX_REG_21_ & ~n89942;
  assign n89945 = ~n89943 & ~n89944;
  assign n89946 = n89223 & ~n89945;
  assign n89947 = ~n83595 & n89726;
  assign n89948 = ~n89939 & ~n89940;
  assign n89949 = ~n89941 & n89948;
  assign n89950 = ~n89946 & n89949;
  assign n16271 = n89947 | ~n89950;
  assign n89952 = P2_P1_INSTQUEUE_REG_7__6_ & n89667;
  assign n89953 = P2_P1_INSTQUEUE_REG_6__6_ & n89669;
  assign n89954 = P2_P1_INSTQUEUE_REG_5__6_ & n89671;
  assign n89955 = P2_P1_INSTQUEUE_REG_4__6_ & n89673;
  assign n89956 = ~n89952 & ~n89953;
  assign n89957 = ~n89954 & n89956;
  assign n89958 = ~n89955 & n89957;
  assign n89959 = P2_P1_INSTQUEUE_REG_3__6_ & n89679;
  assign n89960 = P2_P1_INSTQUEUE_REG_2__6_ & n89681;
  assign n89961 = P2_P1_INSTQUEUE_REG_1__6_ & n89683;
  assign n89962 = P2_P1_INSTQUEUE_REG_0__6_ & n89685;
  assign n89963 = ~n89959 & ~n89960;
  assign n89964 = ~n89961 & n89963;
  assign n89965 = ~n89962 & n89964;
  assign n89966 = P2_P1_INSTQUEUE_REG_15__6_ & n89691;
  assign n89967 = P2_P1_INSTQUEUE_REG_14__6_ & n89693;
  assign n89968 = P2_P1_INSTQUEUE_REG_13__6_ & n89695;
  assign n89969 = P2_P1_INSTQUEUE_REG_12__6_ & n89697;
  assign n89970 = ~n89966 & ~n89967;
  assign n89971 = ~n89968 & n89970;
  assign n89972 = ~n89969 & n89971;
  assign n89973 = P2_P1_INSTQUEUE_REG_11__6_ & n89703;
  assign n89974 = P2_P1_INSTQUEUE_REG_10__6_ & n89705;
  assign n89975 = P2_P1_INSTQUEUE_REG_9__6_ & n89707;
  assign n89976 = P2_P1_INSTQUEUE_REG_8__6_ & n89709;
  assign n89977 = ~n89973 & ~n89974;
  assign n89978 = ~n89975 & n89977;
  assign n89979 = ~n89976 & n89978;
  assign n89980 = n89958 & n89965;
  assign n89981 = n89972 & n89980;
  assign n89982 = n89979 & n89981;
  assign n89983 = n89217 & ~n89982;
  assign n89984 = ~n83535 & n89718;
  assign n89985 = P2_P1_EAX_REG_22_ & ~n89216;
  assign n89986 = P2_P1_EAX_REG_21_ & n89942;
  assign n89987 = ~P2_P1_EAX_REG_22_ & n89986;
  assign n89988 = P2_P1_EAX_REG_22_ & ~n89986;
  assign n89989 = ~n89987 & ~n89988;
  assign n89990 = n89223 & ~n89989;
  assign n89991 = ~n83551 & n89726;
  assign n89992 = ~n89983 & ~n89984;
  assign n89993 = ~n89985 & n89992;
  assign n89994 = ~n89990 & n89993;
  assign n16276 = n89991 | ~n89994;
  assign n89996 = P2_P1_INSTQUEUERD_ADDR_REG_3_ & ~P2_P1_INSTQUEUERD_ADDR_REG_2_;
  assign n89997 = ~n76707 & ~n89996;
  assign n89998 = n76678 & n89997;
  assign n89999 = P2_P1_INSTQUEUE_REG_7__0_ & n89998;
  assign n90000 = n76682 & n89997;
  assign n90001 = P2_P1_INSTQUEUE_REG_6__0_ & n90000;
  assign n90002 = n76687 & n89997;
  assign n90003 = P2_P1_INSTQUEUE_REG_5__0_ & n90002;
  assign n90004 = n76691 & n89997;
  assign n90005 = P2_P1_INSTQUEUE_REG_4__0_ & n90004;
  assign n90006 = ~n89999 & ~n90001;
  assign n90007 = ~n90003 & n90006;
  assign n90008 = ~n90005 & n90007;
  assign n90009 = P2_P1_INSTQUEUERD_ADDR_REG_2_ & n89997;
  assign n90010 = n76677 & n90009;
  assign n90011 = P2_P1_INSTQUEUE_REG_3__0_ & n90010;
  assign n90012 = n76681 & n90009;
  assign n90013 = P2_P1_INSTQUEUE_REG_2__0_ & n90012;
  assign n90014 = n76686 & n90009;
  assign n90015 = P2_P1_INSTQUEUE_REG_1__0_ & n90014;
  assign n90016 = n76690 & n90009;
  assign n90017 = P2_P1_INSTQUEUE_REG_0__0_ & n90016;
  assign n90018 = ~n90011 & ~n90013;
  assign n90019 = ~n90015 & n90018;
  assign n90020 = ~n90017 & n90019;
  assign n90021 = n76678 & ~n89997;
  assign n90022 = P2_P1_INSTQUEUE_REG_15__0_ & n90021;
  assign n90023 = n76682 & ~n89997;
  assign n90024 = P2_P1_INSTQUEUE_REG_14__0_ & n90023;
  assign n90025 = n76687 & ~n89997;
  assign n90026 = P2_P1_INSTQUEUE_REG_13__0_ & n90025;
  assign n90027 = n76691 & ~n89997;
  assign n90028 = P2_P1_INSTQUEUE_REG_12__0_ & n90027;
  assign n90029 = ~n90022 & ~n90024;
  assign n90030 = ~n90026 & n90029;
  assign n90031 = ~n90028 & n90030;
  assign n90032 = P2_P1_INSTQUEUERD_ADDR_REG_2_ & ~n89997;
  assign n90033 = n76677 & n90032;
  assign n90034 = P2_P1_INSTQUEUE_REG_11__0_ & n90033;
  assign n90035 = n76681 & n90032;
  assign n90036 = P2_P1_INSTQUEUE_REG_10__0_ & n90035;
  assign n90037 = n76686 & n90032;
  assign n90038 = P2_P1_INSTQUEUE_REG_9__0_ & n90037;
  assign n90039 = n76690 & n90032;
  assign n90040 = P2_P1_INSTQUEUE_REG_8__0_ & n90039;
  assign n90041 = ~n90034 & ~n90036;
  assign n90042 = ~n90038 & n90041;
  assign n90043 = ~n90040 & n90042;
  assign n90044 = n90008 & n90020;
  assign n90045 = n90031 & n90044;
  assign n90046 = n90043 & n90045;
  assign n90047 = P2_P1_INSTQUEUE_REG_7__7_ & n89667;
  assign n90048 = P2_P1_INSTQUEUE_REG_6__7_ & n89669;
  assign n90049 = P2_P1_INSTQUEUE_REG_5__7_ & n89671;
  assign n90050 = P2_P1_INSTQUEUE_REG_4__7_ & n89673;
  assign n90051 = ~n90047 & ~n90048;
  assign n90052 = ~n90049 & n90051;
  assign n90053 = ~n90050 & n90052;
  assign n90054 = P2_P1_INSTQUEUE_REG_3__7_ & n89679;
  assign n90055 = P2_P1_INSTQUEUE_REG_2__7_ & n89681;
  assign n90056 = P2_P1_INSTQUEUE_REG_1__7_ & n89683;
  assign n90057 = P2_P1_INSTQUEUE_REG_0__7_ & n89685;
  assign n90058 = ~n90054 & ~n90055;
  assign n90059 = ~n90056 & n90058;
  assign n90060 = ~n90057 & n90059;
  assign n90061 = P2_P1_INSTQUEUE_REG_15__7_ & n89691;
  assign n90062 = P2_P1_INSTQUEUE_REG_14__7_ & n89693;
  assign n90063 = P2_P1_INSTQUEUE_REG_13__7_ & n89695;
  assign n90064 = P2_P1_INSTQUEUE_REG_12__7_ & n89697;
  assign n90065 = ~n90061 & ~n90062;
  assign n90066 = ~n90063 & n90065;
  assign n90067 = ~n90064 & n90066;
  assign n90068 = P2_P1_INSTQUEUE_REG_11__7_ & n89703;
  assign n90069 = P2_P1_INSTQUEUE_REG_10__7_ & n89705;
  assign n90070 = P2_P1_INSTQUEUE_REG_9__7_ & n89707;
  assign n90071 = P2_P1_INSTQUEUE_REG_8__7_ & n89709;
  assign n90072 = ~n90068 & ~n90069;
  assign n90073 = ~n90070 & n90072;
  assign n90074 = ~n90071 & n90073;
  assign n90075 = n90053 & n90060;
  assign n90076 = n90067 & n90075;
  assign n90077 = n90074 & n90076;
  assign n90078 = ~n90046 & n90077;
  assign n90079 = n90046 & ~n90077;
  assign n90080 = ~n90078 & ~n90079;
  assign n90081 = n89217 & ~n90080;
  assign n90082 = ~n77700 & n89718;
  assign n90083 = P2_P1_EAX_REG_23_ & ~n89216;
  assign n90084 = P2_P1_EAX_REG_22_ & n89986;
  assign n90085 = ~P2_P1_EAX_REG_23_ & n90084;
  assign n90086 = P2_P1_EAX_REG_23_ & ~n90084;
  assign n90087 = ~n90085 & ~n90086;
  assign n90088 = n89223 & ~n90087;
  assign n90089 = ~n80591 & n89726;
  assign n90090 = ~n90081 & ~n90082;
  assign n90091 = ~n90083 & n90090;
  assign n90092 = ~n90088 & n90091;
  assign n16281 = n90089 | ~n90092;
  assign n90094 = ~n90046 & ~n90077;
  assign n90095 = P2_P1_INSTQUEUE_REG_7__1_ & n89998;
  assign n90096 = P2_P1_INSTQUEUE_REG_6__1_ & n90000;
  assign n90097 = P2_P1_INSTQUEUE_REG_5__1_ & n90002;
  assign n90098 = P2_P1_INSTQUEUE_REG_4__1_ & n90004;
  assign n90099 = ~n90095 & ~n90096;
  assign n90100 = ~n90097 & n90099;
  assign n90101 = ~n90098 & n90100;
  assign n90102 = P2_P1_INSTQUEUE_REG_3__1_ & n90010;
  assign n90103 = P2_P1_INSTQUEUE_REG_2__1_ & n90012;
  assign n90104 = P2_P1_INSTQUEUE_REG_1__1_ & n90014;
  assign n90105 = P2_P1_INSTQUEUE_REG_0__1_ & n90016;
  assign n90106 = ~n90102 & ~n90103;
  assign n90107 = ~n90104 & n90106;
  assign n90108 = ~n90105 & n90107;
  assign n90109 = P2_P1_INSTQUEUE_REG_15__1_ & n90021;
  assign n90110 = P2_P1_INSTQUEUE_REG_14__1_ & n90023;
  assign n90111 = P2_P1_INSTQUEUE_REG_13__1_ & n90025;
  assign n90112 = P2_P1_INSTQUEUE_REG_12__1_ & n90027;
  assign n90113 = ~n90109 & ~n90110;
  assign n90114 = ~n90111 & n90113;
  assign n90115 = ~n90112 & n90114;
  assign n90116 = P2_P1_INSTQUEUE_REG_11__1_ & n90033;
  assign n90117 = P2_P1_INSTQUEUE_REG_10__1_ & n90035;
  assign n90118 = P2_P1_INSTQUEUE_REG_9__1_ & n90037;
  assign n90119 = P2_P1_INSTQUEUE_REG_8__1_ & n90039;
  assign n90120 = ~n90116 & ~n90117;
  assign n90121 = ~n90118 & n90120;
  assign n90122 = ~n90119 & n90121;
  assign n90123 = n90101 & n90108;
  assign n90124 = n90115 & n90123;
  assign n90125 = n90122 & n90124;
  assign n90126 = n90094 & n90125;
  assign n90127 = ~n90094 & ~n90125;
  assign n90128 = ~n90126 & ~n90127;
  assign n90129 = n89217 & ~n90128;
  assign n90130 = ~n88948 & n89718;
  assign n90131 = P2_P1_EAX_REG_24_ & ~n89216;
  assign n90132 = P2_P1_EAX_REG_23_ & n90084;
  assign n90133 = ~P2_P1_EAX_REG_24_ & n90132;
  assign n90134 = P2_P1_EAX_REG_24_ & ~n90132;
  assign n90135 = ~n90133 & ~n90134;
  assign n90136 = n89223 & ~n90135;
  assign n90137 = ~n83819 & n89726;
  assign n90138 = ~n90129 & ~n90130;
  assign n90139 = ~n90131 & n90138;
  assign n90140 = ~n90136 & n90139;
  assign n16286 = n90137 | ~n90140;
  assign n90142 = n90094 & ~n90125;
  assign n90143 = P2_P1_INSTQUEUE_REG_7__2_ & n89998;
  assign n90144 = P2_P1_INSTQUEUE_REG_6__2_ & n90000;
  assign n90145 = P2_P1_INSTQUEUE_REG_5__2_ & n90002;
  assign n90146 = P2_P1_INSTQUEUE_REG_4__2_ & n90004;
  assign n90147 = ~n90143 & ~n90144;
  assign n90148 = ~n90145 & n90147;
  assign n90149 = ~n90146 & n90148;
  assign n90150 = P2_P1_INSTQUEUE_REG_3__2_ & n90010;
  assign n90151 = P2_P1_INSTQUEUE_REG_2__2_ & n90012;
  assign n90152 = P2_P1_INSTQUEUE_REG_1__2_ & n90014;
  assign n90153 = P2_P1_INSTQUEUE_REG_0__2_ & n90016;
  assign n90154 = ~n90150 & ~n90151;
  assign n90155 = ~n90152 & n90154;
  assign n90156 = ~n90153 & n90155;
  assign n90157 = P2_P1_INSTQUEUE_REG_15__2_ & n90021;
  assign n90158 = P2_P1_INSTQUEUE_REG_14__2_ & n90023;
  assign n90159 = P2_P1_INSTQUEUE_REG_13__2_ & n90025;
  assign n90160 = P2_P1_INSTQUEUE_REG_12__2_ & n90027;
  assign n90161 = ~n90157 & ~n90158;
  assign n90162 = ~n90159 & n90161;
  assign n90163 = ~n90160 & n90162;
  assign n90164 = P2_P1_INSTQUEUE_REG_11__2_ & n90033;
  assign n90165 = P2_P1_INSTQUEUE_REG_10__2_ & n90035;
  assign n90166 = P2_P1_INSTQUEUE_REG_9__2_ & n90037;
  assign n90167 = P2_P1_INSTQUEUE_REG_8__2_ & n90039;
  assign n90168 = ~n90164 & ~n90165;
  assign n90169 = ~n90166 & n90168;
  assign n90170 = ~n90167 & n90169;
  assign n90171 = n90149 & n90156;
  assign n90172 = n90163 & n90171;
  assign n90173 = n90170 & n90172;
  assign n90174 = n90142 & n90173;
  assign n90175 = ~n90142 & ~n90173;
  assign n90176 = ~n90174 & ~n90175;
  assign n90177 = n89217 & ~n90176;
  assign n90178 = ~n88931 & n89718;
  assign n90179 = P2_P1_EAX_REG_25_ & ~n89216;
  assign n90180 = P2_P1_EAX_REG_24_ & n90132;
  assign n90181 = ~P2_P1_EAX_REG_25_ & n90180;
  assign n90182 = P2_P1_EAX_REG_25_ & ~n90180;
  assign n90183 = ~n90181 & ~n90182;
  assign n90184 = n89223 & ~n90183;
  assign n90185 = ~n83780 & n89726;
  assign n90186 = ~n90177 & ~n90178;
  assign n90187 = ~n90179 & n90186;
  assign n90188 = ~n90184 & n90187;
  assign n16291 = n90185 | ~n90188;
  assign n90190 = n90142 & ~n90173;
  assign n90191 = P2_P1_INSTQUEUE_REG_7__3_ & n89998;
  assign n90192 = P2_P1_INSTQUEUE_REG_6__3_ & n90000;
  assign n90193 = P2_P1_INSTQUEUE_REG_5__3_ & n90002;
  assign n90194 = P2_P1_INSTQUEUE_REG_4__3_ & n90004;
  assign n90195 = ~n90191 & ~n90192;
  assign n90196 = ~n90193 & n90195;
  assign n90197 = ~n90194 & n90196;
  assign n90198 = P2_P1_INSTQUEUE_REG_3__3_ & n90010;
  assign n90199 = P2_P1_INSTQUEUE_REG_2__3_ & n90012;
  assign n90200 = P2_P1_INSTQUEUE_REG_1__3_ & n90014;
  assign n90201 = P2_P1_INSTQUEUE_REG_0__3_ & n90016;
  assign n90202 = ~n90198 & ~n90199;
  assign n90203 = ~n90200 & n90202;
  assign n90204 = ~n90201 & n90203;
  assign n90205 = P2_P1_INSTQUEUE_REG_15__3_ & n90021;
  assign n90206 = P2_P1_INSTQUEUE_REG_14__3_ & n90023;
  assign n90207 = P2_P1_INSTQUEUE_REG_13__3_ & n90025;
  assign n90208 = P2_P1_INSTQUEUE_REG_12__3_ & n90027;
  assign n90209 = ~n90205 & ~n90206;
  assign n90210 = ~n90207 & n90209;
  assign n90211 = ~n90208 & n90210;
  assign n90212 = P2_P1_INSTQUEUE_REG_11__3_ & n90033;
  assign n90213 = P2_P1_INSTQUEUE_REG_10__3_ & n90035;
  assign n90214 = P2_P1_INSTQUEUE_REG_9__3_ & n90037;
  assign n90215 = P2_P1_INSTQUEUE_REG_8__3_ & n90039;
  assign n90216 = ~n90212 & ~n90213;
  assign n90217 = ~n90214 & n90216;
  assign n90218 = ~n90215 & n90217;
  assign n90219 = n90197 & n90204;
  assign n90220 = n90211 & n90219;
  assign n90221 = n90218 & n90220;
  assign n90222 = n90190 & n90221;
  assign n90223 = ~n90190 & ~n90221;
  assign n90224 = ~n90222 & ~n90223;
  assign n90225 = n89217 & ~n90224;
  assign n90226 = ~n88919 & n89718;
  assign n90227 = P2_P1_EAX_REG_26_ & ~n89216;
  assign n90228 = P2_P1_EAX_REG_25_ & n90180;
  assign n90229 = ~P2_P1_EAX_REG_26_ & n90228;
  assign n90230 = P2_P1_EAX_REG_26_ & ~n90228;
  assign n90231 = ~n90229 & ~n90230;
  assign n90232 = n89223 & ~n90231;
  assign n90233 = ~n83742 & n89726;
  assign n90234 = ~n90225 & ~n90226;
  assign n90235 = ~n90227 & n90234;
  assign n90236 = ~n90232 & n90235;
  assign n16296 = n90233 | ~n90236;
  assign n90238 = n90190 & ~n90221;
  assign n90239 = P2_P1_INSTQUEUE_REG_7__4_ & n89998;
  assign n90240 = P2_P1_INSTQUEUE_REG_6__4_ & n90000;
  assign n90241 = P2_P1_INSTQUEUE_REG_5__4_ & n90002;
  assign n90242 = P2_P1_INSTQUEUE_REG_4__4_ & n90004;
  assign n90243 = ~n90239 & ~n90240;
  assign n90244 = ~n90241 & n90243;
  assign n90245 = ~n90242 & n90244;
  assign n90246 = P2_P1_INSTQUEUE_REG_3__4_ & n90010;
  assign n90247 = P2_P1_INSTQUEUE_REG_2__4_ & n90012;
  assign n90248 = P2_P1_INSTQUEUE_REG_1__4_ & n90014;
  assign n90249 = P2_P1_INSTQUEUE_REG_0__4_ & n90016;
  assign n90250 = ~n90246 & ~n90247;
  assign n90251 = ~n90248 & n90250;
  assign n90252 = ~n90249 & n90251;
  assign n90253 = P2_P1_INSTQUEUE_REG_15__4_ & n90021;
  assign n90254 = P2_P1_INSTQUEUE_REG_14__4_ & n90023;
  assign n90255 = P2_P1_INSTQUEUE_REG_13__4_ & n90025;
  assign n90256 = P2_P1_INSTQUEUE_REG_12__4_ & n90027;
  assign n90257 = ~n90253 & ~n90254;
  assign n90258 = ~n90255 & n90257;
  assign n90259 = ~n90256 & n90258;
  assign n90260 = P2_P1_INSTQUEUE_REG_11__4_ & n90033;
  assign n90261 = P2_P1_INSTQUEUE_REG_10__4_ & n90035;
  assign n90262 = P2_P1_INSTQUEUE_REG_9__4_ & n90037;
  assign n90263 = P2_P1_INSTQUEUE_REG_8__4_ & n90039;
  assign n90264 = ~n90260 & ~n90261;
  assign n90265 = ~n90262 & n90264;
  assign n90266 = ~n90263 & n90265;
  assign n90267 = n90245 & n90252;
  assign n90268 = n90259 & n90267;
  assign n90269 = n90266 & n90268;
  assign n90270 = n90238 & n90269;
  assign n90271 = ~n90238 & ~n90269;
  assign n90272 = ~n90270 & ~n90271;
  assign n90273 = n89217 & ~n90272;
  assign n90274 = ~n88903 & n89718;
  assign n90275 = P2_P1_EAX_REG_27_ & ~n89216;
  assign n90276 = P2_P1_EAX_REG_26_ & n90228;
  assign n90277 = ~P2_P1_EAX_REG_27_ & n90276;
  assign n90278 = P2_P1_EAX_REG_27_ & ~n90276;
  assign n90279 = ~n90277 & ~n90278;
  assign n90280 = n89223 & ~n90279;
  assign n90281 = ~n90275 & ~n90280;
  assign n90282 = ~n83694 & n89726;
  assign n90283 = ~n90273 & ~n90274;
  assign n90284 = n90281 & n90283;
  assign n16301 = n90282 | ~n90284;
  assign n90286 = P2_P1_EAX_REG_28_ & ~n89216;
  assign n90287 = P2_P1_EAX_REG_27_ & n90276;
  assign n90288 = ~P2_P1_EAX_REG_28_ & n90287;
  assign n90289 = P2_P1_EAX_REG_28_ & ~n90287;
  assign n90290 = ~n90288 & ~n90289;
  assign n90291 = n89223 & ~n90290;
  assign n90292 = n90238 & ~n90269;
  assign n90293 = P2_P1_INSTQUEUE_REG_7__5_ & n89998;
  assign n90294 = P2_P1_INSTQUEUE_REG_6__5_ & n90000;
  assign n90295 = P2_P1_INSTQUEUE_REG_5__5_ & n90002;
  assign n90296 = P2_P1_INSTQUEUE_REG_4__5_ & n90004;
  assign n90297 = ~n90293 & ~n90294;
  assign n90298 = ~n90295 & n90297;
  assign n90299 = ~n90296 & n90298;
  assign n90300 = P2_P1_INSTQUEUE_REG_3__5_ & n90010;
  assign n90301 = P2_P1_INSTQUEUE_REG_2__5_ & n90012;
  assign n90302 = P2_P1_INSTQUEUE_REG_1__5_ & n90014;
  assign n90303 = P2_P1_INSTQUEUE_REG_0__5_ & n90016;
  assign n90304 = ~n90300 & ~n90301;
  assign n90305 = ~n90302 & n90304;
  assign n90306 = ~n90303 & n90305;
  assign n90307 = P2_P1_INSTQUEUE_REG_15__5_ & n90021;
  assign n90308 = P2_P1_INSTQUEUE_REG_14__5_ & n90023;
  assign n90309 = P2_P1_INSTQUEUE_REG_13__5_ & n90025;
  assign n90310 = P2_P1_INSTQUEUE_REG_12__5_ & n90027;
  assign n90311 = ~n90307 & ~n90308;
  assign n90312 = ~n90309 & n90311;
  assign n90313 = ~n90310 & n90312;
  assign n90314 = P2_P1_INSTQUEUE_REG_11__5_ & n90033;
  assign n90315 = P2_P1_INSTQUEUE_REG_10__5_ & n90035;
  assign n90316 = P2_P1_INSTQUEUE_REG_9__5_ & n90037;
  assign n90317 = P2_P1_INSTQUEUE_REG_8__5_ & n90039;
  assign n90318 = ~n90314 & ~n90315;
  assign n90319 = ~n90316 & n90318;
  assign n90320 = ~n90317 & n90319;
  assign n90321 = n90299 & n90306;
  assign n90322 = n90313 & n90321;
  assign n90323 = n90320 & n90322;
  assign n90324 = n90292 & n90323;
  assign n90325 = ~n90292 & ~n90323;
  assign n90326 = ~n90324 & ~n90325;
  assign n90327 = n89217 & ~n90326;
  assign n90328 = ~n90286 & ~n90291;
  assign n90329 = ~n90327 & n90328;
  assign n90330 = ~n88888 & n89718;
  assign n90331 = ~n83653 & n89726;
  assign n90332 = n90329 & ~n90330;
  assign n16306 = n90331 | ~n90332;
  assign n90334 = P2_P1_EAX_REG_29_ & ~n89216;
  assign n90335 = P2_P1_EAX_REG_28_ & n90287;
  assign n90336 = ~P2_P1_EAX_REG_29_ & n90335;
  assign n90337 = P2_P1_EAX_REG_29_ & ~n90335;
  assign n90338 = ~n90336 & ~n90337;
  assign n90339 = n89223 & ~n90338;
  assign n90340 = n90292 & ~n90323;
  assign n90341 = P2_P1_INSTQUEUE_REG_7__6_ & n89998;
  assign n90342 = P2_P1_INSTQUEUE_REG_6__6_ & n90000;
  assign n90343 = P2_P1_INSTQUEUE_REG_5__6_ & n90002;
  assign n90344 = P2_P1_INSTQUEUE_REG_4__6_ & n90004;
  assign n90345 = ~n90341 & ~n90342;
  assign n90346 = ~n90343 & n90345;
  assign n90347 = ~n90344 & n90346;
  assign n90348 = P2_P1_INSTQUEUE_REG_3__6_ & n90010;
  assign n90349 = P2_P1_INSTQUEUE_REG_2__6_ & n90012;
  assign n90350 = P2_P1_INSTQUEUE_REG_1__6_ & n90014;
  assign n90351 = P2_P1_INSTQUEUE_REG_0__6_ & n90016;
  assign n90352 = ~n90348 & ~n90349;
  assign n90353 = ~n90350 & n90352;
  assign n90354 = ~n90351 & n90353;
  assign n90355 = P2_P1_INSTQUEUE_REG_15__6_ & n90021;
  assign n90356 = P2_P1_INSTQUEUE_REG_14__6_ & n90023;
  assign n90357 = P2_P1_INSTQUEUE_REG_13__6_ & n90025;
  assign n90358 = P2_P1_INSTQUEUE_REG_12__6_ & n90027;
  assign n90359 = ~n90355 & ~n90356;
  assign n90360 = ~n90357 & n90359;
  assign n90361 = ~n90358 & n90360;
  assign n90362 = P2_P1_INSTQUEUE_REG_11__6_ & n90033;
  assign n90363 = P2_P1_INSTQUEUE_REG_10__6_ & n90035;
  assign n90364 = P2_P1_INSTQUEUE_REG_9__6_ & n90037;
  assign n90365 = P2_P1_INSTQUEUE_REG_8__6_ & n90039;
  assign n90366 = ~n90362 & ~n90363;
  assign n90367 = ~n90364 & n90366;
  assign n90368 = ~n90365 & n90367;
  assign n90369 = n90347 & n90354;
  assign n90370 = n90361 & n90369;
  assign n90371 = n90368 & n90370;
  assign n90372 = n90340 & n90371;
  assign n90373 = ~n90340 & ~n90371;
  assign n90374 = ~n90372 & ~n90373;
  assign n90375 = n89217 & ~n90374;
  assign n90376 = ~n90334 & ~n90339;
  assign n90377 = ~n90375 & n90376;
  assign n90378 = ~n88872 & n89718;
  assign n90379 = ~n83607 & n89726;
  assign n90380 = n90377 & ~n90378;
  assign n16311 = n90379 | ~n90380;
  assign n90382 = P2_P1_EAX_REG_30_ & ~n89216;
  assign n90383 = P2_P1_EAX_REG_29_ & n90335;
  assign n90384 = ~P2_P1_EAX_REG_30_ & n90383;
  assign n90385 = P2_P1_EAX_REG_30_ & ~n90383;
  assign n90386 = ~n90384 & ~n90385;
  assign n90387 = n89223 & ~n90386;
  assign n90388 = n90340 & ~n90371;
  assign n90389 = P2_P1_INSTQUEUE_REG_7__7_ & n89998;
  assign n90390 = P2_P1_INSTQUEUE_REG_6__7_ & n90000;
  assign n90391 = P2_P1_INSTQUEUE_REG_5__7_ & n90002;
  assign n90392 = P2_P1_INSTQUEUE_REG_4__7_ & n90004;
  assign n90393 = ~n90389 & ~n90390;
  assign n90394 = ~n90391 & n90393;
  assign n90395 = ~n90392 & n90394;
  assign n90396 = P2_P1_INSTQUEUE_REG_3__7_ & n90010;
  assign n90397 = P2_P1_INSTQUEUE_REG_2__7_ & n90012;
  assign n90398 = P2_P1_INSTQUEUE_REG_1__7_ & n90014;
  assign n90399 = P2_P1_INSTQUEUE_REG_0__7_ & n90016;
  assign n90400 = ~n90396 & ~n90397;
  assign n90401 = ~n90398 & n90400;
  assign n90402 = ~n90399 & n90401;
  assign n90403 = P2_P1_INSTQUEUE_REG_15__7_ & n90021;
  assign n90404 = P2_P1_INSTQUEUE_REG_14__7_ & n90023;
  assign n90405 = P2_P1_INSTQUEUE_REG_13__7_ & n90025;
  assign n90406 = P2_P1_INSTQUEUE_REG_12__7_ & n90027;
  assign n90407 = ~n90403 & ~n90404;
  assign n90408 = ~n90405 & n90407;
  assign n90409 = ~n90406 & n90408;
  assign n90410 = P2_P1_INSTQUEUE_REG_11__7_ & n90033;
  assign n90411 = P2_P1_INSTQUEUE_REG_10__7_ & n90035;
  assign n90412 = P2_P1_INSTQUEUE_REG_9__7_ & n90037;
  assign n90413 = P2_P1_INSTQUEUE_REG_8__7_ & n90039;
  assign n90414 = ~n90410 & ~n90411;
  assign n90415 = ~n90412 & n90414;
  assign n90416 = ~n90413 & n90415;
  assign n90417 = n90395 & n90402;
  assign n90418 = n90409 & n90417;
  assign n90419 = n90416 & n90418;
  assign n90420 = n90388 & n90419;
  assign n90421 = ~n90388 & ~n90419;
  assign n90422 = ~n90420 & ~n90421;
  assign n90423 = n89217 & ~n90422;
  assign n90424 = ~n90382 & ~n90387;
  assign n90425 = ~n90423 & n90424;
  assign n90426 = ~n88858 & n89718;
  assign n90427 = ~n83565 & n89726;
  assign n90428 = n90425 & ~n90426;
  assign n16316 = n90427 | ~n90428;
  assign n90430 = P2_P1_EAX_REG_30_ & n90383;
  assign n90431 = ~P2_P1_EAX_REG_31_ & n90430;
  assign n90432 = P2_P1_EAX_REG_31_ & ~n90430;
  assign n90433 = ~n90431 & ~n90432;
  assign n90434 = n89223 & ~n90433;
  assign n90435 = P2_P1_EAX_REG_31_ & ~n89216;
  assign n90436 = ~n90434 & ~n90435;
  assign n90437 = ~n83518 & n89726;
  assign n16321 = ~n90436 | n90437;
  assign n90439 = ~n77098 & ~n77192;
  assign n90440 = n77311 & ~n90439;
  assign n90441 = n76828 & n90440;
  assign n90442 = ~P2_P1_EBX_REG_0_ & n90441;
  assign n90443 = ~n76828 & n90440;
  assign n90444 = P2_P1_INSTQUEUE_REG_0__0_ & n90443;
  assign n90445 = P2_P1_EBX_REG_0_ & ~n90440;
  assign n90446 = ~n90442 & ~n90444;
  assign n16326 = n90445 | ~n90446;
  assign n90448 = ~P2_P1_EBX_REG_0_ & P2_P1_EBX_REG_1_;
  assign n90449 = P2_P1_EBX_REG_0_ & ~P2_P1_EBX_REG_1_;
  assign n90450 = ~n90448 & ~n90449;
  assign n90451 = n90441 & ~n90450;
  assign n90452 = P2_P1_INSTQUEUE_REG_0__1_ & n90443;
  assign n90453 = P2_P1_EBX_REG_1_ & ~n90440;
  assign n90454 = ~n90451 & ~n90452;
  assign n16331 = n90453 | ~n90454;
  assign n90456 = P2_P1_EBX_REG_0_ & P2_P1_EBX_REG_1_;
  assign n90457 = ~P2_P1_EBX_REG_2_ & n90456;
  assign n90458 = P2_P1_EBX_REG_2_ & ~n90456;
  assign n90459 = ~n90457 & ~n90458;
  assign n90460 = n90441 & ~n90459;
  assign n90461 = P2_P1_INSTQUEUE_REG_0__2_ & n90443;
  assign n90462 = P2_P1_EBX_REG_2_ & ~n90440;
  assign n90463 = ~n90460 & ~n90461;
  assign n16336 = n90462 | ~n90463;
  assign n90465 = P2_P1_EBX_REG_0_ & P2_P1_EBX_REG_2_;
  assign n90466 = P2_P1_EBX_REG_1_ & n90465;
  assign n90467 = P2_P1_EBX_REG_3_ & ~n90466;
  assign n90468 = ~P2_P1_EBX_REG_3_ & n90466;
  assign n90469 = ~n90467 & ~n90468;
  assign n90470 = n90441 & ~n90469;
  assign n90471 = P2_P1_INSTQUEUE_REG_0__3_ & n90443;
  assign n90472 = P2_P1_EBX_REG_3_ & ~n90440;
  assign n90473 = ~n90470 & ~n90471;
  assign n16341 = n90472 | ~n90473;
  assign n90475 = P2_P1_EBX_REG_3_ & n90466;
  assign n90476 = ~P2_P1_EBX_REG_4_ & n90475;
  assign n90477 = P2_P1_EBX_REG_4_ & ~n90475;
  assign n90478 = ~n90476 & ~n90477;
  assign n90479 = n90441 & ~n90478;
  assign n90480 = P2_P1_INSTQUEUE_REG_0__4_ & n90443;
  assign n90481 = P2_P1_EBX_REG_4_ & ~n90440;
  assign n90482 = ~n90479 & ~n90480;
  assign n16346 = n90481 | ~n90482;
  assign n90484 = P2_P1_EBX_REG_3_ & P2_P1_EBX_REG_4_;
  assign n90485 = n90466 & n90484;
  assign n90486 = P2_P1_EBX_REG_5_ & ~n90485;
  assign n90487 = ~P2_P1_EBX_REG_5_ & n90485;
  assign n90488 = ~n90486 & ~n90487;
  assign n90489 = n90441 & ~n90488;
  assign n90490 = P2_P1_INSTQUEUE_REG_0__5_ & n90443;
  assign n90491 = P2_P1_EBX_REG_5_ & ~n90440;
  assign n90492 = ~n90489 & ~n90490;
  assign n16351 = n90491 | ~n90492;
  assign n90494 = P2_P1_EBX_REG_5_ & n90485;
  assign n90495 = ~P2_P1_EBX_REG_6_ & n90494;
  assign n90496 = P2_P1_EBX_REG_6_ & ~n90494;
  assign n90497 = ~n90495 & ~n90496;
  assign n90498 = n90441 & ~n90497;
  assign n90499 = P2_P1_INSTQUEUE_REG_0__6_ & n90443;
  assign n90500 = P2_P1_EBX_REG_6_ & ~n90440;
  assign n90501 = ~n90498 & ~n90499;
  assign n16356 = n90500 | ~n90501;
  assign n90503 = P2_P1_EBX_REG_5_ & P2_P1_EBX_REG_6_;
  assign n90504 = n90485 & n90503;
  assign n90505 = P2_P1_EBX_REG_7_ & ~n90504;
  assign n90506 = ~P2_P1_EBX_REG_7_ & n90504;
  assign n90507 = ~n90505 & ~n90506;
  assign n90508 = n90441 & ~n90507;
  assign n90509 = P2_P1_INSTQUEUE_REG_0__7_ & n90443;
  assign n90510 = P2_P1_EBX_REG_7_ & ~n90440;
  assign n90511 = ~n90508 & ~n90509;
  assign n16361 = n90510 | ~n90511;
  assign n90513 = P2_P1_EBX_REG_7_ & n90504;
  assign n90514 = ~P2_P1_EBX_REG_8_ & n90513;
  assign n90515 = P2_P1_EBX_REG_8_ & ~n90513;
  assign n90516 = ~n90514 & ~n90515;
  assign n90517 = n90441 & ~n90516;
  assign n90518 = ~n89362 & n90443;
  assign n90519 = P2_P1_EBX_REG_8_ & ~n90440;
  assign n90520 = ~n90517 & ~n90518;
  assign n16366 = n90519 | ~n90520;
  assign n90522 = P2_P1_EBX_REG_7_ & P2_P1_EBX_REG_8_;
  assign n90523 = n90504 & n90522;
  assign n90524 = P2_P1_EBX_REG_9_ & ~n90523;
  assign n90525 = ~P2_P1_EBX_REG_9_ & n90523;
  assign n90526 = ~n90524 & ~n90525;
  assign n90527 = n90441 & ~n90526;
  assign n90528 = ~n89404 & n90443;
  assign n90529 = P2_P1_EBX_REG_9_ & ~n90440;
  assign n90530 = ~n90527 & ~n90528;
  assign n16371 = n90529 | ~n90530;
  assign n90532 = P2_P1_EBX_REG_10_ & ~n90440;
  assign n90533 = ~n89446 & n90443;
  assign n90534 = P2_P1_EBX_REG_9_ & n90523;
  assign n90535 = ~P2_P1_EBX_REG_10_ & n90534;
  assign n90536 = P2_P1_EBX_REG_10_ & ~n90534;
  assign n90537 = ~n90535 & ~n90536;
  assign n90538 = n90441 & ~n90537;
  assign n90539 = ~n90532 & ~n90533;
  assign n16376 = n90538 | ~n90539;
  assign n90541 = P2_P1_EBX_REG_11_ & ~n90440;
  assign n90542 = ~n89488 & n90443;
  assign n90543 = P2_P1_EBX_REG_9_ & P2_P1_EBX_REG_10_;
  assign n90544 = n90523 & n90543;
  assign n90545 = P2_P1_EBX_REG_11_ & ~n90544;
  assign n90546 = ~P2_P1_EBX_REG_11_ & n90544;
  assign n90547 = ~n90545 & ~n90546;
  assign n90548 = n90441 & ~n90547;
  assign n90549 = ~n90541 & ~n90542;
  assign n16381 = n90548 | ~n90549;
  assign n90551 = P2_P1_EBX_REG_12_ & ~n90440;
  assign n90552 = ~n89525 & n90443;
  assign n90553 = P2_P1_EBX_REG_11_ & n90544;
  assign n90554 = ~P2_P1_EBX_REG_12_ & n90553;
  assign n90555 = P2_P1_EBX_REG_12_ & ~n90553;
  assign n90556 = ~n90554 & ~n90555;
  assign n90557 = n90441 & ~n90556;
  assign n90558 = ~n90551 & ~n90552;
  assign n16386 = n90557 | ~n90558;
  assign n90560 = P2_P1_EBX_REG_13_ & ~n90440;
  assign n90561 = ~n89567 & n90443;
  assign n90562 = P2_P1_EBX_REG_11_ & P2_P1_EBX_REG_12_;
  assign n90563 = n90544 & n90562;
  assign n90564 = P2_P1_EBX_REG_13_ & ~n90563;
  assign n90565 = ~P2_P1_EBX_REG_13_ & n90563;
  assign n90566 = ~n90564 & ~n90565;
  assign n90567 = n90441 & ~n90566;
  assign n90568 = ~n90560 & ~n90561;
  assign n16391 = n90567 | ~n90568;
  assign n90570 = P2_P1_EBX_REG_14_ & ~n90440;
  assign n90571 = ~n89609 & n90443;
  assign n90572 = P2_P1_EBX_REG_13_ & n90563;
  assign n90573 = ~P2_P1_EBX_REG_14_ & n90572;
  assign n90574 = P2_P1_EBX_REG_14_ & ~n90572;
  assign n90575 = ~n90573 & ~n90574;
  assign n90576 = n90441 & ~n90575;
  assign n90577 = ~n90570 & ~n90571;
  assign n16396 = n90576 | ~n90577;
  assign n90579 = P2_P1_EBX_REG_15_ & ~n90440;
  assign n90580 = ~n89651 & n90443;
  assign n90581 = P2_P1_EBX_REG_13_ & P2_P1_EBX_REG_14_;
  assign n90582 = n90563 & n90581;
  assign n90583 = P2_P1_EBX_REG_15_ & ~n90582;
  assign n90584 = ~P2_P1_EBX_REG_15_ & n90582;
  assign n90585 = ~n90583 & ~n90584;
  assign n90586 = n90441 & ~n90585;
  assign n90587 = ~n90579 & ~n90580;
  assign n16401 = n90586 | ~n90587;
  assign n90589 = P2_P1_EBX_REG_16_ & ~n90440;
  assign n90590 = ~n89716 & n90443;
  assign n90591 = P2_P1_EBX_REG_15_ & n90582;
  assign n90592 = ~P2_P1_EBX_REG_16_ & n90591;
  assign n90593 = P2_P1_EBX_REG_16_ & ~n90591;
  assign n90594 = ~n90592 & ~n90593;
  assign n90595 = n90441 & ~n90594;
  assign n90596 = ~n90589 & ~n90590;
  assign n16406 = n90595 | ~n90596;
  assign n90598 = P2_P1_EBX_REG_17_ & ~n90440;
  assign n90599 = ~n89762 & n90443;
  assign n90600 = P2_P1_EBX_REG_15_ & P2_P1_EBX_REG_16_;
  assign n90601 = n90582 & n90600;
  assign n90602 = P2_P1_EBX_REG_17_ & ~n90601;
  assign n90603 = ~P2_P1_EBX_REG_17_ & n90601;
  assign n90604 = ~n90602 & ~n90603;
  assign n90605 = n90441 & ~n90604;
  assign n90606 = ~n90598 & ~n90599;
  assign n16411 = n90605 | ~n90606;
  assign n90608 = P2_P1_EBX_REG_18_ & ~n90440;
  assign n90609 = ~n89806 & n90443;
  assign n90610 = P2_P1_EBX_REG_17_ & n90601;
  assign n90611 = ~P2_P1_EBX_REG_18_ & n90610;
  assign n90612 = P2_P1_EBX_REG_18_ & ~n90610;
  assign n90613 = ~n90611 & ~n90612;
  assign n90614 = n90441 & ~n90613;
  assign n90615 = ~n90608 & ~n90609;
  assign n16416 = n90614 | ~n90615;
  assign n90617 = P2_P1_EBX_REG_19_ & ~n90440;
  assign n90618 = ~n89850 & n90443;
  assign n90619 = P2_P1_EBX_REG_17_ & P2_P1_EBX_REG_18_;
  assign n90620 = n90601 & n90619;
  assign n90621 = P2_P1_EBX_REG_19_ & ~n90620;
  assign n90622 = ~P2_P1_EBX_REG_19_ & n90620;
  assign n90623 = ~n90621 & ~n90622;
  assign n90624 = n90441 & ~n90623;
  assign n90625 = ~n90617 & ~n90618;
  assign n16421 = n90624 | ~n90625;
  assign n90627 = P2_P1_EBX_REG_20_ & ~n90440;
  assign n90628 = ~n89894 & n90443;
  assign n90629 = P2_P1_EBX_REG_19_ & n90620;
  assign n90630 = ~P2_P1_EBX_REG_20_ & n90629;
  assign n90631 = P2_P1_EBX_REG_20_ & ~n90629;
  assign n90632 = ~n90630 & ~n90631;
  assign n90633 = n90441 & ~n90632;
  assign n90634 = ~n90627 & ~n90628;
  assign n16426 = n90633 | ~n90634;
  assign n90636 = P2_P1_EBX_REG_21_ & ~n90440;
  assign n90637 = ~n89938 & n90443;
  assign n90638 = P2_P1_EBX_REG_19_ & P2_P1_EBX_REG_20_;
  assign n90639 = n90620 & n90638;
  assign n90640 = P2_P1_EBX_REG_21_ & ~n90639;
  assign n90641 = ~P2_P1_EBX_REG_21_ & n90639;
  assign n90642 = ~n90640 & ~n90641;
  assign n90643 = n90441 & ~n90642;
  assign n90644 = ~n90636 & ~n90637;
  assign n16431 = n90643 | ~n90644;
  assign n90646 = P2_P1_EBX_REG_22_ & ~n90440;
  assign n90647 = ~n89982 & n90443;
  assign n90648 = P2_P1_EBX_REG_21_ & n90639;
  assign n90649 = ~P2_P1_EBX_REG_22_ & n90648;
  assign n90650 = P2_P1_EBX_REG_22_ & ~n90648;
  assign n90651 = ~n90649 & ~n90650;
  assign n90652 = n90441 & ~n90651;
  assign n90653 = ~n90646 & ~n90647;
  assign n16436 = n90652 | ~n90653;
  assign n90655 = P2_P1_EBX_REG_23_ & ~n90440;
  assign n90656 = ~n90080 & n90443;
  assign n90657 = P2_P1_EBX_REG_21_ & P2_P1_EBX_REG_22_;
  assign n90658 = n90639 & n90657;
  assign n90659 = P2_P1_EBX_REG_23_ & ~n90658;
  assign n90660 = ~P2_P1_EBX_REG_23_ & n90658;
  assign n90661 = ~n90659 & ~n90660;
  assign n90662 = n90441 & ~n90661;
  assign n90663 = ~n90655 & ~n90656;
  assign n16441 = n90662 | ~n90663;
  assign n90665 = P2_P1_EBX_REG_24_ & ~n90440;
  assign n90666 = ~n90128 & n90443;
  assign n90667 = P2_P1_EBX_REG_23_ & n90658;
  assign n90668 = ~P2_P1_EBX_REG_24_ & n90667;
  assign n90669 = P2_P1_EBX_REG_24_ & ~n90667;
  assign n90670 = ~n90668 & ~n90669;
  assign n90671 = n90441 & ~n90670;
  assign n90672 = ~n90665 & ~n90666;
  assign n16446 = n90671 | ~n90672;
  assign n90674 = P2_P1_EBX_REG_25_ & ~n90440;
  assign n90675 = ~n90176 & n90443;
  assign n90676 = P2_P1_EBX_REG_23_ & P2_P1_EBX_REG_24_;
  assign n90677 = n90658 & n90676;
  assign n90678 = P2_P1_EBX_REG_25_ & ~n90677;
  assign n90679 = ~P2_P1_EBX_REG_25_ & n90677;
  assign n90680 = ~n90678 & ~n90679;
  assign n90681 = n90441 & ~n90680;
  assign n90682 = ~n90674 & ~n90675;
  assign n16451 = n90681 | ~n90682;
  assign n90684 = P2_P1_EBX_REG_26_ & ~n90440;
  assign n90685 = ~n90224 & n90443;
  assign n90686 = P2_P1_EBX_REG_25_ & n90677;
  assign n90687 = ~P2_P1_EBX_REG_26_ & n90686;
  assign n90688 = P2_P1_EBX_REG_26_ & ~n90686;
  assign n90689 = ~n90687 & ~n90688;
  assign n90690 = n90441 & ~n90689;
  assign n90691 = ~n90684 & ~n90685;
  assign n16456 = n90690 | ~n90691;
  assign n90693 = P2_P1_EBX_REG_27_ & ~n90440;
  assign n90694 = ~n90272 & n90443;
  assign n90695 = P2_P1_EBX_REG_25_ & P2_P1_EBX_REG_26_;
  assign n90696 = n90677 & n90695;
  assign n90697 = P2_P1_EBX_REG_27_ & ~n90696;
  assign n90698 = ~P2_P1_EBX_REG_27_ & n90696;
  assign n90699 = ~n90697 & ~n90698;
  assign n90700 = n90441 & ~n90699;
  assign n90701 = ~n90693 & ~n90694;
  assign n16461 = n90700 | ~n90701;
  assign n90703 = P2_P1_EBX_REG_28_ & ~n90440;
  assign n90704 = ~n90326 & n90443;
  assign n90705 = P2_P1_EBX_REG_27_ & n90696;
  assign n90706 = ~P2_P1_EBX_REG_28_ & n90705;
  assign n90707 = P2_P1_EBX_REG_28_ & ~n90705;
  assign n90708 = ~n90706 & ~n90707;
  assign n90709 = n90441 & ~n90708;
  assign n90710 = ~n90703 & ~n90704;
  assign n16466 = n90709 | ~n90710;
  assign n90712 = P2_P1_EBX_REG_29_ & ~n90440;
  assign n90713 = ~n90374 & n90443;
  assign n90714 = P2_P1_EBX_REG_27_ & P2_P1_EBX_REG_28_;
  assign n90715 = n90696 & n90714;
  assign n90716 = P2_P1_EBX_REG_29_ & ~n90715;
  assign n90717 = ~P2_P1_EBX_REG_29_ & n90715;
  assign n90718 = ~n90716 & ~n90717;
  assign n90719 = n90441 & ~n90718;
  assign n90720 = ~n90712 & ~n90713;
  assign n16471 = n90719 | ~n90720;
  assign n90722 = P2_P1_EBX_REG_30_ & ~n90440;
  assign n90723 = ~n90422 & n90443;
  assign n90724 = P2_P1_EBX_REG_29_ & n90715;
  assign n90725 = ~P2_P1_EBX_REG_30_ & n90724;
  assign n90726 = P2_P1_EBX_REG_30_ & ~n90724;
  assign n90727 = ~n90725 & ~n90726;
  assign n90728 = n90441 & ~n90727;
  assign n90729 = ~n90722 & ~n90723;
  assign n16476 = n90728 | ~n90729;
  assign n90731 = P2_P1_EBX_REG_31_ & ~n90440;
  assign n90732 = P2_P1_EBX_REG_30_ & n90724;
  assign n90733 = ~P2_P1_EBX_REG_31_ & n90732;
  assign n90734 = P2_P1_EBX_REG_31_ & ~n90732;
  assign n90735 = ~n90733 & ~n90734;
  assign n90736 = n90441 & ~n90735;
  assign n16481 = n90731 | n90736;
  assign n90738 = ~n77322 & ~n77361;
  assign n90739 = ~n85231 & n90738;
  assign n90740 = n77189 & n77197;
  assign n90741 = n77311 & ~n90740;
  assign n90742 = n90739 & ~n90741;
  assign n90743 = P2_P1_STATE2_REG_2_ & ~n90742;
  assign n90744 = n77039 & n90743;
  assign n90745 = ~n76672 & n90744;
  assign n90746 = ~P2_P1_EBX_REG_31_ & n90745;
  assign n90747 = n76957 & n90743;
  assign n90748 = ~n76675 & n90747;
  assign n90749 = n76675 & n90747;
  assign n90750 = ~n76672 & n90749;
  assign n90751 = ~n90746 & ~n90748;
  assign n90752 = ~n90750 & n90751;
  assign n90753 = P2_P1_EBX_REG_0_ & ~n90752;
  assign n90754 = n76672 & n90749;
  assign n90755 = P2_P1_REIP_REG_0_ & n90754;
  assign n90756 = P2_P1_EBX_REG_31_ & n90745;
  assign n90757 = P2_P1_EBX_REG_0_ & n90756;
  assign n90758 = n77034 & n90743;
  assign n90759 = ~P2_P1_INSTQUEUERD_ADDR_REG_0_ & n90758;
  assign n90760 = n77030 & n90743;
  assign n90761 = ~P2_P1_INSTQUEUERD_ADDR_REG_0_ & n90760;
  assign n90762 = ~n90759 & ~n90761;
  assign n90763 = ~n90755 & ~n90757;
  assign n90764 = n90762 & n90763;
  assign n90765 = n76672 & n90744;
  assign n90766 = P2_P1_REIP_REG_0_ & n90765;
  assign n90767 = P2_P1_STATE2_REG_1_ & ~n90742;
  assign n90768 = n88812 & n90767;
  assign n90769 = P2_P1_PHYADDRPOINTER_REG_0_ & n90768;
  assign n90770 = P2_P1_REIP_REG_0_ & n90742;
  assign n90771 = P2_P1_STATE2_REG_3_ & ~n90742;
  assign n90772 = P2_P1_PHYADDRPOINTER_REG_0_ & n90771;
  assign n90773 = ~n90770 & ~n90772;
  assign n90774 = ~n88812 & n90767;
  assign n90775 = P2_P1_PHYADDRPOINTER_REG_0_ & n90774;
  assign n90776 = n90773 & ~n90775;
  assign n90777 = ~n90753 & n90764;
  assign n90778 = ~n90766 & n90777;
  assign n90779 = ~n90769 & n90778;
  assign n16486 = ~n90776 | ~n90779;
  assign n90781 = P2_P1_EBX_REG_1_ & ~n90752;
  assign n90782 = ~P2_P1_REIP_REG_1_ & n90754;
  assign n90783 = ~n90450 & n90756;
  assign n90784 = ~n76681 & ~n76686;
  assign n90785 = n90758 & ~n90784;
  assign n90786 = n90760 & ~n90784;
  assign n90787 = ~n90785 & ~n90786;
  assign n90788 = ~n90782 & ~n90783;
  assign n90789 = n90787 & n90788;
  assign n90790 = ~P2_P1_REIP_REG_1_ & n90765;
  assign n90791 = ~P2_P1_PHYADDRPOINTER_REG_1_ & n90768;
  assign n90792 = P2_P1_REIP_REG_1_ & n90742;
  assign n90793 = P2_P1_PHYADDRPOINTER_REG_1_ & n90771;
  assign n90794 = ~n90792 & ~n90793;
  assign n90795 = P2_P1_PHYADDRPOINTER_REG_0_ & P2_P1_PHYADDRPOINTER_REG_1_;
  assign n90796 = ~P2_P1_PHYADDRPOINTER_REG_0_ & ~P2_P1_PHYADDRPOINTER_REG_1_;
  assign n90797 = ~n90795 & ~n90796;
  assign n90798 = n90774 & ~n90797;
  assign n90799 = n90794 & ~n90798;
  assign n90800 = ~n90781 & n90789;
  assign n90801 = ~n90790 & n90800;
  assign n90802 = ~n90791 & n90801;
  assign n16491 = ~n90799 | ~n90802;
  assign n90804 = P2_P1_EBX_REG_2_ & ~n90752;
  assign n90805 = P2_P1_REIP_REG_1_ & ~P2_P1_REIP_REG_2_;
  assign n90806 = ~P2_P1_REIP_REG_1_ & P2_P1_REIP_REG_2_;
  assign n90807 = ~n90805 & ~n90806;
  assign n90808 = n90754 & ~n90807;
  assign n90809 = ~P2_P1_EBX_REG_0_ & ~P2_P1_EBX_REG_1_;
  assign n90810 = P2_P1_EBX_REG_2_ & ~n90809;
  assign n90811 = ~P2_P1_EBX_REG_2_ & n90809;
  assign n90812 = ~n90810 & ~n90811;
  assign n90813 = n90756 & n90812;
  assign n90814 = ~n77159 & n90758;
  assign n90815 = ~n77159 & n90760;
  assign n90816 = ~n90814 & ~n90815;
  assign n90817 = ~n90808 & ~n90813;
  assign n90818 = n90816 & n90817;
  assign n90819 = n90765 & ~n90807;
  assign n90820 = ~n88146 & n90768;
  assign n90821 = P2_P1_REIP_REG_2_ & n90742;
  assign n90822 = P2_P1_PHYADDRPOINTER_REG_2_ & n90771;
  assign n90823 = ~n90821 & ~n90822;
  assign n90824 = ~P2_P1_PHYADDRPOINTER_REG_0_ & P2_P1_PHYADDRPOINTER_REG_1_;
  assign n90825 = ~n88146 & ~n90824;
  assign n90826 = n88146 & n90824;
  assign n90827 = ~n90825 & ~n90826;
  assign n90828 = n90774 & n90827;
  assign n90829 = n90823 & ~n90828;
  assign n90830 = ~n90804 & n90818;
  assign n90831 = ~n90819 & n90830;
  assign n90832 = ~n90820 & n90831;
  assign n16496 = ~n90829 | ~n90832;
  assign n90834 = P2_P1_EBX_REG_3_ & ~n90752;
  assign n90835 = P2_P1_REIP_REG_1_ & P2_P1_REIP_REG_2_;
  assign n90836 = ~P2_P1_REIP_REG_3_ & n90835;
  assign n90837 = P2_P1_REIP_REG_3_ & ~n90835;
  assign n90838 = ~n90836 & ~n90837;
  assign n90839 = n90754 & ~n90838;
  assign n90840 = ~P2_P1_EBX_REG_3_ & n90811;
  assign n90841 = P2_P1_EBX_REG_3_ & ~n90811;
  assign n90842 = ~n90840 & ~n90841;
  assign n90843 = n90756 & n90842;
  assign n90844 = ~P2_P1_INSTQUEUERD_ADDR_REG_3_ & n77207;
  assign n90845 = ~n77208 & ~n90844;
  assign n90846 = n90758 & ~n90845;
  assign n90847 = n90760 & ~n90845;
  assign n90848 = ~n90846 & ~n90847;
  assign n90849 = ~n90839 & ~n90843;
  assign n90850 = n90848 & n90849;
  assign n90851 = n90765 & ~n90838;
  assign n90852 = ~n88168 & n90768;
  assign n90853 = P2_P1_REIP_REG_3_ & n90742;
  assign n90854 = P2_P1_PHYADDRPOINTER_REG_3_ & n90771;
  assign n90855 = ~n90853 & ~n90854;
  assign n90856 = n88168 & n90826;
  assign n90857 = ~n88168 & ~n90826;
  assign n90858 = ~n90856 & ~n90857;
  assign n90859 = n90774 & n90858;
  assign n90860 = n90855 & ~n90859;
  assign n90861 = ~n90834 & n90850;
  assign n90862 = ~n90851 & n90861;
  assign n90863 = ~n90852 & n90862;
  assign n16501 = ~n90860 | ~n90863;
  assign n90865 = P2_P1_INSTQUEUERD_ADDR_REG_3_ & n77207;
  assign n90866 = ~P2_P1_INSTQUEUERD_ADDR_REG_4_ & n90865;
  assign n90867 = P2_P1_INSTQUEUERD_ADDR_REG_4_ & ~n90865;
  assign n90868 = ~n90866 & ~n90867;
  assign n90869 = n90760 & ~n90868;
  assign n90870 = n90758 & ~n90868;
  assign n90871 = ~n90869 & ~n90870;
  assign n90872 = P2_P1_EBX_REG_4_ & ~n90752;
  assign n90873 = P2_P1_EBX_REG_4_ & ~n90840;
  assign n90874 = ~P2_P1_EBX_REG_3_ & ~P2_P1_EBX_REG_4_;
  assign n90875 = n90811 & n90874;
  assign n90876 = ~n90873 & ~n90875;
  assign n90877 = n90756 & n90876;
  assign n90878 = n85230 & ~n90742;
  assign n90879 = P2_P1_REIP_REG_3_ & n90835;
  assign n90880 = ~P2_P1_REIP_REG_4_ & n90879;
  assign n90881 = P2_P1_REIP_REG_4_ & ~n90879;
  assign n90882 = ~n90880 & ~n90881;
  assign n90883 = n90754 & ~n90882;
  assign n90884 = ~n90877 & ~n90878;
  assign n90885 = ~n90883 & n90884;
  assign n90886 = n90765 & ~n90882;
  assign n90887 = ~n88189 & n90768;
  assign n90888 = n90871 & ~n90872;
  assign n90889 = n90885 & n90888;
  assign n90890 = ~n90886 & n90889;
  assign n90891 = ~n90887 & n90890;
  assign n90892 = P2_P1_REIP_REG_4_ & n90742;
  assign n90893 = P2_P1_PHYADDRPOINTER_REG_4_ & n90771;
  assign n90894 = ~n90892 & ~n90893;
  assign n90895 = ~n88189 & ~n90856;
  assign n90896 = n88168 & n88189;
  assign n90897 = n90826 & n90896;
  assign n90898 = ~n90895 & ~n90897;
  assign n90899 = n90774 & n90898;
  assign n90900 = n90894 & ~n90899;
  assign n16506 = ~n90891 | ~n90900;
  assign n90902 = P2_P1_INSTQUEUERD_ADDR_REG_4_ & n90865;
  assign n90903 = n90760 & n90902;
  assign n90904 = n90758 & n90902;
  assign n90905 = ~n90903 & ~n90904;
  assign n90906 = P2_P1_EBX_REG_5_ & ~n90752;
  assign n90907 = ~P2_P1_EBX_REG_5_ & n90875;
  assign n90908 = P2_P1_EBX_REG_5_ & ~n90875;
  assign n90909 = ~n90907 & ~n90908;
  assign n90910 = n90756 & n90909;
  assign n90911 = P2_P1_REIP_REG_4_ & n90879;
  assign n90912 = ~P2_P1_REIP_REG_5_ & n90911;
  assign n90913 = P2_P1_REIP_REG_5_ & ~n90911;
  assign n90914 = ~n90912 & ~n90913;
  assign n90915 = n90754 & ~n90914;
  assign n90916 = ~n90878 & ~n90910;
  assign n90917 = ~n90915 & n90916;
  assign n90918 = n90765 & ~n90914;
  assign n90919 = ~n88212 & n90768;
  assign n90920 = n90905 & ~n90906;
  assign n90921 = n90917 & n90920;
  assign n90922 = ~n90918 & n90921;
  assign n90923 = ~n90919 & n90922;
  assign n90924 = P2_P1_REIP_REG_5_ & n90742;
  assign n90925 = P2_P1_PHYADDRPOINTER_REG_5_ & n90771;
  assign n90926 = ~n90924 & ~n90925;
  assign n90927 = n88212 & n90897;
  assign n90928 = ~n88212 & ~n90897;
  assign n90929 = ~n90927 & ~n90928;
  assign n90930 = n90774 & n90929;
  assign n90931 = n90926 & ~n90930;
  assign n16511 = ~n90923 | ~n90931;
  assign n90933 = P2_P1_REIP_REG_5_ & n90911;
  assign n90934 = ~P2_P1_REIP_REG_6_ & n90933;
  assign n90935 = P2_P1_REIP_REG_6_ & ~n90933;
  assign n90936 = ~n90934 & ~n90935;
  assign n90937 = n90765 & ~n90936;
  assign n90938 = P2_P1_EBX_REG_6_ & ~n90752;
  assign n90939 = P2_P1_EBX_REG_6_ & ~n90907;
  assign n90940 = ~P2_P1_EBX_REG_5_ & ~P2_P1_EBX_REG_6_;
  assign n90941 = n90875 & n90940;
  assign n90942 = ~n90939 & ~n90941;
  assign n90943 = n90756 & n90942;
  assign n90944 = n90754 & ~n90936;
  assign n90945 = ~n90878 & ~n90943;
  assign n90946 = ~n90944 & n90945;
  assign n90947 = ~n88235 & ~n90927;
  assign n90948 = n88212 & n88235;
  assign n90949 = n90897 & n90948;
  assign n90950 = ~n90947 & ~n90949;
  assign n90951 = n90774 & n90950;
  assign n90952 = P2_P1_REIP_REG_6_ & n90742;
  assign n90953 = P2_P1_PHYADDRPOINTER_REG_6_ & n90771;
  assign n90954 = ~n90952 & ~n90953;
  assign n90955 = ~n88235 & n90768;
  assign n90956 = n90954 & ~n90955;
  assign n90957 = ~n90937 & ~n90938;
  assign n90958 = n90946 & n90957;
  assign n90959 = ~n90951 & n90958;
  assign n16516 = ~n90956 | ~n90959;
  assign n90961 = P2_P1_REIP_REG_6_ & n90933;
  assign n90962 = ~P2_P1_REIP_REG_7_ & n90961;
  assign n90963 = P2_P1_REIP_REG_7_ & ~n90961;
  assign n90964 = ~n90962 & ~n90963;
  assign n90965 = n90765 & ~n90964;
  assign n90966 = P2_P1_EBX_REG_7_ & ~n90752;
  assign n90967 = ~P2_P1_EBX_REG_7_ & n90941;
  assign n90968 = P2_P1_EBX_REG_7_ & ~n90941;
  assign n90969 = ~n90967 & ~n90968;
  assign n90970 = n90756 & n90969;
  assign n90971 = n90754 & ~n90964;
  assign n90972 = ~n90878 & ~n90970;
  assign n90973 = ~n90971 & n90972;
  assign n90974 = n88258 & n90949;
  assign n90975 = ~n88258 & ~n90949;
  assign n90976 = ~n90974 & ~n90975;
  assign n90977 = n90774 & n90976;
  assign n90978 = P2_P1_REIP_REG_7_ & n90742;
  assign n90979 = P2_P1_PHYADDRPOINTER_REG_7_ & n90771;
  assign n90980 = ~n90978 & ~n90979;
  assign n90981 = ~n88258 & n90768;
  assign n90982 = n90980 & ~n90981;
  assign n90983 = ~n90965 & ~n90966;
  assign n90984 = n90973 & n90983;
  assign n90985 = ~n90977 & n90984;
  assign n16521 = ~n90982 | ~n90985;
  assign n90987 = P2_P1_REIP_REG_7_ & n90961;
  assign n90988 = ~P2_P1_REIP_REG_8_ & n90987;
  assign n90989 = P2_P1_REIP_REG_8_ & ~n90987;
  assign n90990 = ~n90988 & ~n90989;
  assign n90991 = n90765 & ~n90990;
  assign n90992 = P2_P1_EBX_REG_8_ & ~n90752;
  assign n90993 = P2_P1_EBX_REG_8_ & ~n90967;
  assign n90994 = ~P2_P1_EBX_REG_7_ & ~P2_P1_EBX_REG_8_;
  assign n90995 = n90941 & n90994;
  assign n90996 = ~n90993 & ~n90995;
  assign n90997 = n90756 & n90996;
  assign n90998 = n90754 & ~n90990;
  assign n90999 = ~n90878 & ~n90997;
  assign n91000 = ~n90998 & n90999;
  assign n91001 = ~n88281 & ~n90974;
  assign n91002 = n88258 & n88281;
  assign n91003 = n90949 & n91002;
  assign n91004 = ~n91001 & ~n91003;
  assign n91005 = n90774 & n91004;
  assign n91006 = P2_P1_REIP_REG_8_ & n90742;
  assign n91007 = P2_P1_PHYADDRPOINTER_REG_8_ & n90771;
  assign n91008 = ~n91006 & ~n91007;
  assign n91009 = ~n88281 & n90768;
  assign n91010 = n91008 & ~n91009;
  assign n91011 = ~n90991 & ~n90992;
  assign n91012 = n91000 & n91011;
  assign n91013 = ~n91005 & n91012;
  assign n16526 = ~n91010 | ~n91013;
  assign n91015 = P2_P1_REIP_REG_8_ & n90987;
  assign n91016 = ~P2_P1_REIP_REG_9_ & n91015;
  assign n91017 = P2_P1_REIP_REG_9_ & ~n91015;
  assign n91018 = ~n91016 & ~n91017;
  assign n91019 = n90765 & ~n91018;
  assign n91020 = P2_P1_EBX_REG_9_ & ~n90752;
  assign n91021 = ~P2_P1_EBX_REG_9_ & n90995;
  assign n91022 = P2_P1_EBX_REG_9_ & ~n90995;
  assign n91023 = ~n91021 & ~n91022;
  assign n91024 = n90756 & n91023;
  assign n91025 = n90754 & ~n91018;
  assign n91026 = ~n90878 & ~n91024;
  assign n91027 = ~n91025 & n91026;
  assign n91028 = n88304 & n91003;
  assign n91029 = ~n88304 & ~n91003;
  assign n91030 = ~n91028 & ~n91029;
  assign n91031 = n90774 & n91030;
  assign n91032 = P2_P1_REIP_REG_9_ & n90742;
  assign n91033 = P2_P1_PHYADDRPOINTER_REG_9_ & n90771;
  assign n91034 = ~n91032 & ~n91033;
  assign n91035 = ~n88304 & n90768;
  assign n91036 = n91034 & ~n91035;
  assign n91037 = ~n91019 & ~n91020;
  assign n91038 = n91027 & n91037;
  assign n91039 = ~n91031 & n91038;
  assign n16531 = ~n91036 | ~n91039;
  assign n91041 = P2_P1_REIP_REG_9_ & n91015;
  assign n91042 = ~P2_P1_REIP_REG_10_ & n91041;
  assign n91043 = P2_P1_REIP_REG_10_ & ~n91041;
  assign n91044 = ~n91042 & ~n91043;
  assign n91045 = n90765 & ~n91044;
  assign n91046 = P2_P1_EBX_REG_10_ & ~n90752;
  assign n91047 = P2_P1_EBX_REG_10_ & ~n91021;
  assign n91048 = ~P2_P1_EBX_REG_9_ & ~P2_P1_EBX_REG_10_;
  assign n91049 = n90995 & n91048;
  assign n91050 = ~n91047 & ~n91049;
  assign n91051 = n90756 & n91050;
  assign n91052 = n90754 & ~n91044;
  assign n91053 = ~n90878 & ~n91051;
  assign n91054 = ~n91052 & n91053;
  assign n91055 = ~n88327 & ~n91028;
  assign n91056 = n88304 & n88327;
  assign n91057 = n91003 & n91056;
  assign n91058 = ~n91055 & ~n91057;
  assign n91059 = n90774 & n91058;
  assign n91060 = P2_P1_REIP_REG_10_ & n90742;
  assign n91061 = P2_P1_PHYADDRPOINTER_REG_10_ & n90771;
  assign n91062 = ~n91060 & ~n91061;
  assign n91063 = ~n88327 & n90768;
  assign n91064 = n91062 & ~n91063;
  assign n91065 = ~n91045 & ~n91046;
  assign n91066 = n91054 & n91065;
  assign n91067 = ~n91059 & n91066;
  assign n16536 = ~n91064 | ~n91067;
  assign n91069 = P2_P1_REIP_REG_10_ & n91041;
  assign n91070 = ~P2_P1_REIP_REG_11_ & n91069;
  assign n91071 = P2_P1_REIP_REG_11_ & ~n91069;
  assign n91072 = ~n91070 & ~n91071;
  assign n91073 = n90765 & ~n91072;
  assign n91074 = P2_P1_EBX_REG_11_ & ~n90752;
  assign n91075 = ~P2_P1_EBX_REG_11_ & n91049;
  assign n91076 = P2_P1_EBX_REG_11_ & ~n91049;
  assign n91077 = ~n91075 & ~n91076;
  assign n91078 = n90756 & n91077;
  assign n91079 = n90754 & ~n91072;
  assign n91080 = ~n90878 & ~n91078;
  assign n91081 = ~n91079 & n91080;
  assign n91082 = n88350 & n91057;
  assign n91083 = ~n88350 & ~n91057;
  assign n91084 = ~n91082 & ~n91083;
  assign n91085 = n90774 & n91084;
  assign n91086 = P2_P1_REIP_REG_11_ & n90742;
  assign n91087 = P2_P1_PHYADDRPOINTER_REG_11_ & n90771;
  assign n91088 = ~n91086 & ~n91087;
  assign n91089 = ~n88350 & n90768;
  assign n91090 = n91088 & ~n91089;
  assign n91091 = ~n91073 & ~n91074;
  assign n91092 = n91081 & n91091;
  assign n91093 = ~n91085 & n91092;
  assign n16541 = ~n91090 | ~n91093;
  assign n91095 = P2_P1_REIP_REG_11_ & n91069;
  assign n91096 = ~P2_P1_REIP_REG_12_ & n91095;
  assign n91097 = P2_P1_REIP_REG_12_ & ~n91095;
  assign n91098 = ~n91096 & ~n91097;
  assign n91099 = n90765 & ~n91098;
  assign n91100 = P2_P1_EBX_REG_12_ & ~n90752;
  assign n91101 = P2_P1_EBX_REG_12_ & ~n91075;
  assign n91102 = ~P2_P1_EBX_REG_11_ & ~P2_P1_EBX_REG_12_;
  assign n91103 = n91049 & n91102;
  assign n91104 = ~n91101 & ~n91103;
  assign n91105 = n90756 & n91104;
  assign n91106 = n90754 & ~n91098;
  assign n91107 = ~n90878 & ~n91105;
  assign n91108 = ~n91106 & n91107;
  assign n91109 = ~n88373 & ~n91082;
  assign n91110 = n88350 & n88373;
  assign n91111 = n91057 & n91110;
  assign n91112 = ~n91109 & ~n91111;
  assign n91113 = n90774 & n91112;
  assign n91114 = P2_P1_REIP_REG_12_ & n90742;
  assign n91115 = P2_P1_PHYADDRPOINTER_REG_12_ & n90771;
  assign n91116 = ~n91114 & ~n91115;
  assign n91117 = ~n88373 & n90768;
  assign n91118 = n91116 & ~n91117;
  assign n91119 = ~n91099 & ~n91100;
  assign n91120 = n91108 & n91119;
  assign n91121 = ~n91113 & n91120;
  assign n16546 = ~n91118 | ~n91121;
  assign n91123 = P2_P1_REIP_REG_12_ & n91095;
  assign n91124 = ~P2_P1_REIP_REG_13_ & n91123;
  assign n91125 = P2_P1_REIP_REG_13_ & ~n91123;
  assign n91126 = ~n91124 & ~n91125;
  assign n91127 = n90765 & ~n91126;
  assign n91128 = P2_P1_EBX_REG_13_ & ~n90752;
  assign n91129 = ~P2_P1_EBX_REG_13_ & n91103;
  assign n91130 = P2_P1_EBX_REG_13_ & ~n91103;
  assign n91131 = ~n91129 & ~n91130;
  assign n91132 = n90756 & n91131;
  assign n91133 = n90754 & ~n91126;
  assign n91134 = ~n90878 & ~n91132;
  assign n91135 = ~n91133 & n91134;
  assign n91136 = n88396 & n91111;
  assign n91137 = ~n88396 & ~n91111;
  assign n91138 = ~n91136 & ~n91137;
  assign n91139 = n90774 & n91138;
  assign n91140 = P2_P1_REIP_REG_13_ & n90742;
  assign n91141 = P2_P1_PHYADDRPOINTER_REG_13_ & n90771;
  assign n91142 = ~n91140 & ~n91141;
  assign n91143 = ~n88396 & n90768;
  assign n91144 = n91142 & ~n91143;
  assign n91145 = ~n91127 & ~n91128;
  assign n91146 = n91135 & n91145;
  assign n91147 = ~n91139 & n91146;
  assign n16551 = ~n91144 | ~n91147;
  assign n91149 = P2_P1_REIP_REG_13_ & n91123;
  assign n91150 = ~P2_P1_REIP_REG_14_ & n91149;
  assign n91151 = P2_P1_REIP_REG_14_ & ~n91149;
  assign n91152 = ~n91150 & ~n91151;
  assign n91153 = n90765 & ~n91152;
  assign n91154 = P2_P1_EBX_REG_14_ & ~n90752;
  assign n91155 = P2_P1_EBX_REG_14_ & ~n91129;
  assign n91156 = ~P2_P1_EBX_REG_13_ & ~P2_P1_EBX_REG_14_;
  assign n91157 = n91103 & n91156;
  assign n91158 = ~n91155 & ~n91157;
  assign n91159 = n90756 & n91158;
  assign n91160 = n90754 & ~n91152;
  assign n91161 = ~n90878 & ~n91159;
  assign n91162 = ~n91160 & n91161;
  assign n91163 = ~n88419 & ~n91136;
  assign n91164 = n88396 & n88419;
  assign n91165 = n91111 & n91164;
  assign n91166 = ~n91163 & ~n91165;
  assign n91167 = n90774 & n91166;
  assign n91168 = P2_P1_REIP_REG_14_ & n90742;
  assign n91169 = P2_P1_PHYADDRPOINTER_REG_14_ & n90771;
  assign n91170 = ~n91168 & ~n91169;
  assign n91171 = ~n88419 & n90768;
  assign n91172 = n91170 & ~n91171;
  assign n91173 = ~n91153 & ~n91154;
  assign n91174 = n91162 & n91173;
  assign n91175 = ~n91167 & n91174;
  assign n16556 = ~n91172 | ~n91175;
  assign n91177 = P2_P1_REIP_REG_14_ & n91149;
  assign n91178 = ~P2_P1_REIP_REG_15_ & n91177;
  assign n91179 = P2_P1_REIP_REG_15_ & ~n91177;
  assign n91180 = ~n91178 & ~n91179;
  assign n91181 = n90765 & ~n91180;
  assign n91182 = P2_P1_EBX_REG_15_ & ~n90752;
  assign n91183 = ~P2_P1_EBX_REG_15_ & n91157;
  assign n91184 = P2_P1_EBX_REG_15_ & ~n91157;
  assign n91185 = ~n91183 & ~n91184;
  assign n91186 = n90756 & n91185;
  assign n91187 = n90754 & ~n91180;
  assign n91188 = ~n90878 & ~n91186;
  assign n91189 = ~n91187 & n91188;
  assign n91190 = n88442 & n91165;
  assign n91191 = ~n88442 & ~n91165;
  assign n91192 = ~n91190 & ~n91191;
  assign n91193 = n90774 & n91192;
  assign n91194 = P2_P1_REIP_REG_15_ & n90742;
  assign n91195 = P2_P1_PHYADDRPOINTER_REG_15_ & n90771;
  assign n91196 = ~n91194 & ~n91195;
  assign n91197 = ~n88442 & n90768;
  assign n91198 = n91196 & ~n91197;
  assign n91199 = ~n91181 & ~n91182;
  assign n91200 = n91189 & n91199;
  assign n91201 = ~n91193 & n91200;
  assign n16561 = ~n91198 | ~n91201;
  assign n91203 = P2_P1_REIP_REG_15_ & n91177;
  assign n91204 = ~P2_P1_REIP_REG_16_ & n91203;
  assign n91205 = P2_P1_REIP_REG_16_ & ~n91203;
  assign n91206 = ~n91204 & ~n91205;
  assign n91207 = n90765 & ~n91206;
  assign n91208 = P2_P1_EBX_REG_16_ & ~n90752;
  assign n91209 = P2_P1_EBX_REG_16_ & ~n91183;
  assign n91210 = ~P2_P1_EBX_REG_15_ & ~P2_P1_EBX_REG_16_;
  assign n91211 = n91157 & n91210;
  assign n91212 = ~n91209 & ~n91211;
  assign n91213 = n90756 & n91212;
  assign n91214 = n90754 & ~n91206;
  assign n91215 = ~n90878 & ~n91213;
  assign n91216 = ~n91214 & n91215;
  assign n91217 = ~n88465 & ~n91190;
  assign n91218 = n88442 & n88465;
  assign n91219 = n91165 & n91218;
  assign n91220 = ~n91217 & ~n91219;
  assign n91221 = n90774 & n91220;
  assign n91222 = P2_P1_REIP_REG_16_ & n90742;
  assign n91223 = P2_P1_PHYADDRPOINTER_REG_16_ & n90771;
  assign n91224 = ~n91222 & ~n91223;
  assign n91225 = ~n88465 & n90768;
  assign n91226 = n91224 & ~n91225;
  assign n91227 = ~n91207 & ~n91208;
  assign n91228 = n91216 & n91227;
  assign n91229 = ~n91221 & n91228;
  assign n16566 = ~n91226 | ~n91229;
  assign n91231 = P2_P1_REIP_REG_16_ & n91203;
  assign n91232 = ~P2_P1_REIP_REG_17_ & n91231;
  assign n91233 = P2_P1_REIP_REG_17_ & ~n91231;
  assign n91234 = ~n91232 & ~n91233;
  assign n91235 = n90765 & ~n91234;
  assign n91236 = P2_P1_EBX_REG_17_ & ~n90752;
  assign n91237 = ~P2_P1_EBX_REG_17_ & n91211;
  assign n91238 = P2_P1_EBX_REG_17_ & ~n91211;
  assign n91239 = ~n91237 & ~n91238;
  assign n91240 = n90756 & n91239;
  assign n91241 = n90754 & ~n91234;
  assign n91242 = ~n90878 & ~n91240;
  assign n91243 = ~n91241 & n91242;
  assign n91244 = n88488 & n91219;
  assign n91245 = ~n88488 & ~n91219;
  assign n91246 = ~n91244 & ~n91245;
  assign n91247 = n90774 & n91246;
  assign n91248 = P2_P1_REIP_REG_17_ & n90742;
  assign n91249 = P2_P1_PHYADDRPOINTER_REG_17_ & n90771;
  assign n91250 = ~n91248 & ~n91249;
  assign n91251 = ~n88488 & n90768;
  assign n91252 = n91250 & ~n91251;
  assign n91253 = ~n91235 & ~n91236;
  assign n91254 = n91243 & n91253;
  assign n91255 = ~n91247 & n91254;
  assign n16571 = ~n91252 | ~n91255;
  assign n91257 = P2_P1_REIP_REG_17_ & n91231;
  assign n91258 = ~P2_P1_REIP_REG_18_ & n91257;
  assign n91259 = P2_P1_REIP_REG_18_ & ~n91257;
  assign n91260 = ~n91258 & ~n91259;
  assign n91261 = n90765 & ~n91260;
  assign n91262 = P2_P1_EBX_REG_18_ & ~n90752;
  assign n91263 = P2_P1_EBX_REG_18_ & ~n91237;
  assign n91264 = ~P2_P1_EBX_REG_17_ & ~P2_P1_EBX_REG_18_;
  assign n91265 = n91211 & n91264;
  assign n91266 = ~n91263 & ~n91265;
  assign n91267 = n90756 & n91266;
  assign n91268 = n90754 & ~n91260;
  assign n91269 = ~n90878 & ~n91267;
  assign n91270 = ~n91268 & n91269;
  assign n91271 = ~n88511 & ~n91244;
  assign n91272 = n88488 & n88511;
  assign n91273 = n91219 & n91272;
  assign n91274 = ~n91271 & ~n91273;
  assign n91275 = n90774 & n91274;
  assign n91276 = P2_P1_REIP_REG_18_ & n90742;
  assign n91277 = P2_P1_PHYADDRPOINTER_REG_18_ & n90771;
  assign n91278 = ~n91276 & ~n91277;
  assign n91279 = ~n88511 & n90768;
  assign n91280 = n91278 & ~n91279;
  assign n91281 = ~n91261 & ~n91262;
  assign n91282 = n91270 & n91281;
  assign n91283 = ~n91275 & n91282;
  assign n16576 = ~n91280 | ~n91283;
  assign n91285 = P2_P1_REIP_REG_18_ & n91257;
  assign n91286 = ~P2_P1_REIP_REG_19_ & n91285;
  assign n91287 = P2_P1_REIP_REG_19_ & ~n91285;
  assign n91288 = ~n91286 & ~n91287;
  assign n91289 = n90765 & ~n91288;
  assign n91290 = P2_P1_EBX_REG_19_ & ~n90752;
  assign n91291 = ~P2_P1_EBX_REG_19_ & n91265;
  assign n91292 = P2_P1_EBX_REG_19_ & ~n91265;
  assign n91293 = ~n91291 & ~n91292;
  assign n91294 = n90756 & n91293;
  assign n91295 = n90754 & ~n91288;
  assign n91296 = ~n90878 & ~n91294;
  assign n91297 = ~n91295 & n91296;
  assign n91298 = n88534 & n91273;
  assign n91299 = ~n88534 & ~n91273;
  assign n91300 = ~n91298 & ~n91299;
  assign n91301 = n90774 & n91300;
  assign n91302 = P2_P1_REIP_REG_19_ & n90742;
  assign n91303 = P2_P1_PHYADDRPOINTER_REG_19_ & n90771;
  assign n91304 = ~n91302 & ~n91303;
  assign n91305 = ~n88534 & n90768;
  assign n91306 = n91304 & ~n91305;
  assign n91307 = ~n91289 & ~n91290;
  assign n91308 = n91297 & n91307;
  assign n91309 = ~n91301 & n91308;
  assign n16581 = ~n91306 | ~n91309;
  assign n91311 = P2_P1_REIP_REG_19_ & n91285;
  assign n91312 = ~P2_P1_REIP_REG_20_ & n91311;
  assign n91313 = P2_P1_REIP_REG_20_ & ~n91311;
  assign n91314 = ~n91312 & ~n91313;
  assign n91315 = n90765 & ~n91314;
  assign n91316 = P2_P1_EBX_REG_20_ & ~n90752;
  assign n91317 = n90754 & ~n91314;
  assign n91318 = P2_P1_EBX_REG_20_ & ~n91291;
  assign n91319 = ~P2_P1_EBX_REG_19_ & ~P2_P1_EBX_REG_20_;
  assign n91320 = n91265 & n91319;
  assign n91321 = ~n91318 & ~n91320;
  assign n91322 = n90756 & n91321;
  assign n91323 = ~n91317 & ~n91322;
  assign n91324 = ~n88557 & ~n91298;
  assign n91325 = n88534 & n88557;
  assign n91326 = n91273 & n91325;
  assign n91327 = ~n91324 & ~n91326;
  assign n91328 = n90774 & n91327;
  assign n91329 = P2_P1_REIP_REG_20_ & n90742;
  assign n91330 = P2_P1_PHYADDRPOINTER_REG_20_ & n90771;
  assign n91331 = ~n91329 & ~n91330;
  assign n91332 = ~n88557 & n90768;
  assign n91333 = n91331 & ~n91332;
  assign n91334 = ~n91315 & ~n91316;
  assign n91335 = n91323 & n91334;
  assign n91336 = ~n91328 & n91335;
  assign n16586 = ~n91333 | ~n91336;
  assign n91338 = P2_P1_REIP_REG_20_ & n91311;
  assign n91339 = ~P2_P1_REIP_REG_21_ & n91338;
  assign n91340 = P2_P1_REIP_REG_21_ & ~n91338;
  assign n91341 = ~n91339 & ~n91340;
  assign n91342 = n90765 & ~n91341;
  assign n91343 = P2_P1_EBX_REG_21_ & ~n90752;
  assign n91344 = n90754 & ~n91341;
  assign n91345 = ~P2_P1_EBX_REG_21_ & n91320;
  assign n91346 = P2_P1_EBX_REG_21_ & ~n91320;
  assign n91347 = ~n91345 & ~n91346;
  assign n91348 = n90756 & n91347;
  assign n91349 = ~n91344 & ~n91348;
  assign n91350 = n88580 & n91326;
  assign n91351 = ~n88580 & ~n91326;
  assign n91352 = ~n91350 & ~n91351;
  assign n91353 = n90774 & n91352;
  assign n91354 = P2_P1_REIP_REG_21_ & n90742;
  assign n91355 = P2_P1_PHYADDRPOINTER_REG_21_ & n90771;
  assign n91356 = ~n91354 & ~n91355;
  assign n91357 = ~n88580 & n90768;
  assign n91358 = n91356 & ~n91357;
  assign n91359 = ~n91342 & ~n91343;
  assign n91360 = n91349 & n91359;
  assign n91361 = ~n91353 & n91360;
  assign n16591 = ~n91358 | ~n91361;
  assign n91363 = P2_P1_REIP_REG_21_ & n91338;
  assign n91364 = ~P2_P1_REIP_REG_22_ & n91363;
  assign n91365 = P2_P1_REIP_REG_22_ & ~n91363;
  assign n91366 = ~n91364 & ~n91365;
  assign n91367 = n90765 & ~n91366;
  assign n91368 = P2_P1_EBX_REG_22_ & ~n90752;
  assign n91369 = n90754 & ~n91366;
  assign n91370 = P2_P1_EBX_REG_22_ & ~n91345;
  assign n91371 = ~P2_P1_EBX_REG_21_ & ~P2_P1_EBX_REG_22_;
  assign n91372 = n91320 & n91371;
  assign n91373 = ~n91370 & ~n91372;
  assign n91374 = n90756 & n91373;
  assign n91375 = ~n91369 & ~n91374;
  assign n91376 = ~n88604 & ~n91350;
  assign n91377 = n88580 & n88604;
  assign n91378 = n91326 & n91377;
  assign n91379 = ~n91376 & ~n91378;
  assign n91380 = n90774 & n91379;
  assign n91381 = P2_P1_REIP_REG_22_ & n90742;
  assign n91382 = P2_P1_PHYADDRPOINTER_REG_22_ & n90771;
  assign n91383 = ~n91381 & ~n91382;
  assign n91384 = ~n88604 & n90768;
  assign n91385 = n91383 & ~n91384;
  assign n91386 = ~n91367 & ~n91368;
  assign n91387 = n91375 & n91386;
  assign n91388 = ~n91380 & n91387;
  assign n16596 = ~n91385 | ~n91388;
  assign n91390 = P2_P1_REIP_REG_22_ & n91363;
  assign n91391 = ~P2_P1_REIP_REG_23_ & n91390;
  assign n91392 = P2_P1_REIP_REG_23_ & ~n91390;
  assign n91393 = ~n91391 & ~n91392;
  assign n91394 = n90765 & ~n91393;
  assign n91395 = P2_P1_EBX_REG_23_ & ~n90752;
  assign n91396 = n90754 & ~n91393;
  assign n91397 = ~P2_P1_EBX_REG_23_ & n91372;
  assign n91398 = P2_P1_EBX_REG_23_ & ~n91372;
  assign n91399 = ~n91397 & ~n91398;
  assign n91400 = n90756 & n91399;
  assign n91401 = ~n91396 & ~n91400;
  assign n91402 = n88627 & n91378;
  assign n91403 = ~n88627 & ~n91378;
  assign n91404 = ~n91402 & ~n91403;
  assign n91405 = n90774 & n91404;
  assign n91406 = P2_P1_REIP_REG_23_ & n90742;
  assign n91407 = P2_P1_PHYADDRPOINTER_REG_23_ & n90771;
  assign n91408 = ~n91406 & ~n91407;
  assign n91409 = ~n88627 & n90768;
  assign n91410 = n91408 & ~n91409;
  assign n91411 = ~n91394 & ~n91395;
  assign n91412 = n91401 & n91411;
  assign n91413 = ~n91405 & n91412;
  assign n16601 = ~n91410 | ~n91413;
  assign n91415 = P2_P1_REIP_REG_23_ & n91390;
  assign n91416 = ~P2_P1_REIP_REG_24_ & n91415;
  assign n91417 = P2_P1_REIP_REG_24_ & ~n91415;
  assign n91418 = ~n91416 & ~n91417;
  assign n91419 = n90765 & ~n91418;
  assign n91420 = P2_P1_EBX_REG_24_ & ~n90752;
  assign n91421 = n90754 & ~n91418;
  assign n91422 = P2_P1_EBX_REG_24_ & ~n91397;
  assign n91423 = ~P2_P1_EBX_REG_23_ & ~P2_P1_EBX_REG_24_;
  assign n91424 = n91372 & n91423;
  assign n91425 = ~n91422 & ~n91424;
  assign n91426 = n90756 & n91425;
  assign n91427 = ~n91421 & ~n91426;
  assign n91428 = ~n88650 & ~n91402;
  assign n91429 = n88627 & n88650;
  assign n91430 = n91378 & n91429;
  assign n91431 = ~n91428 & ~n91430;
  assign n91432 = n90774 & n91431;
  assign n91433 = P2_P1_REIP_REG_24_ & n90742;
  assign n91434 = P2_P1_PHYADDRPOINTER_REG_24_ & n90771;
  assign n91435 = ~n91433 & ~n91434;
  assign n91436 = ~n88650 & n90768;
  assign n91437 = n91435 & ~n91436;
  assign n91438 = ~n91419 & ~n91420;
  assign n91439 = n91427 & n91438;
  assign n91440 = ~n91432 & n91439;
  assign n16606 = ~n91437 | ~n91440;
  assign n91442 = P2_P1_REIP_REG_24_ & n91415;
  assign n91443 = ~P2_P1_REIP_REG_25_ & n91442;
  assign n91444 = P2_P1_REIP_REG_25_ & ~n91442;
  assign n91445 = ~n91443 & ~n91444;
  assign n91446 = n90765 & ~n91445;
  assign n91447 = P2_P1_EBX_REG_25_ & ~n90752;
  assign n91448 = n90754 & ~n91445;
  assign n91449 = ~P2_P1_EBX_REG_25_ & n91424;
  assign n91450 = P2_P1_EBX_REG_25_ & ~n91424;
  assign n91451 = ~n91449 & ~n91450;
  assign n91452 = n90756 & n91451;
  assign n91453 = ~n91448 & ~n91452;
  assign n91454 = n88673 & n91430;
  assign n91455 = ~n88673 & ~n91430;
  assign n91456 = ~n91454 & ~n91455;
  assign n91457 = n90774 & n91456;
  assign n91458 = P2_P1_REIP_REG_25_ & n90742;
  assign n91459 = P2_P1_PHYADDRPOINTER_REG_25_ & n90771;
  assign n91460 = ~n91458 & ~n91459;
  assign n91461 = ~n88673 & n90768;
  assign n91462 = n91460 & ~n91461;
  assign n91463 = ~n91446 & ~n91447;
  assign n91464 = n91453 & n91463;
  assign n91465 = ~n91457 & n91464;
  assign n16611 = ~n91462 | ~n91465;
  assign n91467 = P2_P1_REIP_REG_25_ & n91442;
  assign n91468 = ~P2_P1_REIP_REG_26_ & n91467;
  assign n91469 = P2_P1_REIP_REG_26_ & ~n91467;
  assign n91470 = ~n91468 & ~n91469;
  assign n91471 = n90765 & ~n91470;
  assign n91472 = P2_P1_EBX_REG_26_ & ~n90752;
  assign n91473 = n90754 & ~n91470;
  assign n91474 = P2_P1_EBX_REG_26_ & ~n91449;
  assign n91475 = ~P2_P1_EBX_REG_25_ & ~P2_P1_EBX_REG_26_;
  assign n91476 = n91424 & n91475;
  assign n91477 = ~n91474 & ~n91476;
  assign n91478 = n90756 & n91477;
  assign n91479 = ~n91473 & ~n91478;
  assign n91480 = ~n88696 & ~n91454;
  assign n91481 = n88673 & n88696;
  assign n91482 = n91430 & n91481;
  assign n91483 = ~n91480 & ~n91482;
  assign n91484 = n90774 & n91483;
  assign n91485 = P2_P1_REIP_REG_26_ & n90742;
  assign n91486 = P2_P1_PHYADDRPOINTER_REG_26_ & n90771;
  assign n91487 = ~n91485 & ~n91486;
  assign n91488 = ~n88696 & n90768;
  assign n91489 = n91487 & ~n91488;
  assign n91490 = ~n91471 & ~n91472;
  assign n91491 = n91479 & n91490;
  assign n91492 = ~n91484 & n91491;
  assign n16616 = ~n91489 | ~n91492;
  assign n91494 = P2_P1_REIP_REG_26_ & n91467;
  assign n91495 = ~P2_P1_REIP_REG_27_ & n91494;
  assign n91496 = P2_P1_REIP_REG_27_ & ~n91494;
  assign n91497 = ~n91495 & ~n91496;
  assign n91498 = n90765 & ~n91497;
  assign n91499 = P2_P1_EBX_REG_27_ & ~n90752;
  assign n91500 = n90754 & ~n91497;
  assign n91501 = ~P2_P1_EBX_REG_27_ & n91476;
  assign n91502 = P2_P1_EBX_REG_27_ & ~n91476;
  assign n91503 = ~n91501 & ~n91502;
  assign n91504 = n90756 & n91503;
  assign n91505 = ~n91500 & ~n91504;
  assign n91506 = n88719 & n91482;
  assign n91507 = ~n88719 & ~n91482;
  assign n91508 = ~n91506 & ~n91507;
  assign n91509 = n90774 & n91508;
  assign n91510 = P2_P1_REIP_REG_27_ & n90742;
  assign n91511 = P2_P1_PHYADDRPOINTER_REG_27_ & n90771;
  assign n91512 = ~n91510 & ~n91511;
  assign n91513 = ~n88719 & n90768;
  assign n91514 = n91512 & ~n91513;
  assign n91515 = ~n91498 & ~n91499;
  assign n91516 = n91505 & n91515;
  assign n91517 = ~n91509 & n91516;
  assign n16621 = ~n91514 | ~n91517;
  assign n91519 = P2_P1_REIP_REG_27_ & n91494;
  assign n91520 = ~P2_P1_REIP_REG_28_ & n91519;
  assign n91521 = P2_P1_REIP_REG_28_ & ~n91519;
  assign n91522 = ~n91520 & ~n91521;
  assign n91523 = n90765 & ~n91522;
  assign n91524 = P2_P1_EBX_REG_28_ & ~n90752;
  assign n91525 = n90754 & ~n91522;
  assign n91526 = P2_P1_EBX_REG_28_ & ~n91501;
  assign n91527 = ~P2_P1_EBX_REG_27_ & ~P2_P1_EBX_REG_28_;
  assign n91528 = n91476 & n91527;
  assign n91529 = ~n91526 & ~n91528;
  assign n91530 = n90756 & n91529;
  assign n91531 = ~n91525 & ~n91530;
  assign n91532 = ~n88743 & ~n91506;
  assign n91533 = n88719 & n88743;
  assign n91534 = n91482 & n91533;
  assign n91535 = ~n91532 & ~n91534;
  assign n91536 = n90774 & n91535;
  assign n91537 = P2_P1_REIP_REG_28_ & n90742;
  assign n91538 = P2_P1_PHYADDRPOINTER_REG_28_ & n90771;
  assign n91539 = ~n91537 & ~n91538;
  assign n91540 = ~n88743 & n90768;
  assign n91541 = n91539 & ~n91540;
  assign n91542 = ~n91523 & ~n91524;
  assign n91543 = n91531 & n91542;
  assign n91544 = ~n91536 & n91543;
  assign n16626 = ~n91541 | ~n91544;
  assign n91546 = P2_P1_REIP_REG_28_ & n91519;
  assign n91547 = ~P2_P1_REIP_REG_29_ & n91546;
  assign n91548 = P2_P1_REIP_REG_29_ & ~n91546;
  assign n91549 = ~n91547 & ~n91548;
  assign n91550 = n90765 & ~n91549;
  assign n91551 = P2_P1_EBX_REG_29_ & ~n90752;
  assign n91552 = n90754 & ~n91549;
  assign n91553 = P2_P1_EBX_REG_29_ & ~n91528;
  assign n91554 = ~P2_P1_EBX_REG_29_ & n91528;
  assign n91555 = ~n91553 & ~n91554;
  assign n91556 = n90756 & n91555;
  assign n91557 = ~n91552 & ~n91556;
  assign n91558 = ~n88766 & ~n91534;
  assign n91559 = n88766 & n91534;
  assign n91560 = ~n91558 & ~n91559;
  assign n91561 = n90774 & n91560;
  assign n91562 = P2_P1_REIP_REG_29_ & n90742;
  assign n91563 = P2_P1_PHYADDRPOINTER_REG_29_ & n90771;
  assign n91564 = ~n91562 & ~n91563;
  assign n91565 = ~n88766 & n90768;
  assign n91566 = n91564 & ~n91565;
  assign n91567 = ~n91550 & ~n91551;
  assign n91568 = n91557 & n91567;
  assign n91569 = ~n91561 & n91568;
  assign n16631 = ~n91566 | ~n91569;
  assign n91571 = P2_P1_REIP_REG_29_ & n91546;
  assign n91572 = ~P2_P1_REIP_REG_30_ & n91571;
  assign n91573 = P2_P1_REIP_REG_30_ & ~n91571;
  assign n91574 = ~n91572 & ~n91573;
  assign n91575 = n90765 & ~n91574;
  assign n91576 = P2_P1_EBX_REG_30_ & ~n90752;
  assign n91577 = n90754 & ~n91574;
  assign n91578 = ~P2_P1_EBX_REG_30_ & n91554;
  assign n91579 = P2_P1_EBX_REG_30_ & ~n91554;
  assign n91580 = ~n91578 & ~n91579;
  assign n91581 = n90756 & n91580;
  assign n91582 = ~n91577 & ~n91581;
  assign n91583 = n88789 & n91559;
  assign n91584 = ~n88789 & ~n91559;
  assign n91585 = ~n91583 & ~n91584;
  assign n91586 = n90774 & n91585;
  assign n91587 = P2_P1_REIP_REG_30_ & n90742;
  assign n91588 = P2_P1_PHYADDRPOINTER_REG_30_ & n90771;
  assign n91589 = ~n91587 & ~n91588;
  assign n91590 = ~n88789 & n90768;
  assign n91591 = n91589 & ~n91590;
  assign n91592 = ~n91575 & ~n91576;
  assign n91593 = n91582 & n91592;
  assign n91594 = ~n91586 & n91593;
  assign n16636 = ~n91591 | ~n91594;
  assign n91596 = P2_P1_REIP_REG_30_ & n91571;
  assign n91597 = ~P2_P1_REIP_REG_31_ & n91596;
  assign n91598 = P2_P1_REIP_REG_31_ & ~n91596;
  assign n91599 = ~n91597 & ~n91598;
  assign n91600 = n90765 & ~n91599;
  assign n91601 = P2_P1_EBX_REG_31_ & ~n90752;
  assign n91602 = n90754 & ~n91599;
  assign n91603 = P2_P1_EBX_REG_31_ & n91578;
  assign n91604 = ~P2_P1_EBX_REG_31_ & ~n91578;
  assign n91605 = ~n91603 & ~n91604;
  assign n91606 = n90756 & ~n91605;
  assign n91607 = ~n91602 & ~n91606;
  assign n91608 = P2_P1_REIP_REG_31_ & n90742;
  assign n91609 = P2_P1_PHYADDRPOINTER_REG_31_ & n90771;
  assign n91610 = ~n91608 & ~n91609;
  assign n91611 = ~n88812 & n90768;
  assign n91612 = n91610 & ~n91611;
  assign n91613 = ~n88812 & n91583;
  assign n91614 = n88812 & ~n91583;
  assign n91615 = ~n91613 & ~n91614;
  assign n91616 = n90774 & ~n91615;
  assign n91617 = ~n91600 & ~n91601;
  assign n91618 = n91607 & n91617;
  assign n91619 = n91612 & n91618;
  assign n16641 = n91616 | ~n91619;
  assign n91621 = ~P2_P1_DATAWIDTH_REG_1_ & ~P2_P1_REIP_REG_1_;
  assign n91622 = ~P2_P1_DATAWIDTH_REG_30_ & ~P2_P1_DATAWIDTH_REG_31_;
  assign n91623 = P2_P1_DATAWIDTH_REG_0_ & P2_P1_DATAWIDTH_REG_1_;
  assign n91624 = ~P2_P1_DATAWIDTH_REG_28_ & ~P2_P1_DATAWIDTH_REG_29_;
  assign n91625 = ~P2_P1_DATAWIDTH_REG_26_ & ~P2_P1_DATAWIDTH_REG_27_;
  assign n91626 = n91622 & ~n91623;
  assign n91627 = n91624 & n91626;
  assign n91628 = n91625 & n91627;
  assign n91629 = ~P2_P1_DATAWIDTH_REG_22_ & ~P2_P1_DATAWIDTH_REG_23_;
  assign n91630 = ~P2_P1_DATAWIDTH_REG_24_ & n91629;
  assign n91631 = ~P2_P1_DATAWIDTH_REG_25_ & n91630;
  assign n91632 = ~P2_P1_DATAWIDTH_REG_18_ & ~P2_P1_DATAWIDTH_REG_19_;
  assign n91633 = ~P2_P1_DATAWIDTH_REG_20_ & n91632;
  assign n91634 = ~P2_P1_DATAWIDTH_REG_21_ & n91633;
  assign n91635 = n91631 & n91634;
  assign n91636 = ~P2_P1_DATAWIDTH_REG_14_ & ~P2_P1_DATAWIDTH_REG_15_;
  assign n91637 = ~P2_P1_DATAWIDTH_REG_16_ & n91636;
  assign n91638 = ~P2_P1_DATAWIDTH_REG_17_ & n91637;
  assign n91639 = ~P2_P1_DATAWIDTH_REG_10_ & ~P2_P1_DATAWIDTH_REG_11_;
  assign n91640 = ~P2_P1_DATAWIDTH_REG_12_ & n91639;
  assign n91641 = ~P2_P1_DATAWIDTH_REG_13_ & n91640;
  assign n91642 = n91638 & n91641;
  assign n91643 = ~P2_P1_DATAWIDTH_REG_6_ & ~P2_P1_DATAWIDTH_REG_7_;
  assign n91644 = ~P2_P1_DATAWIDTH_REG_8_ & n91643;
  assign n91645 = ~P2_P1_DATAWIDTH_REG_9_ & n91644;
  assign n91646 = ~P2_P1_DATAWIDTH_REG_2_ & ~P2_P1_DATAWIDTH_REG_3_;
  assign n91647 = ~P2_P1_DATAWIDTH_REG_4_ & n91646;
  assign n91648 = ~P2_P1_DATAWIDTH_REG_5_ & n91647;
  assign n91649 = n91645 & n91648;
  assign n91650 = n91628 & n91635;
  assign n91651 = n91642 & n91650;
  assign n91652 = n91649 & n91651;
  assign n91653 = n91621 & n91652;
  assign n91654 = P2_P1_BYTEENABLE_REG_3_ & ~n91652;
  assign n91655 = ~P2_P1_DATAWIDTH_REG_0_ & ~P2_P1_REIP_REG_0_;
  assign n91656 = ~P2_P1_DATAWIDTH_REG_1_ & n91655;
  assign n91657 = n91652 & n91656;
  assign n91658 = ~n91653 & ~n91654;
  assign n16646 = n91657 | ~n91658;
  assign n91660 = P2_P1_REIP_REG_0_ & P2_P1_REIP_REG_1_;
  assign n91661 = P2_P1_DATAWIDTH_REG_0_ & ~P2_P1_REIP_REG_0_;
  assign n91662 = ~P2_P1_DATAWIDTH_REG_0_ & ~P2_P1_DATAWIDTH_REG_1_;
  assign n91663 = ~n91661 & ~n91662;
  assign n91664 = ~P2_P1_REIP_REG_1_ & ~n91663;
  assign n91665 = ~n91660 & ~n91664;
  assign n91666 = n91652 & ~n91665;
  assign n91667 = P2_P1_BYTEENABLE_REG_2_ & ~n91652;
  assign n16651 = n91666 | n91667;
  assign n91669 = P2_P1_REIP_REG_1_ & n91652;
  assign n91670 = P2_P1_BYTEENABLE_REG_1_ & ~n91652;
  assign n91671 = ~n91669 & ~n91670;
  assign n16656 = n91657 | ~n91671;
  assign n91673 = ~P2_P1_REIP_REG_0_ & ~P2_P1_REIP_REG_1_;
  assign n91674 = n91652 & ~n91673;
  assign n91675 = P2_P1_BYTEENABLE_REG_0_ & ~n91652;
  assign n16661 = n91674 | n91675;
  assign n91677 = P2_P1_W_R_N_REG & ~n76415;
  assign n91678 = ~P2_P1_READREQUEST_REG & n76415;
  assign n16666 = n91677 | n91678;
  assign n91680 = n77079 & n77311;
  assign n91681 = ~n77027 & n77311;
  assign n91682 = P2_P1_FLUSH_REG & ~n91681;
  assign n16671 = n91680 | n91682;
  assign n91684 = P2_P1_MORE_REG & ~n91681;
  assign n91685 = ~n77073 & n91681;
  assign n16676 = n91684 | n91685;
  assign n91687 = BS & ~n76632;
  assign n91688 = P2_P1_STATEBS16_REG & n76632;
  assign n91689 = ~P2_P1_STATE_REG_0_ & n76587;
  assign n91690 = ~n91687 & ~n91688;
  assign n16681 = n91689 | ~n91690;
  assign n91692 = ~n76957 & ~n77030;
  assign n91693 = ~n76675 & ~n91692;
  assign n91694 = ~P2_P1_STATEBS16_REG & n76957;
  assign n91695 = ~n76584 & ~n91694;
  assign n91696 = P2_P1_STATE2_REG_2_ & ~n91693;
  assign n91697 = n91695 & n91696;
  assign n91698 = P2_P1_STATE2_REG_0_ & ~n91697;
  assign n91699 = ~n77327 & ~n91698;
  assign n91700 = ~n76584 & n76669;
  assign n91701 = ~n77317 & ~n91700;
  assign n91702 = ~P2_P1_STATE2_REG_0_ & ~n91701;
  assign n91703 = ~n77389 & ~n91702;
  assign n91704 = ~n90741 & n91703;
  assign n91705 = ~n91699 & ~n91704;
  assign n91706 = P2_P1_REQUESTPENDING_REG & n91704;
  assign n16686 = n91705 | n91706;
  assign n91708 = P2_P1_D_C_N_REG & ~n76415;
  assign n91709 = ~P2_P1_CODEFETCH_REG & n76415;
  assign n91710 = ~n91708 & ~n91709;
  assign n16691 = n91689 | ~n91710;
  assign n91712 = P2_P1_MEMORYFETCH_REG & n76415;
  assign n91713 = P2_P1_M_IO_N_REG & ~n76415;
  assign n16696 = n91712 | n91713;
  assign n91715 = P2_P1_STATE2_REG_0_ & n85230;
  assign n91716 = n77026 & n77311;
  assign n91717 = P2_P1_CODEFETCH_REG & ~n91716;
  assign n16701 = n91715 | n91717;
  assign n91719 = P2_P1_STATE_REG_0_ & P2_P1_ADS_N_REG;
  assign n16706 = ~n76632 | n91719;
  assign n91721 = P2_P1_STATE2_REG_2_ & ~n77039;
  assign n91722 = ~n77034 & n91721;
  assign n91723 = ~n85230 & ~n90741;
  assign n91724 = ~n91722 & ~n91723;
  assign n91725 = P2_P1_READREQUEST_REG & n91723;
  assign n16711 = n91724 | n91725;
  assign n91727 = P2_P1_STATE2_REG_2_ & n76956;
  assign n91728 = ~n91723 & ~n91727;
  assign n91729 = P2_P1_MEMORYFETCH_REG & n91723;
  assign n16716 = n91728 | n91729;
  assign n2011 = ~P3_STATE_REG;
  assign n3236 = ~P4_STATE_REG;
  always @ (posedge clock) begin
    P1_BUF1_REG_0_ <= n121;
    P1_BUF1_REG_1_ <= n126;
    P1_BUF1_REG_2_ <= n131;
    P1_BUF1_REG_3_ <= n136;
    P1_BUF1_REG_4_ <= n141;
    P1_BUF1_REG_5_ <= n146;
    P1_BUF1_REG_6_ <= n151;
    P1_BUF1_REG_7_ <= n156;
    P1_BUF1_REG_8_ <= n161;
    P1_BUF1_REG_9_ <= n166;
    P1_BUF1_REG_10_ <= n171;
    P1_BUF1_REG_11_ <= n176;
    P1_BUF1_REG_12_ <= n181;
    P1_BUF1_REG_13_ <= n186;
    P1_BUF1_REG_14_ <= n191;
    P1_BUF1_REG_15_ <= n196;
    P1_BUF1_REG_16_ <= n201;
    P1_BUF1_REG_17_ <= n206;
    P1_BUF1_REG_18_ <= n211;
    P1_BUF1_REG_19_ <= n216;
    P1_BUF1_REG_20_ <= n221;
    P1_BUF1_REG_21_ <= n226;
    P1_BUF1_REG_22_ <= n231;
    P1_BUF1_REG_23_ <= n236;
    P1_BUF1_REG_24_ <= n241;
    P1_BUF1_REG_25_ <= n246;
    P1_BUF1_REG_26_ <= n251;
    P1_BUF1_REG_27_ <= n256;
    P1_BUF1_REG_28_ <= n261;
    P1_BUF1_REG_29_ <= n266;
    P1_BUF1_REG_30_ <= n271;
    P1_BUF1_REG_31_ <= n276;
    P1_BUF2_REG_0_ <= n281;
    P1_BUF2_REG_1_ <= n286;
    P1_BUF2_REG_2_ <= n291;
    P1_BUF2_REG_3_ <= n296;
    P1_BUF2_REG_4_ <= n301;
    P1_BUF2_REG_5_ <= n306;
    P1_BUF2_REG_6_ <= n311;
    P1_BUF2_REG_7_ <= n316;
    P1_BUF2_REG_8_ <= n321;
    P1_BUF2_REG_9_ <= n326;
    P1_BUF2_REG_10_ <= n331;
    P1_BUF2_REG_11_ <= n336;
    P1_BUF2_REG_12_ <= n341;
    P1_BUF2_REG_13_ <= n346;
    P1_BUF2_REG_14_ <= n351;
    P1_BUF2_REG_15_ <= n356;
    P1_BUF2_REG_16_ <= n361;
    P1_BUF2_REG_17_ <= n366;
    P1_BUF2_REG_18_ <= n371;
    P1_BUF2_REG_19_ <= n376;
    P1_BUF2_REG_20_ <= n381;
    P1_BUF2_REG_21_ <= n386;
    P1_BUF2_REG_22_ <= n391;
    P1_BUF2_REG_23_ <= n396;
    P1_BUF2_REG_24_ <= n401;
    P1_BUF2_REG_25_ <= n406;
    P1_BUF2_REG_26_ <= n411;
    P1_BUF2_REG_27_ <= n416;
    P1_BUF2_REG_28_ <= n421;
    P1_BUF2_REG_29_ <= n426;
    P1_BUF2_REG_30_ <= n431;
    P1_BUF2_REG_31_ <= n436;
    P1_READY12_REG <= n441;
    P1_READY21_REG <= n446;
    P1_READY22_REG <= n451;
    P1_READY11_REG <= n456;
    P2_BUF1_REG_0_ <= n461;
    P2_BUF1_REG_1_ <= n466;
    P2_BUF1_REG_2_ <= n471;
    P2_BUF1_REG_3_ <= n476;
    P2_BUF1_REG_4_ <= n481;
    P2_BUF1_REG_5_ <= n486;
    P2_BUF1_REG_6_ <= n491;
    P2_BUF1_REG_7_ <= n496;
    P2_BUF1_REG_8_ <= n501;
    P2_BUF1_REG_9_ <= n506;
    P2_BUF1_REG_10_ <= n511;
    P2_BUF1_REG_11_ <= n516;
    P2_BUF1_REG_12_ <= n521;
    P2_BUF1_REG_13_ <= n526;
    P2_BUF1_REG_14_ <= n531;
    P2_BUF1_REG_15_ <= n536;
    P2_BUF1_REG_16_ <= n541;
    P2_BUF1_REG_17_ <= n546;
    P2_BUF1_REG_18_ <= n551;
    P2_BUF1_REG_19_ <= n556;
    P2_BUF1_REG_20_ <= n561;
    P2_BUF1_REG_21_ <= n566;
    P2_BUF1_REG_22_ <= n571;
    P2_BUF1_REG_23_ <= n576;
    P2_BUF1_REG_24_ <= n581;
    P2_BUF1_REG_25_ <= n586;
    P2_BUF1_REG_26_ <= n591;
    P2_BUF1_REG_27_ <= n596;
    P2_BUF1_REG_28_ <= n601;
    P2_BUF1_REG_29_ <= n606;
    P2_BUF1_REG_30_ <= n611;
    P2_BUF1_REG_31_ <= n616;
    P2_BUF2_REG_0_ <= n621;
    P2_BUF2_REG_1_ <= n626;
    P2_BUF2_REG_2_ <= n631;
    P2_BUF2_REG_3_ <= n636;
    P2_BUF2_REG_4_ <= n641;
    P2_BUF2_REG_5_ <= n646;
    P2_BUF2_REG_6_ <= n651;
    P2_BUF2_REG_7_ <= n656;
    P2_BUF2_REG_8_ <= n661;
    P2_BUF2_REG_9_ <= n666;
    P2_BUF2_REG_10_ <= n671;
    P2_BUF2_REG_11_ <= n676;
    P2_BUF2_REG_12_ <= n681;
    P2_BUF2_REG_13_ <= n686;
    P2_BUF2_REG_14_ <= n691;
    P2_BUF2_REG_15_ <= n696;
    P2_BUF2_REG_16_ <= n701;
    P2_BUF2_REG_17_ <= n706;
    P2_BUF2_REG_18_ <= n711;
    P2_BUF2_REG_19_ <= n716;
    P2_BUF2_REG_20_ <= n721;
    P2_BUF2_REG_21_ <= n726;
    P2_BUF2_REG_22_ <= n731;
    P2_BUF2_REG_23_ <= n736;
    P2_BUF2_REG_24_ <= n741;
    P2_BUF2_REG_25_ <= n746;
    P2_BUF2_REG_26_ <= n751;
    P2_BUF2_REG_27_ <= n756;
    P2_BUF2_REG_28_ <= n761;
    P2_BUF2_REG_29_ <= n766;
    P2_BUF2_REG_30_ <= n771;
    P2_BUF2_REG_31_ <= n776;
    P2_READY12_REG <= n781;
    P2_READY21_REG <= n786;
    P2_READY22_REG <= n791;
    P2_READY11_REG <= n796;
    P3_IR_REG_0_ <= n801;
    P3_IR_REG_1_ <= n806;
    P3_IR_REG_2_ <= n811;
    P3_IR_REG_3_ <= n816;
    P3_IR_REG_4_ <= n821;
    P3_IR_REG_5_ <= n826;
    P3_IR_REG_6_ <= n831;
    P3_IR_REG_7_ <= n836;
    P3_IR_REG_8_ <= n841;
    P3_IR_REG_9_ <= n846;
    P3_IR_REG_10_ <= n851;
    P3_IR_REG_11_ <= n856;
    P3_IR_REG_12_ <= n861;
    P3_IR_REG_13_ <= n866;
    P3_IR_REG_14_ <= n871;
    P3_IR_REG_15_ <= n876;
    P3_IR_REG_16_ <= n881;
    P3_IR_REG_17_ <= n886;
    P3_IR_REG_18_ <= n891;
    P3_IR_REG_19_ <= n896;
    P3_IR_REG_20_ <= n901;
    P3_IR_REG_21_ <= n906;
    P3_IR_REG_22_ <= n911;
    P3_IR_REG_23_ <= n916;
    P3_IR_REG_24_ <= n921;
    P3_IR_REG_25_ <= n926;
    P3_IR_REG_26_ <= n931;
    P3_IR_REG_27_ <= n936;
    P3_IR_REG_28_ <= n941;
    P3_IR_REG_29_ <= n946;
    P3_IR_REG_30_ <= n951;
    P3_IR_REG_31_ <= n956;
    P3_D_REG_0_ <= n961;
    P3_D_REG_1_ <= n966;
    P3_D_REG_2_ <= n971;
    P3_D_REG_3_ <= n976;
    P3_D_REG_4_ <= n981;
    P3_D_REG_5_ <= n986;
    P3_D_REG_6_ <= n991;
    P3_D_REG_7_ <= n996;
    P3_D_REG_8_ <= n1001;
    P3_D_REG_9_ <= n1006;
    P3_D_REG_10_ <= n1011;
    P3_D_REG_11_ <= n1016;
    P3_D_REG_12_ <= n1021;
    P3_D_REG_13_ <= n1026;
    P3_D_REG_14_ <= n1031;
    P3_D_REG_15_ <= n1036;
    P3_D_REG_16_ <= n1041;
    P3_D_REG_17_ <= n1046;
    P3_D_REG_18_ <= n1051;
    P3_D_REG_19_ <= n1056;
    P3_D_REG_20_ <= n1061;
    P3_D_REG_21_ <= n1066;
    P3_D_REG_22_ <= n1071;
    P3_D_REG_23_ <= n1076;
    P3_D_REG_24_ <= n1081;
    P3_D_REG_25_ <= n1086;
    P3_D_REG_26_ <= n1091;
    P3_D_REG_27_ <= n1096;
    P3_D_REG_28_ <= n1101;
    P3_D_REG_29_ <= n1106;
    P3_D_REG_30_ <= n1111;
    P3_D_REG_31_ <= n1116;
    P3_REG0_REG_0_ <= n1121;
    P3_REG0_REG_1_ <= n1126;
    P3_REG0_REG_2_ <= n1131;
    P3_REG0_REG_3_ <= n1136;
    P3_REG0_REG_4_ <= n1141;
    P3_REG0_REG_5_ <= n1146;
    P3_REG0_REG_6_ <= n1151;
    P3_REG0_REG_7_ <= n1156;
    P3_REG0_REG_8_ <= n1161;
    P3_REG0_REG_9_ <= n1166;
    P3_REG0_REG_10_ <= n1171;
    P3_REG0_REG_11_ <= n1176;
    P3_REG0_REG_12_ <= n1181;
    P3_REG0_REG_13_ <= n1186;
    P3_REG0_REG_14_ <= n1191;
    P3_REG0_REG_15_ <= n1196;
    P3_REG0_REG_16_ <= n1201;
    P3_REG0_REG_17_ <= n1206;
    P3_REG0_REG_18_ <= n1211;
    P3_REG0_REG_19_ <= n1216;
    P3_REG0_REG_20_ <= n1221;
    P3_REG0_REG_21_ <= n1226;
    P3_REG0_REG_22_ <= n1231;
    P3_REG0_REG_23_ <= n1236;
    P3_REG0_REG_24_ <= n1241;
    P3_REG0_REG_25_ <= n1246;
    P3_REG0_REG_26_ <= n1251;
    P3_REG0_REG_27_ <= n1256;
    P3_REG0_REG_28_ <= n1261;
    P3_REG0_REG_29_ <= n1266;
    P3_REG0_REG_30_ <= n1271;
    P3_REG0_REG_31_ <= n1276;
    P3_REG1_REG_0_ <= n1281;
    P3_REG1_REG_1_ <= n1286;
    P3_REG1_REG_2_ <= n1291;
    P3_REG1_REG_3_ <= n1296;
    P3_REG1_REG_4_ <= n1301;
    P3_REG1_REG_5_ <= n1306;
    P3_REG1_REG_6_ <= n1311;
    P3_REG1_REG_7_ <= n1316;
    P3_REG1_REG_8_ <= n1321;
    P3_REG1_REG_9_ <= n1326;
    P3_REG1_REG_10_ <= n1331;
    P3_REG1_REG_11_ <= n1336;
    P3_REG1_REG_12_ <= n1341;
    P3_REG1_REG_13_ <= n1346;
    P3_REG1_REG_14_ <= n1351;
    P3_REG1_REG_15_ <= n1356;
    P3_REG1_REG_16_ <= n1361;
    P3_REG1_REG_17_ <= n1366;
    P3_REG1_REG_18_ <= n1371;
    P3_REG1_REG_19_ <= n1376;
    P3_REG1_REG_20_ <= n1381;
    P3_REG1_REG_21_ <= n1386;
    P3_REG1_REG_22_ <= n1391;
    P3_REG1_REG_23_ <= n1396;
    P3_REG1_REG_24_ <= n1401;
    P3_REG1_REG_25_ <= n1406;
    P3_REG1_REG_26_ <= n1411;
    P3_REG1_REG_27_ <= n1416;
    P3_REG1_REG_28_ <= n1421;
    P3_REG1_REG_29_ <= n1426;
    P3_REG1_REG_30_ <= n1431;
    P3_REG1_REG_31_ <= n1436;
    P3_REG2_REG_0_ <= n1441;
    P3_REG2_REG_1_ <= n1446;
    P3_REG2_REG_2_ <= n1451;
    P3_REG2_REG_3_ <= n1456;
    P3_REG2_REG_4_ <= n1461;
    P3_REG2_REG_5_ <= n1466;
    P3_REG2_REG_6_ <= n1471;
    P3_REG2_REG_7_ <= n1476;
    P3_REG2_REG_8_ <= n1481;
    P3_REG2_REG_9_ <= n1486;
    P3_REG2_REG_10_ <= n1491;
    P3_REG2_REG_11_ <= n1496;
    P3_REG2_REG_12_ <= n1501;
    P3_REG2_REG_13_ <= n1506;
    P3_REG2_REG_14_ <= n1511;
    P3_REG2_REG_15_ <= n1516;
    P3_REG2_REG_16_ <= n1521;
    P3_REG2_REG_17_ <= n1526;
    P3_REG2_REG_18_ <= n1531;
    P3_REG2_REG_19_ <= n1536;
    P3_REG2_REG_20_ <= n1541;
    P3_REG2_REG_21_ <= n1546;
    P3_REG2_REG_22_ <= n1551;
    P3_REG2_REG_23_ <= n1556;
    P3_REG2_REG_24_ <= n1561;
    P3_REG2_REG_25_ <= n1566;
    P3_REG2_REG_26_ <= n1571;
    P3_REG2_REG_27_ <= n1576;
    P3_REG2_REG_28_ <= n1581;
    P3_REG2_REG_29_ <= n1586;
    P3_REG2_REG_30_ <= n1591;
    P3_REG2_REG_31_ <= n1596;
    P3_ADDR_REG_19_ <= n1601;
    P3_ADDR_REG_18_ <= n1606;
    P3_ADDR_REG_17_ <= n1611;
    P3_ADDR_REG_16_ <= n1616;
    P3_ADDR_REG_15_ <= n1621;
    P3_ADDR_REG_14_ <= n1626;
    P3_ADDR_REG_13_ <= n1631;
    P3_ADDR_REG_12_ <= n1636;
    P3_ADDR_REG_11_ <= n1641;
    P3_ADDR_REG_10_ <= n1646;
    P3_ADDR_REG_9_ <= n1651;
    P3_ADDR_REG_8_ <= n1656;
    P3_ADDR_REG_7_ <= n1661;
    P3_ADDR_REG_6_ <= n1666;
    P3_ADDR_REG_5_ <= n1671;
    P3_ADDR_REG_4_ <= n1676;
    P3_ADDR_REG_3_ <= n1681;
    P3_ADDR_REG_2_ <= n1686;
    P3_ADDR_REG_1_ <= n1691;
    P3_ADDR_REG_0_ <= n1696;
    P3_DATAO_REG_0_ <= n1701;
    P3_DATAO_REG_1_ <= n1706;
    P3_DATAO_REG_2_ <= n1711;
    P3_DATAO_REG_3_ <= n1716;
    P3_DATAO_REG_4_ <= n1721;
    P3_DATAO_REG_5_ <= n1726;
    P3_DATAO_REG_6_ <= n1731;
    P3_DATAO_REG_7_ <= n1736;
    P3_DATAO_REG_8_ <= n1741;
    P3_DATAO_REG_9_ <= n1746;
    P3_DATAO_REG_10_ <= n1751;
    P3_DATAO_REG_11_ <= n1756;
    P3_DATAO_REG_12_ <= n1761;
    P3_DATAO_REG_13_ <= n1766;
    P3_DATAO_REG_14_ <= n1771;
    P3_DATAO_REG_15_ <= n1776;
    P3_DATAO_REG_16_ <= n1781;
    P3_DATAO_REG_17_ <= n1786;
    P3_DATAO_REG_18_ <= n1791;
    P3_DATAO_REG_19_ <= n1796;
    P3_DATAO_REG_20_ <= n1801;
    P3_DATAO_REG_21_ <= n1806;
    P3_DATAO_REG_22_ <= n1811;
    P3_DATAO_REG_23_ <= n1816;
    P3_DATAO_REG_24_ <= n1821;
    P3_DATAO_REG_25_ <= n1826;
    P3_DATAO_REG_26_ <= n1831;
    P3_DATAO_REG_27_ <= n1836;
    P3_DATAO_REG_28_ <= n1841;
    P3_DATAO_REG_29_ <= n1846;
    P3_DATAO_REG_30_ <= n1851;
    P3_DATAO_REG_31_ <= n1856;
    P3_B_REG <= n1861;
    P3_REG3_REG_15_ <= n1866;
    P3_REG3_REG_26_ <= n1871;
    P3_REG3_REG_6_ <= n1876;
    P3_REG3_REG_18_ <= n1881;
    P3_REG3_REG_2_ <= n1886;
    P3_REG3_REG_11_ <= n1891;
    P3_REG3_REG_22_ <= n1896;
    P3_REG3_REG_13_ <= n1901;
    P3_REG3_REG_20_ <= n1906;
    P3_REG3_REG_0_ <= n1911;
    P3_REG3_REG_9_ <= n1916;
    P3_REG3_REG_4_ <= n1921;
    P3_REG3_REG_24_ <= n1926;
    P3_REG3_REG_17_ <= n1931;
    P3_REG3_REG_5_ <= n1936;
    P3_REG3_REG_16_ <= n1941;
    P3_REG3_REG_25_ <= n1946;
    P3_REG3_REG_12_ <= n1951;
    P3_REG3_REG_21_ <= n1956;
    P3_REG3_REG_1_ <= n1961;
    P3_REG3_REG_8_ <= n1966;
    P3_REG3_REG_28_ <= n1971;
    P3_REG3_REG_19_ <= n1976;
    P3_REG3_REG_3_ <= n1981;
    P3_REG3_REG_10_ <= n1986;
    P3_REG3_REG_23_ <= n1991;
    P3_REG3_REG_14_ <= n1996;
    P3_REG3_REG_27_ <= n2001;
    P3_REG3_REG_7_ <= n2006;
    P3_STATE_REG <= n2011;
    P3_RD_REG <= n2016;
    P3_WR_REG <= n2021;
    P4_IR_REG_0_ <= n2026;
    P4_IR_REG_1_ <= n2031;
    P4_IR_REG_2_ <= n2036;
    P4_IR_REG_3_ <= n2041;
    P4_IR_REG_4_ <= n2046;
    P4_IR_REG_5_ <= n2051;
    P4_IR_REG_6_ <= n2056;
    P4_IR_REG_7_ <= n2061;
    P4_IR_REG_8_ <= n2066;
    P4_IR_REG_9_ <= n2071;
    P4_IR_REG_10_ <= n2076;
    P4_IR_REG_11_ <= n2081;
    P4_IR_REG_12_ <= n2086;
    P4_IR_REG_13_ <= n2091;
    P4_IR_REG_14_ <= n2096;
    P4_IR_REG_15_ <= n2101;
    P4_IR_REG_16_ <= n2106;
    P4_IR_REG_17_ <= n2111;
    P4_IR_REG_18_ <= n2116;
    P4_IR_REG_19_ <= n2121;
    P4_IR_REG_20_ <= n2126;
    P4_IR_REG_21_ <= n2131;
    P4_IR_REG_22_ <= n2136;
    P4_IR_REG_23_ <= n2141;
    P4_IR_REG_24_ <= n2146;
    P4_IR_REG_25_ <= n2151;
    P4_IR_REG_26_ <= n2156;
    P4_IR_REG_27_ <= n2161;
    P4_IR_REG_28_ <= n2166;
    P4_IR_REG_29_ <= n2171;
    P4_IR_REG_30_ <= n2176;
    P4_IR_REG_31_ <= n2181;
    P4_D_REG_0_ <= n2186;
    P4_D_REG_1_ <= n2191;
    P4_D_REG_2_ <= n2196;
    P4_D_REG_3_ <= n2201;
    P4_D_REG_4_ <= n2206;
    P4_D_REG_5_ <= n2211;
    P4_D_REG_6_ <= n2216;
    P4_D_REG_7_ <= n2221;
    P4_D_REG_8_ <= n2226;
    P4_D_REG_9_ <= n2231;
    P4_D_REG_10_ <= n2236;
    P4_D_REG_11_ <= n2241;
    P4_D_REG_12_ <= n2246;
    P4_D_REG_13_ <= n2251;
    P4_D_REG_14_ <= n2256;
    P4_D_REG_15_ <= n2261;
    P4_D_REG_16_ <= n2266;
    P4_D_REG_17_ <= n2271;
    P4_D_REG_18_ <= n2276;
    P4_D_REG_19_ <= n2281;
    P4_D_REG_20_ <= n2286;
    P4_D_REG_21_ <= n2291;
    P4_D_REG_22_ <= n2296;
    P4_D_REG_23_ <= n2301;
    P4_D_REG_24_ <= n2306;
    P4_D_REG_25_ <= n2311;
    P4_D_REG_26_ <= n2316;
    P4_D_REG_27_ <= n2321;
    P4_D_REG_28_ <= n2326;
    P4_D_REG_29_ <= n2331;
    P4_D_REG_30_ <= n2336;
    P4_D_REG_31_ <= n2341;
    P4_REG0_REG_0_ <= n2346;
    P4_REG0_REG_1_ <= n2351;
    P4_REG0_REG_2_ <= n2356;
    P4_REG0_REG_3_ <= n2361;
    P4_REG0_REG_4_ <= n2366;
    P4_REG0_REG_5_ <= n2371;
    P4_REG0_REG_6_ <= n2376;
    P4_REG0_REG_7_ <= n2381;
    P4_REG0_REG_8_ <= n2386;
    P4_REG0_REG_9_ <= n2391;
    P4_REG0_REG_10_ <= n2396;
    P4_REG0_REG_11_ <= n2401;
    P4_REG0_REG_12_ <= n2406;
    P4_REG0_REG_13_ <= n2411;
    P4_REG0_REG_14_ <= n2416;
    P4_REG0_REG_15_ <= n2421;
    P4_REG0_REG_16_ <= n2426;
    P4_REG0_REG_17_ <= n2431;
    P4_REG0_REG_18_ <= n2436;
    P4_REG0_REG_19_ <= n2441;
    P4_REG0_REG_20_ <= n2446;
    P4_REG0_REG_21_ <= n2451;
    P4_REG0_REG_22_ <= n2456;
    P4_REG0_REG_23_ <= n2461;
    P4_REG0_REG_24_ <= n2466;
    P4_REG0_REG_25_ <= n2471;
    P4_REG0_REG_26_ <= n2476;
    P4_REG0_REG_27_ <= n2481;
    P4_REG0_REG_28_ <= n2486;
    P4_REG0_REG_29_ <= n2491;
    P4_REG0_REG_30_ <= n2496;
    P4_REG0_REG_31_ <= n2501;
    P4_REG1_REG_0_ <= n2506;
    P4_REG1_REG_1_ <= n2511;
    P4_REG1_REG_2_ <= n2516;
    P4_REG1_REG_3_ <= n2521;
    P4_REG1_REG_4_ <= n2526;
    P4_REG1_REG_5_ <= n2531;
    P4_REG1_REG_6_ <= n2536;
    P4_REG1_REG_7_ <= n2541;
    P4_REG1_REG_8_ <= n2546;
    P4_REG1_REG_9_ <= n2551;
    P4_REG1_REG_10_ <= n2556;
    P4_REG1_REG_11_ <= n2561;
    P4_REG1_REG_12_ <= n2566;
    P4_REG1_REG_13_ <= n2571;
    P4_REG1_REG_14_ <= n2576;
    P4_REG1_REG_15_ <= n2581;
    P4_REG1_REG_16_ <= n2586;
    P4_REG1_REG_17_ <= n2591;
    P4_REG1_REG_18_ <= n2596;
    P4_REG1_REG_19_ <= n2601;
    P4_REG1_REG_20_ <= n2606;
    P4_REG1_REG_21_ <= n2611;
    P4_REG1_REG_22_ <= n2616;
    P4_REG1_REG_23_ <= n2621;
    P4_REG1_REG_24_ <= n2626;
    P4_REG1_REG_25_ <= n2631;
    P4_REG1_REG_26_ <= n2636;
    P4_REG1_REG_27_ <= n2641;
    P4_REG1_REG_28_ <= n2646;
    P4_REG1_REG_29_ <= n2651;
    P4_REG1_REG_30_ <= n2656;
    P4_REG1_REG_31_ <= n2661;
    P4_REG2_REG_0_ <= n2666;
    P4_REG2_REG_1_ <= n2671;
    P4_REG2_REG_2_ <= n2676;
    P4_REG2_REG_3_ <= n2681;
    P4_REG2_REG_4_ <= n2686;
    P4_REG2_REG_5_ <= n2691;
    P4_REG2_REG_6_ <= n2696;
    P4_REG2_REG_7_ <= n2701;
    P4_REG2_REG_8_ <= n2706;
    P4_REG2_REG_9_ <= n2711;
    P4_REG2_REG_10_ <= n2716;
    P4_REG2_REG_11_ <= n2721;
    P4_REG2_REG_12_ <= n2726;
    P4_REG2_REG_13_ <= n2731;
    P4_REG2_REG_14_ <= n2736;
    P4_REG2_REG_15_ <= n2741;
    P4_REG2_REG_16_ <= n2746;
    P4_REG2_REG_17_ <= n2751;
    P4_REG2_REG_18_ <= n2756;
    P4_REG2_REG_19_ <= n2761;
    P4_REG2_REG_20_ <= n2766;
    P4_REG2_REG_21_ <= n2771;
    P4_REG2_REG_22_ <= n2776;
    P4_REG2_REG_23_ <= n2781;
    P4_REG2_REG_24_ <= n2786;
    P4_REG2_REG_25_ <= n2791;
    P4_REG2_REG_26_ <= n2796;
    P4_REG2_REG_27_ <= n2801;
    P4_REG2_REG_28_ <= n2806;
    P4_REG2_REG_29_ <= n2811;
    P4_REG2_REG_30_ <= n2816;
    P4_REG2_REG_31_ <= n2821;
    P4_ADDR_REG_19_ <= n2826;
    P4_ADDR_REG_18_ <= n2831;
    P4_ADDR_REG_17_ <= n2836;
    P4_ADDR_REG_16_ <= n2841;
    P4_ADDR_REG_15_ <= n2846;
    P4_ADDR_REG_14_ <= n2851;
    P4_ADDR_REG_13_ <= n2856;
    P4_ADDR_REG_12_ <= n2861;
    P4_ADDR_REG_11_ <= n2866;
    P4_ADDR_REG_10_ <= n2871;
    P4_ADDR_REG_9_ <= n2876;
    P4_ADDR_REG_8_ <= n2881;
    P4_ADDR_REG_7_ <= n2886;
    P4_ADDR_REG_6_ <= n2891;
    P4_ADDR_REG_5_ <= n2896;
    P4_ADDR_REG_4_ <= n2901;
    P4_ADDR_REG_3_ <= n2906;
    P4_ADDR_REG_2_ <= n2911;
    P4_ADDR_REG_1_ <= n2916;
    P4_ADDR_REG_0_ <= n2921;
    P4_DATAO_REG_0_ <= n2926;
    P4_DATAO_REG_1_ <= n2931;
    P4_DATAO_REG_2_ <= n2936;
    P4_DATAO_REG_3_ <= n2941;
    P4_DATAO_REG_4_ <= n2946;
    P4_DATAO_REG_5_ <= n2951;
    P4_DATAO_REG_6_ <= n2956;
    P4_DATAO_REG_7_ <= n2961;
    P4_DATAO_REG_8_ <= n2966;
    P4_DATAO_REG_9_ <= n2971;
    P4_DATAO_REG_10_ <= n2976;
    P4_DATAO_REG_11_ <= n2981;
    P4_DATAO_REG_12_ <= n2986;
    P4_DATAO_REG_13_ <= n2991;
    P4_DATAO_REG_14_ <= n2996;
    P4_DATAO_REG_15_ <= n3001;
    P4_DATAO_REG_16_ <= n3006;
    P4_DATAO_REG_17_ <= n3011;
    P4_DATAO_REG_18_ <= n3016;
    P4_DATAO_REG_19_ <= n3021;
    P4_DATAO_REG_20_ <= n3026;
    P4_DATAO_REG_21_ <= n3031;
    P4_DATAO_REG_22_ <= n3036;
    P4_DATAO_REG_23_ <= n3041;
    P4_DATAO_REG_24_ <= n3046;
    P4_DATAO_REG_25_ <= n3051;
    P4_DATAO_REG_26_ <= n3056;
    P4_DATAO_REG_27_ <= n3061;
    P4_DATAO_REG_28_ <= n3066;
    P4_DATAO_REG_29_ <= n3071;
    P4_DATAO_REG_30_ <= n3076;
    P4_DATAO_REG_31_ <= n3081;
    P4_B_REG <= n3086;
    P4_REG3_REG_15_ <= n3091;
    P4_REG3_REG_26_ <= n3096;
    P4_REG3_REG_6_ <= n3101;
    P4_REG3_REG_18_ <= n3106;
    P4_REG3_REG_2_ <= n3111;
    P4_REG3_REG_11_ <= n3116;
    P4_REG3_REG_22_ <= n3121;
    P4_REG3_REG_13_ <= n3126;
    P4_REG3_REG_20_ <= n3131;
    P4_REG3_REG_0_ <= n3136;
    P4_REG3_REG_9_ <= n3141;
    P4_REG3_REG_4_ <= n3146;
    P4_REG3_REG_24_ <= n3151;
    P4_REG3_REG_17_ <= n3156;
    P4_REG3_REG_5_ <= n3161;
    P4_REG3_REG_16_ <= n3166;
    P4_REG3_REG_25_ <= n3171;
    P4_REG3_REG_12_ <= n3176;
    P4_REG3_REG_21_ <= n3181;
    P4_REG3_REG_1_ <= n3186;
    P4_REG3_REG_8_ <= n3191;
    P4_REG3_REG_28_ <= n3196;
    P4_REG3_REG_19_ <= n3201;
    P4_REG3_REG_3_ <= n3206;
    P4_REG3_REG_10_ <= n3211;
    P4_REG3_REG_23_ <= n3216;
    P4_REG3_REG_14_ <= n3221;
    P4_REG3_REG_27_ <= n3226;
    P4_REG3_REG_7_ <= n3231;
    P4_STATE_REG <= n3236;
    P4_RD_REG <= n3241;
    P4_WR_REG <= n3246;
    P1_P3_BE_N_REG_3_ <= n3251;
    P1_P3_BE_N_REG_2_ <= n3256;
    P1_P3_BE_N_REG_1_ <= n3261;
    P1_P3_BE_N_REG_0_ <= n3266;
    P1_P3_ADDRESS_REG_29_ <= n3271;
    P1_P3_ADDRESS_REG_28_ <= n3276;
    P1_P3_ADDRESS_REG_27_ <= n3281;
    P1_P3_ADDRESS_REG_26_ <= n3286;
    P1_P3_ADDRESS_REG_25_ <= n3291;
    P1_P3_ADDRESS_REG_24_ <= n3296;
    P1_P3_ADDRESS_REG_23_ <= n3301;
    P1_P3_ADDRESS_REG_22_ <= n3306;
    P1_P3_ADDRESS_REG_21_ <= n3311;
    P1_P3_ADDRESS_REG_20_ <= n3316;
    P1_P3_ADDRESS_REG_19_ <= n3321;
    P1_P3_ADDRESS_REG_18_ <= n3326;
    P1_P3_ADDRESS_REG_17_ <= n3331;
    P1_P3_ADDRESS_REG_16_ <= n3336;
    P1_P3_ADDRESS_REG_15_ <= n3341;
    P1_P3_ADDRESS_REG_14_ <= n3346;
    P1_P3_ADDRESS_REG_13_ <= n3351;
    P1_P3_ADDRESS_REG_12_ <= n3356;
    P1_P3_ADDRESS_REG_11_ <= n3361;
    P1_P3_ADDRESS_REG_10_ <= n3366;
    P1_P3_ADDRESS_REG_9_ <= n3371;
    P1_P3_ADDRESS_REG_8_ <= n3376;
    P1_P3_ADDRESS_REG_7_ <= n3381;
    P1_P3_ADDRESS_REG_6_ <= n3386;
    P1_P3_ADDRESS_REG_5_ <= n3391;
    P1_P3_ADDRESS_REG_4_ <= n3396;
    P1_P3_ADDRESS_REG_3_ <= n3401;
    P1_P3_ADDRESS_REG_2_ <= n3406;
    P1_P3_ADDRESS_REG_1_ <= n3411;
    P1_P3_ADDRESS_REG_0_ <= n3416;
    P1_P3_STATE_REG_2_ <= n3421;
    P1_P3_STATE_REG_1_ <= n3426;
    P1_P3_STATE_REG_0_ <= n3431;
    P1_P3_DATAWIDTH_REG_0_ <= n3436;
    P1_P3_DATAWIDTH_REG_1_ <= n3441;
    P1_P3_DATAWIDTH_REG_2_ <= n3446;
    P1_P3_DATAWIDTH_REG_3_ <= n3451;
    P1_P3_DATAWIDTH_REG_4_ <= n3456;
    P1_P3_DATAWIDTH_REG_5_ <= n3461;
    P1_P3_DATAWIDTH_REG_6_ <= n3466;
    P1_P3_DATAWIDTH_REG_7_ <= n3471;
    P1_P3_DATAWIDTH_REG_8_ <= n3476;
    P1_P3_DATAWIDTH_REG_9_ <= n3481;
    P1_P3_DATAWIDTH_REG_10_ <= n3486;
    P1_P3_DATAWIDTH_REG_11_ <= n3491;
    P1_P3_DATAWIDTH_REG_12_ <= n3496;
    P1_P3_DATAWIDTH_REG_13_ <= n3501;
    P1_P3_DATAWIDTH_REG_14_ <= n3506;
    P1_P3_DATAWIDTH_REG_15_ <= n3511;
    P1_P3_DATAWIDTH_REG_16_ <= n3516;
    P1_P3_DATAWIDTH_REG_17_ <= n3521;
    P1_P3_DATAWIDTH_REG_18_ <= n3526;
    P1_P3_DATAWIDTH_REG_19_ <= n3531;
    P1_P3_DATAWIDTH_REG_20_ <= n3536;
    P1_P3_DATAWIDTH_REG_21_ <= n3541;
    P1_P3_DATAWIDTH_REG_22_ <= n3546;
    P1_P3_DATAWIDTH_REG_23_ <= n3551;
    P1_P3_DATAWIDTH_REG_24_ <= n3556;
    P1_P3_DATAWIDTH_REG_25_ <= n3561;
    P1_P3_DATAWIDTH_REG_26_ <= n3566;
    P1_P3_DATAWIDTH_REG_27_ <= n3571;
    P1_P3_DATAWIDTH_REG_28_ <= n3576;
    P1_P3_DATAWIDTH_REG_29_ <= n3581;
    P1_P3_DATAWIDTH_REG_30_ <= n3586;
    P1_P3_DATAWIDTH_REG_31_ <= n3591;
    P1_P3_STATE2_REG_3_ <= n3596;
    P1_P3_STATE2_REG_2_ <= n3601;
    P1_P3_STATE2_REG_1_ <= n3606;
    P1_P3_STATE2_REG_0_ <= n3611;
    P1_P3_INSTQUEUE_REG_15__7_ <= n3616;
    P1_P3_INSTQUEUE_REG_15__6_ <= n3621;
    P1_P3_INSTQUEUE_REG_15__5_ <= n3626;
    P1_P3_INSTQUEUE_REG_15__4_ <= n3631;
    P1_P3_INSTQUEUE_REG_15__3_ <= n3636;
    P1_P3_INSTQUEUE_REG_15__2_ <= n3641;
    P1_P3_INSTQUEUE_REG_15__1_ <= n3646;
    P1_P3_INSTQUEUE_REG_15__0_ <= n3651;
    P1_P3_INSTQUEUE_REG_14__7_ <= n3656;
    P1_P3_INSTQUEUE_REG_14__6_ <= n3661;
    P1_P3_INSTQUEUE_REG_14__5_ <= n3666;
    P1_P3_INSTQUEUE_REG_14__4_ <= n3671;
    P1_P3_INSTQUEUE_REG_14__3_ <= n3676;
    P1_P3_INSTQUEUE_REG_14__2_ <= n3681;
    P1_P3_INSTQUEUE_REG_14__1_ <= n3686;
    P1_P3_INSTQUEUE_REG_14__0_ <= n3691;
    P1_P3_INSTQUEUE_REG_13__7_ <= n3696;
    P1_P3_INSTQUEUE_REG_13__6_ <= n3701;
    P1_P3_INSTQUEUE_REG_13__5_ <= n3706;
    P1_P3_INSTQUEUE_REG_13__4_ <= n3711;
    P1_P3_INSTQUEUE_REG_13__3_ <= n3716;
    P1_P3_INSTQUEUE_REG_13__2_ <= n3721;
    P1_P3_INSTQUEUE_REG_13__1_ <= n3726;
    P1_P3_INSTQUEUE_REG_13__0_ <= n3731;
    P1_P3_INSTQUEUE_REG_12__7_ <= n3736;
    P1_P3_INSTQUEUE_REG_12__6_ <= n3741;
    P1_P3_INSTQUEUE_REG_12__5_ <= n3746;
    P1_P3_INSTQUEUE_REG_12__4_ <= n3751;
    P1_P3_INSTQUEUE_REG_12__3_ <= n3756;
    P1_P3_INSTQUEUE_REG_12__2_ <= n3761;
    P1_P3_INSTQUEUE_REG_12__1_ <= n3766;
    P1_P3_INSTQUEUE_REG_12__0_ <= n3771;
    P1_P3_INSTQUEUE_REG_11__7_ <= n3776;
    P1_P3_INSTQUEUE_REG_11__6_ <= n3781;
    P1_P3_INSTQUEUE_REG_11__5_ <= n3786;
    P1_P3_INSTQUEUE_REG_11__4_ <= n3791;
    P1_P3_INSTQUEUE_REG_11__3_ <= n3796;
    P1_P3_INSTQUEUE_REG_11__2_ <= n3801;
    P1_P3_INSTQUEUE_REG_11__1_ <= n3806;
    P1_P3_INSTQUEUE_REG_11__0_ <= n3811;
    P1_P3_INSTQUEUE_REG_10__7_ <= n3816;
    P1_P3_INSTQUEUE_REG_10__6_ <= n3821;
    P1_P3_INSTQUEUE_REG_10__5_ <= n3826;
    P1_P3_INSTQUEUE_REG_10__4_ <= n3831;
    P1_P3_INSTQUEUE_REG_10__3_ <= n3836;
    P1_P3_INSTQUEUE_REG_10__2_ <= n3841;
    P1_P3_INSTQUEUE_REG_10__1_ <= n3846;
    P1_P3_INSTQUEUE_REG_10__0_ <= n3851;
    P1_P3_INSTQUEUE_REG_9__7_ <= n3856;
    P1_P3_INSTQUEUE_REG_9__6_ <= n3861;
    P1_P3_INSTQUEUE_REG_9__5_ <= n3866;
    P1_P3_INSTQUEUE_REG_9__4_ <= n3871;
    P1_P3_INSTQUEUE_REG_9__3_ <= n3876;
    P1_P3_INSTQUEUE_REG_9__2_ <= n3881;
    P1_P3_INSTQUEUE_REG_9__1_ <= n3886;
    P1_P3_INSTQUEUE_REG_9__0_ <= n3891;
    P1_P3_INSTQUEUE_REG_8__7_ <= n3896;
    P1_P3_INSTQUEUE_REG_8__6_ <= n3901;
    P1_P3_INSTQUEUE_REG_8__5_ <= n3906;
    P1_P3_INSTQUEUE_REG_8__4_ <= n3911;
    P1_P3_INSTQUEUE_REG_8__3_ <= n3916;
    P1_P3_INSTQUEUE_REG_8__2_ <= n3921;
    P1_P3_INSTQUEUE_REG_8__1_ <= n3926;
    P1_P3_INSTQUEUE_REG_8__0_ <= n3931;
    P1_P3_INSTQUEUE_REG_7__7_ <= n3936;
    P1_P3_INSTQUEUE_REG_7__6_ <= n3941;
    P1_P3_INSTQUEUE_REG_7__5_ <= n3946;
    P1_P3_INSTQUEUE_REG_7__4_ <= n3951;
    P1_P3_INSTQUEUE_REG_7__3_ <= n3956;
    P1_P3_INSTQUEUE_REG_7__2_ <= n3961;
    P1_P3_INSTQUEUE_REG_7__1_ <= n3966;
    P1_P3_INSTQUEUE_REG_7__0_ <= n3971;
    P1_P3_INSTQUEUE_REG_6__7_ <= n3976;
    P1_P3_INSTQUEUE_REG_6__6_ <= n3981;
    P1_P3_INSTQUEUE_REG_6__5_ <= n3986;
    P1_P3_INSTQUEUE_REG_6__4_ <= n3991;
    P1_P3_INSTQUEUE_REG_6__3_ <= n3996;
    P1_P3_INSTQUEUE_REG_6__2_ <= n4001;
    P1_P3_INSTQUEUE_REG_6__1_ <= n4006;
    P1_P3_INSTQUEUE_REG_6__0_ <= n4011;
    P1_P3_INSTQUEUE_REG_5__7_ <= n4016;
    P1_P3_INSTQUEUE_REG_5__6_ <= n4021;
    P1_P3_INSTQUEUE_REG_5__5_ <= n4026;
    P1_P3_INSTQUEUE_REG_5__4_ <= n4031;
    P1_P3_INSTQUEUE_REG_5__3_ <= n4036;
    P1_P3_INSTQUEUE_REG_5__2_ <= n4041;
    P1_P3_INSTQUEUE_REG_5__1_ <= n4046;
    P1_P3_INSTQUEUE_REG_5__0_ <= n4051;
    P1_P3_INSTQUEUE_REG_4__7_ <= n4056;
    P1_P3_INSTQUEUE_REG_4__6_ <= n4061;
    P1_P3_INSTQUEUE_REG_4__5_ <= n4066;
    P1_P3_INSTQUEUE_REG_4__4_ <= n4071;
    P1_P3_INSTQUEUE_REG_4__3_ <= n4076;
    P1_P3_INSTQUEUE_REG_4__2_ <= n4081;
    P1_P3_INSTQUEUE_REG_4__1_ <= n4086;
    P1_P3_INSTQUEUE_REG_4__0_ <= n4091;
    P1_P3_INSTQUEUE_REG_3__7_ <= n4096;
    P1_P3_INSTQUEUE_REG_3__6_ <= n4101;
    P1_P3_INSTQUEUE_REG_3__5_ <= n4106;
    P1_P3_INSTQUEUE_REG_3__4_ <= n4111;
    P1_P3_INSTQUEUE_REG_3__3_ <= n4116;
    P1_P3_INSTQUEUE_REG_3__2_ <= n4121;
    P1_P3_INSTQUEUE_REG_3__1_ <= n4126;
    P1_P3_INSTQUEUE_REG_3__0_ <= n4131;
    P1_P3_INSTQUEUE_REG_2__7_ <= n4136;
    P1_P3_INSTQUEUE_REG_2__6_ <= n4141;
    P1_P3_INSTQUEUE_REG_2__5_ <= n4146;
    P1_P3_INSTQUEUE_REG_2__4_ <= n4151;
    P1_P3_INSTQUEUE_REG_2__3_ <= n4156;
    P1_P3_INSTQUEUE_REG_2__2_ <= n4161;
    P1_P3_INSTQUEUE_REG_2__1_ <= n4166;
    P1_P3_INSTQUEUE_REG_2__0_ <= n4171;
    P1_P3_INSTQUEUE_REG_1__7_ <= n4176;
    P1_P3_INSTQUEUE_REG_1__6_ <= n4181;
    P1_P3_INSTQUEUE_REG_1__5_ <= n4186;
    P1_P3_INSTQUEUE_REG_1__4_ <= n4191;
    P1_P3_INSTQUEUE_REG_1__3_ <= n4196;
    P1_P3_INSTQUEUE_REG_1__2_ <= n4201;
    P1_P3_INSTQUEUE_REG_1__1_ <= n4206;
    P1_P3_INSTQUEUE_REG_1__0_ <= n4211;
    P1_P3_INSTQUEUE_REG_0__7_ <= n4216;
    P1_P3_INSTQUEUE_REG_0__6_ <= n4221;
    P1_P3_INSTQUEUE_REG_0__5_ <= n4226;
    P1_P3_INSTQUEUE_REG_0__4_ <= n4231;
    P1_P3_INSTQUEUE_REG_0__3_ <= n4236;
    P1_P3_INSTQUEUE_REG_0__2_ <= n4241;
    P1_P3_INSTQUEUE_REG_0__1_ <= n4246;
    P1_P3_INSTQUEUE_REG_0__0_ <= n4251;
    P1_P3_INSTQUEUERD_ADDR_REG_4_ <= n4256;
    P1_P3_INSTQUEUERD_ADDR_REG_3_ <= n4261;
    P1_P3_INSTQUEUERD_ADDR_REG_2_ <= n4266;
    P1_P3_INSTQUEUERD_ADDR_REG_1_ <= n4271;
    P1_P3_INSTQUEUERD_ADDR_REG_0_ <= n4276;
    P1_P3_INSTQUEUEWR_ADDR_REG_4_ <= n4281;
    P1_P3_INSTQUEUEWR_ADDR_REG_3_ <= n4286;
    P1_P3_INSTQUEUEWR_ADDR_REG_2_ <= n4291;
    P1_P3_INSTQUEUEWR_ADDR_REG_1_ <= n4296;
    P1_P3_INSTQUEUEWR_ADDR_REG_0_ <= n4301;
    P1_P3_INSTADDRPOINTER_REG_0_ <= n4306;
    P1_P3_INSTADDRPOINTER_REG_1_ <= n4311;
    P1_P3_INSTADDRPOINTER_REG_2_ <= n4316;
    P1_P3_INSTADDRPOINTER_REG_3_ <= n4321;
    P1_P3_INSTADDRPOINTER_REG_4_ <= n4326;
    P1_P3_INSTADDRPOINTER_REG_5_ <= n4331;
    P1_P3_INSTADDRPOINTER_REG_6_ <= n4336;
    P1_P3_INSTADDRPOINTER_REG_7_ <= n4341;
    P1_P3_INSTADDRPOINTER_REG_8_ <= n4346;
    P1_P3_INSTADDRPOINTER_REG_9_ <= n4351;
    P1_P3_INSTADDRPOINTER_REG_10_ <= n4356;
    P1_P3_INSTADDRPOINTER_REG_11_ <= n4361;
    P1_P3_INSTADDRPOINTER_REG_12_ <= n4366;
    P1_P3_INSTADDRPOINTER_REG_13_ <= n4371;
    P1_P3_INSTADDRPOINTER_REG_14_ <= n4376;
    P1_P3_INSTADDRPOINTER_REG_15_ <= n4381;
    P1_P3_INSTADDRPOINTER_REG_16_ <= n4386;
    P1_P3_INSTADDRPOINTER_REG_17_ <= n4391;
    P1_P3_INSTADDRPOINTER_REG_18_ <= n4396;
    P1_P3_INSTADDRPOINTER_REG_19_ <= n4401;
    P1_P3_INSTADDRPOINTER_REG_20_ <= n4406;
    P1_P3_INSTADDRPOINTER_REG_21_ <= n4411;
    P1_P3_INSTADDRPOINTER_REG_22_ <= n4416;
    P1_P3_INSTADDRPOINTER_REG_23_ <= n4421;
    P1_P3_INSTADDRPOINTER_REG_24_ <= n4426;
    P1_P3_INSTADDRPOINTER_REG_25_ <= n4431;
    P1_P3_INSTADDRPOINTER_REG_26_ <= n4436;
    P1_P3_INSTADDRPOINTER_REG_27_ <= n4441;
    P1_P3_INSTADDRPOINTER_REG_28_ <= n4446;
    P1_P3_INSTADDRPOINTER_REG_29_ <= n4451;
    P1_P3_INSTADDRPOINTER_REG_30_ <= n4456;
    P1_P3_INSTADDRPOINTER_REG_31_ <= n4461;
    P1_P3_PHYADDRPOINTER_REG_0_ <= n4466;
    P1_P3_PHYADDRPOINTER_REG_1_ <= n4471;
    P1_P3_PHYADDRPOINTER_REG_2_ <= n4476;
    P1_P3_PHYADDRPOINTER_REG_3_ <= n4481;
    P1_P3_PHYADDRPOINTER_REG_4_ <= n4486;
    P1_P3_PHYADDRPOINTER_REG_5_ <= n4491;
    P1_P3_PHYADDRPOINTER_REG_6_ <= n4496;
    P1_P3_PHYADDRPOINTER_REG_7_ <= n4501;
    P1_P3_PHYADDRPOINTER_REG_8_ <= n4506;
    P1_P3_PHYADDRPOINTER_REG_9_ <= n4511;
    P1_P3_PHYADDRPOINTER_REG_10_ <= n4516;
    P1_P3_PHYADDRPOINTER_REG_11_ <= n4521;
    P1_P3_PHYADDRPOINTER_REG_12_ <= n4526;
    P1_P3_PHYADDRPOINTER_REG_13_ <= n4531;
    P1_P3_PHYADDRPOINTER_REG_14_ <= n4536;
    P1_P3_PHYADDRPOINTER_REG_15_ <= n4541;
    P1_P3_PHYADDRPOINTER_REG_16_ <= n4546;
    P1_P3_PHYADDRPOINTER_REG_17_ <= n4551;
    P1_P3_PHYADDRPOINTER_REG_18_ <= n4556;
    P1_P3_PHYADDRPOINTER_REG_19_ <= n4561;
    P1_P3_PHYADDRPOINTER_REG_20_ <= n4566;
    P1_P3_PHYADDRPOINTER_REG_21_ <= n4571;
    P1_P3_PHYADDRPOINTER_REG_22_ <= n4576;
    P1_P3_PHYADDRPOINTER_REG_23_ <= n4581;
    P1_P3_PHYADDRPOINTER_REG_24_ <= n4586;
    P1_P3_PHYADDRPOINTER_REG_25_ <= n4591;
    P1_P3_PHYADDRPOINTER_REG_26_ <= n4596;
    P1_P3_PHYADDRPOINTER_REG_27_ <= n4601;
    P1_P3_PHYADDRPOINTER_REG_28_ <= n4606;
    P1_P3_PHYADDRPOINTER_REG_29_ <= n4611;
    P1_P3_PHYADDRPOINTER_REG_30_ <= n4616;
    P1_P3_PHYADDRPOINTER_REG_31_ <= n4621;
    P1_P3_LWORD_REG_15_ <= n4626;
    P1_P3_LWORD_REG_14_ <= n4631;
    P1_P3_LWORD_REG_13_ <= n4636;
    P1_P3_LWORD_REG_12_ <= n4641;
    P1_P3_LWORD_REG_11_ <= n4646;
    P1_P3_LWORD_REG_10_ <= n4651;
    P1_P3_LWORD_REG_9_ <= n4656;
    P1_P3_LWORD_REG_8_ <= n4661;
    P1_P3_LWORD_REG_7_ <= n4666;
    P1_P3_LWORD_REG_6_ <= n4671;
    P1_P3_LWORD_REG_5_ <= n4676;
    P1_P3_LWORD_REG_4_ <= n4681;
    P1_P3_LWORD_REG_3_ <= n4686;
    P1_P3_LWORD_REG_2_ <= n4691;
    P1_P3_LWORD_REG_1_ <= n4696;
    P1_P3_LWORD_REG_0_ <= n4701;
    P1_P3_UWORD_REG_14_ <= n4706;
    P1_P3_UWORD_REG_13_ <= n4711;
    P1_P3_UWORD_REG_12_ <= n4716;
    P1_P3_UWORD_REG_11_ <= n4721;
    P1_P3_UWORD_REG_10_ <= n4726;
    P1_P3_UWORD_REG_9_ <= n4731;
    P1_P3_UWORD_REG_8_ <= n4736;
    P1_P3_UWORD_REG_7_ <= n4741;
    P1_P3_UWORD_REG_6_ <= n4746;
    P1_P3_UWORD_REG_5_ <= n4751;
    P1_P3_UWORD_REG_4_ <= n4756;
    P1_P3_UWORD_REG_3_ <= n4761;
    P1_P3_UWORD_REG_2_ <= n4766;
    P1_P3_UWORD_REG_1_ <= n4771;
    P1_P3_UWORD_REG_0_ <= n4776;
    P1_P3_DATAO_REG_0_ <= n4781;
    P1_P3_DATAO_REG_1_ <= n4786;
    P1_P3_DATAO_REG_2_ <= n4791;
    P1_P3_DATAO_REG_3_ <= n4796;
    P1_P3_DATAO_REG_4_ <= n4801;
    P1_P3_DATAO_REG_5_ <= n4806;
    P1_P3_DATAO_REG_6_ <= n4811;
    P1_P3_DATAO_REG_7_ <= n4816;
    P1_P3_DATAO_REG_8_ <= n4821;
    P1_P3_DATAO_REG_9_ <= n4826;
    P1_P3_DATAO_REG_10_ <= n4831;
    P1_P3_DATAO_REG_11_ <= n4836;
    P1_P3_DATAO_REG_12_ <= n4841;
    P1_P3_DATAO_REG_13_ <= n4846;
    P1_P3_DATAO_REG_14_ <= n4851;
    P1_P3_DATAO_REG_15_ <= n4856;
    P1_P3_DATAO_REG_16_ <= n4861;
    P1_P3_DATAO_REG_17_ <= n4866;
    P1_P3_DATAO_REG_18_ <= n4871;
    P1_P3_DATAO_REG_19_ <= n4876;
    P1_P3_DATAO_REG_20_ <= n4881;
    P1_P3_DATAO_REG_21_ <= n4886;
    P1_P3_DATAO_REG_22_ <= n4891;
    P1_P3_DATAO_REG_23_ <= n4896;
    P1_P3_DATAO_REG_24_ <= n4901;
    P1_P3_DATAO_REG_25_ <= n4906;
    P1_P3_DATAO_REG_26_ <= n4911;
    P1_P3_DATAO_REG_27_ <= n4916;
    P1_P3_DATAO_REG_28_ <= n4921;
    P1_P3_DATAO_REG_29_ <= n4926;
    P1_P3_DATAO_REG_30_ <= n4931;
    P1_P3_DATAO_REG_31_ <= n4936;
    P1_P3_EAX_REG_0_ <= n4941;
    P1_P3_EAX_REG_1_ <= n4946;
    P1_P3_EAX_REG_2_ <= n4951;
    P1_P3_EAX_REG_3_ <= n4956;
    P1_P3_EAX_REG_4_ <= n4961;
    P1_P3_EAX_REG_5_ <= n4966;
    P1_P3_EAX_REG_6_ <= n4971;
    P1_P3_EAX_REG_7_ <= n4976;
    P1_P3_EAX_REG_8_ <= n4981;
    P1_P3_EAX_REG_9_ <= n4986;
    P1_P3_EAX_REG_10_ <= n4991;
    P1_P3_EAX_REG_11_ <= n4996;
    P1_P3_EAX_REG_12_ <= n5001;
    P1_P3_EAX_REG_13_ <= n5006;
    P1_P3_EAX_REG_14_ <= n5011;
    P1_P3_EAX_REG_15_ <= n5016;
    P1_P3_EAX_REG_16_ <= n5021;
    P1_P3_EAX_REG_17_ <= n5026;
    P1_P3_EAX_REG_18_ <= n5031;
    P1_P3_EAX_REG_19_ <= n5036;
    P1_P3_EAX_REG_20_ <= n5041;
    P1_P3_EAX_REG_21_ <= n5046;
    P1_P3_EAX_REG_22_ <= n5051;
    P1_P3_EAX_REG_23_ <= n5056;
    P1_P3_EAX_REG_24_ <= n5061;
    P1_P3_EAX_REG_25_ <= n5066;
    P1_P3_EAX_REG_26_ <= n5071;
    P1_P3_EAX_REG_27_ <= n5076;
    P1_P3_EAX_REG_28_ <= n5081;
    P1_P3_EAX_REG_29_ <= n5086;
    P1_P3_EAX_REG_30_ <= n5091;
    P1_P3_EAX_REG_31_ <= n5096;
    P1_P3_EBX_REG_0_ <= n5101;
    P1_P3_EBX_REG_1_ <= n5106;
    P1_P3_EBX_REG_2_ <= n5111;
    P1_P3_EBX_REG_3_ <= n5116;
    P1_P3_EBX_REG_4_ <= n5121;
    P1_P3_EBX_REG_5_ <= n5126;
    P1_P3_EBX_REG_6_ <= n5131;
    P1_P3_EBX_REG_7_ <= n5136;
    P1_P3_EBX_REG_8_ <= n5141;
    P1_P3_EBX_REG_9_ <= n5146;
    P1_P3_EBX_REG_10_ <= n5151;
    P1_P3_EBX_REG_11_ <= n5156;
    P1_P3_EBX_REG_12_ <= n5161;
    P1_P3_EBX_REG_13_ <= n5166;
    P1_P3_EBX_REG_14_ <= n5171;
    P1_P3_EBX_REG_15_ <= n5176;
    P1_P3_EBX_REG_16_ <= n5181;
    P1_P3_EBX_REG_17_ <= n5186;
    P1_P3_EBX_REG_18_ <= n5191;
    P1_P3_EBX_REG_19_ <= n5196;
    P1_P3_EBX_REG_20_ <= n5201;
    P1_P3_EBX_REG_21_ <= n5206;
    P1_P3_EBX_REG_22_ <= n5211;
    P1_P3_EBX_REG_23_ <= n5216;
    P1_P3_EBX_REG_24_ <= n5221;
    P1_P3_EBX_REG_25_ <= n5226;
    P1_P3_EBX_REG_26_ <= n5231;
    P1_P3_EBX_REG_27_ <= n5236;
    P1_P3_EBX_REG_28_ <= n5241;
    P1_P3_EBX_REG_29_ <= n5246;
    P1_P3_EBX_REG_30_ <= n5251;
    P1_P3_EBX_REG_31_ <= n5256;
    P1_P3_REIP_REG_0_ <= n5261;
    P1_P3_REIP_REG_1_ <= n5266;
    P1_P3_REIP_REG_2_ <= n5271;
    P1_P3_REIP_REG_3_ <= n5276;
    P1_P3_REIP_REG_4_ <= n5281;
    P1_P3_REIP_REG_5_ <= n5286;
    P1_P3_REIP_REG_6_ <= n5291;
    P1_P3_REIP_REG_7_ <= n5296;
    P1_P3_REIP_REG_8_ <= n5301;
    P1_P3_REIP_REG_9_ <= n5306;
    P1_P3_REIP_REG_10_ <= n5311;
    P1_P3_REIP_REG_11_ <= n5316;
    P1_P3_REIP_REG_12_ <= n5321;
    P1_P3_REIP_REG_13_ <= n5326;
    P1_P3_REIP_REG_14_ <= n5331;
    P1_P3_REIP_REG_15_ <= n5336;
    P1_P3_REIP_REG_16_ <= n5341;
    P1_P3_REIP_REG_17_ <= n5346;
    P1_P3_REIP_REG_18_ <= n5351;
    P1_P3_REIP_REG_19_ <= n5356;
    P1_P3_REIP_REG_20_ <= n5361;
    P1_P3_REIP_REG_21_ <= n5366;
    P1_P3_REIP_REG_22_ <= n5371;
    P1_P3_REIP_REG_23_ <= n5376;
    P1_P3_REIP_REG_24_ <= n5381;
    P1_P3_REIP_REG_25_ <= n5386;
    P1_P3_REIP_REG_26_ <= n5391;
    P1_P3_REIP_REG_27_ <= n5396;
    P1_P3_REIP_REG_28_ <= n5401;
    P1_P3_REIP_REG_29_ <= n5406;
    P1_P3_REIP_REG_30_ <= n5411;
    P1_P3_REIP_REG_31_ <= n5416;
    P1_P3_BYTEENABLE_REG_3_ <= n5421;
    P1_P3_BYTEENABLE_REG_2_ <= n5426;
    P1_P3_BYTEENABLE_REG_1_ <= n5431;
    P1_P3_BYTEENABLE_REG_0_ <= n5436;
    P1_P3_W_R_N_REG <= n5441;
    P1_P3_FLUSH_REG <= n5446;
    P1_P3_MORE_REG <= n5451;
    P1_P3_STATEBS16_REG <= n5456;
    P1_P3_REQUESTPENDING_REG <= n5461;
    P1_P3_D_C_N_REG <= n5466;
    P1_P3_M_IO_N_REG <= n5471;
    P1_P3_CODEFETCH_REG <= n5476;
    P1_P3_ADS_N_REG <= n5481;
    P1_P3_READREQUEST_REG <= n5486;
    P1_P3_MEMORYFETCH_REG <= n5491;
    P1_P2_BE_N_REG_3_ <= n5496;
    P1_P2_BE_N_REG_2_ <= n5501;
    P1_P2_BE_N_REG_1_ <= n5506;
    P1_P2_BE_N_REG_0_ <= n5511;
    P1_P2_ADDRESS_REG_29_ <= n5516;
    P1_P2_ADDRESS_REG_28_ <= n5521;
    P1_P2_ADDRESS_REG_27_ <= n5526;
    P1_P2_ADDRESS_REG_26_ <= n5531;
    P1_P2_ADDRESS_REG_25_ <= n5536;
    P1_P2_ADDRESS_REG_24_ <= n5541;
    P1_P2_ADDRESS_REG_23_ <= n5546;
    P1_P2_ADDRESS_REG_22_ <= n5551;
    P1_P2_ADDRESS_REG_21_ <= n5556;
    P1_P2_ADDRESS_REG_20_ <= n5561;
    P1_P2_ADDRESS_REG_19_ <= n5566;
    P1_P2_ADDRESS_REG_18_ <= n5571;
    P1_P2_ADDRESS_REG_17_ <= n5576;
    P1_P2_ADDRESS_REG_16_ <= n5581;
    P1_P2_ADDRESS_REG_15_ <= n5586;
    P1_P2_ADDRESS_REG_14_ <= n5591;
    P1_P2_ADDRESS_REG_13_ <= n5596;
    P1_P2_ADDRESS_REG_12_ <= n5601;
    P1_P2_ADDRESS_REG_11_ <= n5606;
    P1_P2_ADDRESS_REG_10_ <= n5611;
    P1_P2_ADDRESS_REG_9_ <= n5616;
    P1_P2_ADDRESS_REG_8_ <= n5621;
    P1_P2_ADDRESS_REG_7_ <= n5626;
    P1_P2_ADDRESS_REG_6_ <= n5631;
    P1_P2_ADDRESS_REG_5_ <= n5636;
    P1_P2_ADDRESS_REG_4_ <= n5641;
    P1_P2_ADDRESS_REG_3_ <= n5646;
    P1_P2_ADDRESS_REG_2_ <= n5651;
    P1_P2_ADDRESS_REG_1_ <= n5656;
    P1_P2_ADDRESS_REG_0_ <= n5661;
    P1_P2_STATE_REG_2_ <= n5666;
    P1_P2_STATE_REG_1_ <= n5671;
    P1_P2_STATE_REG_0_ <= n5676;
    P1_P2_DATAWIDTH_REG_0_ <= n5681;
    P1_P2_DATAWIDTH_REG_1_ <= n5686;
    P1_P2_DATAWIDTH_REG_2_ <= n5691;
    P1_P2_DATAWIDTH_REG_3_ <= n5696;
    P1_P2_DATAWIDTH_REG_4_ <= n5701;
    P1_P2_DATAWIDTH_REG_5_ <= n5706;
    P1_P2_DATAWIDTH_REG_6_ <= n5711;
    P1_P2_DATAWIDTH_REG_7_ <= n5716;
    P1_P2_DATAWIDTH_REG_8_ <= n5721;
    P1_P2_DATAWIDTH_REG_9_ <= n5726;
    P1_P2_DATAWIDTH_REG_10_ <= n5731;
    P1_P2_DATAWIDTH_REG_11_ <= n5736;
    P1_P2_DATAWIDTH_REG_12_ <= n5741;
    P1_P2_DATAWIDTH_REG_13_ <= n5746;
    P1_P2_DATAWIDTH_REG_14_ <= n5751;
    P1_P2_DATAWIDTH_REG_15_ <= n5756;
    P1_P2_DATAWIDTH_REG_16_ <= n5761;
    P1_P2_DATAWIDTH_REG_17_ <= n5766;
    P1_P2_DATAWIDTH_REG_18_ <= n5771;
    P1_P2_DATAWIDTH_REG_19_ <= n5776;
    P1_P2_DATAWIDTH_REG_20_ <= n5781;
    P1_P2_DATAWIDTH_REG_21_ <= n5786;
    P1_P2_DATAWIDTH_REG_22_ <= n5791;
    P1_P2_DATAWIDTH_REG_23_ <= n5796;
    P1_P2_DATAWIDTH_REG_24_ <= n5801;
    P1_P2_DATAWIDTH_REG_25_ <= n5806;
    P1_P2_DATAWIDTH_REG_26_ <= n5811;
    P1_P2_DATAWIDTH_REG_27_ <= n5816;
    P1_P2_DATAWIDTH_REG_28_ <= n5821;
    P1_P2_DATAWIDTH_REG_29_ <= n5826;
    P1_P2_DATAWIDTH_REG_30_ <= n5831;
    P1_P2_DATAWIDTH_REG_31_ <= n5836;
    P1_P2_STATE2_REG_3_ <= n5841;
    P1_P2_STATE2_REG_2_ <= n5846;
    P1_P2_STATE2_REG_1_ <= n5851;
    P1_P2_STATE2_REG_0_ <= n5856;
    P1_P2_INSTQUEUE_REG_15__7_ <= n5861;
    P1_P2_INSTQUEUE_REG_15__6_ <= n5866;
    P1_P2_INSTQUEUE_REG_15__5_ <= n5871;
    P1_P2_INSTQUEUE_REG_15__4_ <= n5876;
    P1_P2_INSTQUEUE_REG_15__3_ <= n5881;
    P1_P2_INSTQUEUE_REG_15__2_ <= n5886;
    P1_P2_INSTQUEUE_REG_15__1_ <= n5891;
    P1_P2_INSTQUEUE_REG_15__0_ <= n5896;
    P1_P2_INSTQUEUE_REG_14__7_ <= n5901;
    P1_P2_INSTQUEUE_REG_14__6_ <= n5906;
    P1_P2_INSTQUEUE_REG_14__5_ <= n5911;
    P1_P2_INSTQUEUE_REG_14__4_ <= n5916;
    P1_P2_INSTQUEUE_REG_14__3_ <= n5921;
    P1_P2_INSTQUEUE_REG_14__2_ <= n5926;
    P1_P2_INSTQUEUE_REG_14__1_ <= n5931;
    P1_P2_INSTQUEUE_REG_14__0_ <= n5936;
    P1_P2_INSTQUEUE_REG_13__7_ <= n5941;
    P1_P2_INSTQUEUE_REG_13__6_ <= n5946;
    P1_P2_INSTQUEUE_REG_13__5_ <= n5951;
    P1_P2_INSTQUEUE_REG_13__4_ <= n5956;
    P1_P2_INSTQUEUE_REG_13__3_ <= n5961;
    P1_P2_INSTQUEUE_REG_13__2_ <= n5966;
    P1_P2_INSTQUEUE_REG_13__1_ <= n5971;
    P1_P2_INSTQUEUE_REG_13__0_ <= n5976;
    P1_P2_INSTQUEUE_REG_12__7_ <= n5981;
    P1_P2_INSTQUEUE_REG_12__6_ <= n5986;
    P1_P2_INSTQUEUE_REG_12__5_ <= n5991;
    P1_P2_INSTQUEUE_REG_12__4_ <= n5996;
    P1_P2_INSTQUEUE_REG_12__3_ <= n6001;
    P1_P2_INSTQUEUE_REG_12__2_ <= n6006;
    P1_P2_INSTQUEUE_REG_12__1_ <= n6011;
    P1_P2_INSTQUEUE_REG_12__0_ <= n6016;
    P1_P2_INSTQUEUE_REG_11__7_ <= n6021;
    P1_P2_INSTQUEUE_REG_11__6_ <= n6026;
    P1_P2_INSTQUEUE_REG_11__5_ <= n6031;
    P1_P2_INSTQUEUE_REG_11__4_ <= n6036;
    P1_P2_INSTQUEUE_REG_11__3_ <= n6041;
    P1_P2_INSTQUEUE_REG_11__2_ <= n6046;
    P1_P2_INSTQUEUE_REG_11__1_ <= n6051;
    P1_P2_INSTQUEUE_REG_11__0_ <= n6056;
    P1_P2_INSTQUEUE_REG_10__7_ <= n6061;
    P1_P2_INSTQUEUE_REG_10__6_ <= n6066;
    P1_P2_INSTQUEUE_REG_10__5_ <= n6071;
    P1_P2_INSTQUEUE_REG_10__4_ <= n6076;
    P1_P2_INSTQUEUE_REG_10__3_ <= n6081;
    P1_P2_INSTQUEUE_REG_10__2_ <= n6086;
    P1_P2_INSTQUEUE_REG_10__1_ <= n6091;
    P1_P2_INSTQUEUE_REG_10__0_ <= n6096;
    P1_P2_INSTQUEUE_REG_9__7_ <= n6101;
    P1_P2_INSTQUEUE_REG_9__6_ <= n6106;
    P1_P2_INSTQUEUE_REG_9__5_ <= n6111;
    P1_P2_INSTQUEUE_REG_9__4_ <= n6116;
    P1_P2_INSTQUEUE_REG_9__3_ <= n6121;
    P1_P2_INSTQUEUE_REG_9__2_ <= n6126;
    P1_P2_INSTQUEUE_REG_9__1_ <= n6131;
    P1_P2_INSTQUEUE_REG_9__0_ <= n6136;
    P1_P2_INSTQUEUE_REG_8__7_ <= n6141;
    P1_P2_INSTQUEUE_REG_8__6_ <= n6146;
    P1_P2_INSTQUEUE_REG_8__5_ <= n6151;
    P1_P2_INSTQUEUE_REG_8__4_ <= n6156;
    P1_P2_INSTQUEUE_REG_8__3_ <= n6161;
    P1_P2_INSTQUEUE_REG_8__2_ <= n6166;
    P1_P2_INSTQUEUE_REG_8__1_ <= n6171;
    P1_P2_INSTQUEUE_REG_8__0_ <= n6176;
    P1_P2_INSTQUEUE_REG_7__7_ <= n6181;
    P1_P2_INSTQUEUE_REG_7__6_ <= n6186;
    P1_P2_INSTQUEUE_REG_7__5_ <= n6191;
    P1_P2_INSTQUEUE_REG_7__4_ <= n6196;
    P1_P2_INSTQUEUE_REG_7__3_ <= n6201;
    P1_P2_INSTQUEUE_REG_7__2_ <= n6206;
    P1_P2_INSTQUEUE_REG_7__1_ <= n6211;
    P1_P2_INSTQUEUE_REG_7__0_ <= n6216;
    P1_P2_INSTQUEUE_REG_6__7_ <= n6221;
    P1_P2_INSTQUEUE_REG_6__6_ <= n6226;
    P1_P2_INSTQUEUE_REG_6__5_ <= n6231;
    P1_P2_INSTQUEUE_REG_6__4_ <= n6236;
    P1_P2_INSTQUEUE_REG_6__3_ <= n6241;
    P1_P2_INSTQUEUE_REG_6__2_ <= n6246;
    P1_P2_INSTQUEUE_REG_6__1_ <= n6251;
    P1_P2_INSTQUEUE_REG_6__0_ <= n6256;
    P1_P2_INSTQUEUE_REG_5__7_ <= n6261;
    P1_P2_INSTQUEUE_REG_5__6_ <= n6266;
    P1_P2_INSTQUEUE_REG_5__5_ <= n6271;
    P1_P2_INSTQUEUE_REG_5__4_ <= n6276;
    P1_P2_INSTQUEUE_REG_5__3_ <= n6281;
    P1_P2_INSTQUEUE_REG_5__2_ <= n6286;
    P1_P2_INSTQUEUE_REG_5__1_ <= n6291;
    P1_P2_INSTQUEUE_REG_5__0_ <= n6296;
    P1_P2_INSTQUEUE_REG_4__7_ <= n6301;
    P1_P2_INSTQUEUE_REG_4__6_ <= n6306;
    P1_P2_INSTQUEUE_REG_4__5_ <= n6311;
    P1_P2_INSTQUEUE_REG_4__4_ <= n6316;
    P1_P2_INSTQUEUE_REG_4__3_ <= n6321;
    P1_P2_INSTQUEUE_REG_4__2_ <= n6326;
    P1_P2_INSTQUEUE_REG_4__1_ <= n6331;
    P1_P2_INSTQUEUE_REG_4__0_ <= n6336;
    P1_P2_INSTQUEUE_REG_3__7_ <= n6341;
    P1_P2_INSTQUEUE_REG_3__6_ <= n6346;
    P1_P2_INSTQUEUE_REG_3__5_ <= n6351;
    P1_P2_INSTQUEUE_REG_3__4_ <= n6356;
    P1_P2_INSTQUEUE_REG_3__3_ <= n6361;
    P1_P2_INSTQUEUE_REG_3__2_ <= n6366;
    P1_P2_INSTQUEUE_REG_3__1_ <= n6371;
    P1_P2_INSTQUEUE_REG_3__0_ <= n6376;
    P1_P2_INSTQUEUE_REG_2__7_ <= n6381;
    P1_P2_INSTQUEUE_REG_2__6_ <= n6386;
    P1_P2_INSTQUEUE_REG_2__5_ <= n6391;
    P1_P2_INSTQUEUE_REG_2__4_ <= n6396;
    P1_P2_INSTQUEUE_REG_2__3_ <= n6401;
    P1_P2_INSTQUEUE_REG_2__2_ <= n6406;
    P1_P2_INSTQUEUE_REG_2__1_ <= n6411;
    P1_P2_INSTQUEUE_REG_2__0_ <= n6416;
    P1_P2_INSTQUEUE_REG_1__7_ <= n6421;
    P1_P2_INSTQUEUE_REG_1__6_ <= n6426;
    P1_P2_INSTQUEUE_REG_1__5_ <= n6431;
    P1_P2_INSTQUEUE_REG_1__4_ <= n6436;
    P1_P2_INSTQUEUE_REG_1__3_ <= n6441;
    P1_P2_INSTQUEUE_REG_1__2_ <= n6446;
    P1_P2_INSTQUEUE_REG_1__1_ <= n6451;
    P1_P2_INSTQUEUE_REG_1__0_ <= n6456;
    P1_P2_INSTQUEUE_REG_0__7_ <= n6461;
    P1_P2_INSTQUEUE_REG_0__6_ <= n6466;
    P1_P2_INSTQUEUE_REG_0__5_ <= n6471;
    P1_P2_INSTQUEUE_REG_0__4_ <= n6476;
    P1_P2_INSTQUEUE_REG_0__3_ <= n6481;
    P1_P2_INSTQUEUE_REG_0__2_ <= n6486;
    P1_P2_INSTQUEUE_REG_0__1_ <= n6491;
    P1_P2_INSTQUEUE_REG_0__0_ <= n6496;
    P1_P2_INSTQUEUERD_ADDR_REG_4_ <= n6501;
    P1_P2_INSTQUEUERD_ADDR_REG_3_ <= n6506;
    P1_P2_INSTQUEUERD_ADDR_REG_2_ <= n6511;
    P1_P2_INSTQUEUERD_ADDR_REG_1_ <= n6516;
    P1_P2_INSTQUEUERD_ADDR_REG_0_ <= n6521;
    P1_P2_INSTQUEUEWR_ADDR_REG_4_ <= n6526;
    P1_P2_INSTQUEUEWR_ADDR_REG_3_ <= n6531;
    P1_P2_INSTQUEUEWR_ADDR_REG_2_ <= n6536;
    P1_P2_INSTQUEUEWR_ADDR_REG_1_ <= n6541;
    P1_P2_INSTQUEUEWR_ADDR_REG_0_ <= n6546;
    P1_P2_INSTADDRPOINTER_REG_0_ <= n6551;
    P1_P2_INSTADDRPOINTER_REG_1_ <= n6556;
    P1_P2_INSTADDRPOINTER_REG_2_ <= n6561;
    P1_P2_INSTADDRPOINTER_REG_3_ <= n6566;
    P1_P2_INSTADDRPOINTER_REG_4_ <= n6571;
    P1_P2_INSTADDRPOINTER_REG_5_ <= n6576;
    P1_P2_INSTADDRPOINTER_REG_6_ <= n6581;
    P1_P2_INSTADDRPOINTER_REG_7_ <= n6586;
    P1_P2_INSTADDRPOINTER_REG_8_ <= n6591;
    P1_P2_INSTADDRPOINTER_REG_9_ <= n6596;
    P1_P2_INSTADDRPOINTER_REG_10_ <= n6601;
    P1_P2_INSTADDRPOINTER_REG_11_ <= n6606;
    P1_P2_INSTADDRPOINTER_REG_12_ <= n6611;
    P1_P2_INSTADDRPOINTER_REG_13_ <= n6616;
    P1_P2_INSTADDRPOINTER_REG_14_ <= n6621;
    P1_P2_INSTADDRPOINTER_REG_15_ <= n6626;
    P1_P2_INSTADDRPOINTER_REG_16_ <= n6631;
    P1_P2_INSTADDRPOINTER_REG_17_ <= n6636;
    P1_P2_INSTADDRPOINTER_REG_18_ <= n6641;
    P1_P2_INSTADDRPOINTER_REG_19_ <= n6646;
    P1_P2_INSTADDRPOINTER_REG_20_ <= n6651;
    P1_P2_INSTADDRPOINTER_REG_21_ <= n6656;
    P1_P2_INSTADDRPOINTER_REG_22_ <= n6661;
    P1_P2_INSTADDRPOINTER_REG_23_ <= n6666;
    P1_P2_INSTADDRPOINTER_REG_24_ <= n6671;
    P1_P2_INSTADDRPOINTER_REG_25_ <= n6676;
    P1_P2_INSTADDRPOINTER_REG_26_ <= n6681;
    P1_P2_INSTADDRPOINTER_REG_27_ <= n6686;
    P1_P2_INSTADDRPOINTER_REG_28_ <= n6691;
    P1_P2_INSTADDRPOINTER_REG_29_ <= n6696;
    P1_P2_INSTADDRPOINTER_REG_30_ <= n6701;
    P1_P2_INSTADDRPOINTER_REG_31_ <= n6706;
    P1_P2_PHYADDRPOINTER_REG_0_ <= n6711;
    P1_P2_PHYADDRPOINTER_REG_1_ <= n6716;
    P1_P2_PHYADDRPOINTER_REG_2_ <= n6721;
    P1_P2_PHYADDRPOINTER_REG_3_ <= n6726;
    P1_P2_PHYADDRPOINTER_REG_4_ <= n6731;
    P1_P2_PHYADDRPOINTER_REG_5_ <= n6736;
    P1_P2_PHYADDRPOINTER_REG_6_ <= n6741;
    P1_P2_PHYADDRPOINTER_REG_7_ <= n6746;
    P1_P2_PHYADDRPOINTER_REG_8_ <= n6751;
    P1_P2_PHYADDRPOINTER_REG_9_ <= n6756;
    P1_P2_PHYADDRPOINTER_REG_10_ <= n6761;
    P1_P2_PHYADDRPOINTER_REG_11_ <= n6766;
    P1_P2_PHYADDRPOINTER_REG_12_ <= n6771;
    P1_P2_PHYADDRPOINTER_REG_13_ <= n6776;
    P1_P2_PHYADDRPOINTER_REG_14_ <= n6781;
    P1_P2_PHYADDRPOINTER_REG_15_ <= n6786;
    P1_P2_PHYADDRPOINTER_REG_16_ <= n6791;
    P1_P2_PHYADDRPOINTER_REG_17_ <= n6796;
    P1_P2_PHYADDRPOINTER_REG_18_ <= n6801;
    P1_P2_PHYADDRPOINTER_REG_19_ <= n6806;
    P1_P2_PHYADDRPOINTER_REG_20_ <= n6811;
    P1_P2_PHYADDRPOINTER_REG_21_ <= n6816;
    P1_P2_PHYADDRPOINTER_REG_22_ <= n6821;
    P1_P2_PHYADDRPOINTER_REG_23_ <= n6826;
    P1_P2_PHYADDRPOINTER_REG_24_ <= n6831;
    P1_P2_PHYADDRPOINTER_REG_25_ <= n6836;
    P1_P2_PHYADDRPOINTER_REG_26_ <= n6841;
    P1_P2_PHYADDRPOINTER_REG_27_ <= n6846;
    P1_P2_PHYADDRPOINTER_REG_28_ <= n6851;
    P1_P2_PHYADDRPOINTER_REG_29_ <= n6856;
    P1_P2_PHYADDRPOINTER_REG_30_ <= n6861;
    P1_P2_PHYADDRPOINTER_REG_31_ <= n6866;
    P1_P2_LWORD_REG_15_ <= n6871;
    P1_P2_LWORD_REG_14_ <= n6876;
    P1_P2_LWORD_REG_13_ <= n6881;
    P1_P2_LWORD_REG_12_ <= n6886;
    P1_P2_LWORD_REG_11_ <= n6891;
    P1_P2_LWORD_REG_10_ <= n6896;
    P1_P2_LWORD_REG_9_ <= n6901;
    P1_P2_LWORD_REG_8_ <= n6906;
    P1_P2_LWORD_REG_7_ <= n6911;
    P1_P2_LWORD_REG_6_ <= n6916;
    P1_P2_LWORD_REG_5_ <= n6921;
    P1_P2_LWORD_REG_4_ <= n6926;
    P1_P2_LWORD_REG_3_ <= n6931;
    P1_P2_LWORD_REG_2_ <= n6936;
    P1_P2_LWORD_REG_1_ <= n6941;
    P1_P2_LWORD_REG_0_ <= n6946;
    P1_P2_UWORD_REG_14_ <= n6951;
    P1_P2_UWORD_REG_13_ <= n6956;
    P1_P2_UWORD_REG_12_ <= n6961;
    P1_P2_UWORD_REG_11_ <= n6966;
    P1_P2_UWORD_REG_10_ <= n6971;
    P1_P2_UWORD_REG_9_ <= n6976;
    P1_P2_UWORD_REG_8_ <= n6981;
    P1_P2_UWORD_REG_7_ <= n6986;
    P1_P2_UWORD_REG_6_ <= n6991;
    P1_P2_UWORD_REG_5_ <= n6996;
    P1_P2_UWORD_REG_4_ <= n7001;
    P1_P2_UWORD_REG_3_ <= n7006;
    P1_P2_UWORD_REG_2_ <= n7011;
    P1_P2_UWORD_REG_1_ <= n7016;
    P1_P2_UWORD_REG_0_ <= n7021;
    P1_P2_DATAO_REG_0_ <= n7026;
    P1_P2_DATAO_REG_1_ <= n7031;
    P1_P2_DATAO_REG_2_ <= n7036;
    P1_P2_DATAO_REG_3_ <= n7041;
    P1_P2_DATAO_REG_4_ <= n7046;
    P1_P2_DATAO_REG_5_ <= n7051;
    P1_P2_DATAO_REG_6_ <= n7056;
    P1_P2_DATAO_REG_7_ <= n7061;
    P1_P2_DATAO_REG_8_ <= n7066;
    P1_P2_DATAO_REG_9_ <= n7071;
    P1_P2_DATAO_REG_10_ <= n7076;
    P1_P2_DATAO_REG_11_ <= n7081;
    P1_P2_DATAO_REG_12_ <= n7086;
    P1_P2_DATAO_REG_13_ <= n7091;
    P1_P2_DATAO_REG_14_ <= n7096;
    P1_P2_DATAO_REG_15_ <= n7101;
    P1_P2_DATAO_REG_16_ <= n7106;
    P1_P2_DATAO_REG_17_ <= n7111;
    P1_P2_DATAO_REG_18_ <= n7116;
    P1_P2_DATAO_REG_19_ <= n7121;
    P1_P2_DATAO_REG_20_ <= n7126;
    P1_P2_DATAO_REG_21_ <= n7131;
    P1_P2_DATAO_REG_22_ <= n7136;
    P1_P2_DATAO_REG_23_ <= n7141;
    P1_P2_DATAO_REG_24_ <= n7146;
    P1_P2_DATAO_REG_25_ <= n7151;
    P1_P2_DATAO_REG_26_ <= n7156;
    P1_P2_DATAO_REG_27_ <= n7161;
    P1_P2_DATAO_REG_28_ <= n7166;
    P1_P2_DATAO_REG_29_ <= n7171;
    P1_P2_DATAO_REG_30_ <= n7176;
    P1_P2_DATAO_REG_31_ <= n7181;
    P1_P2_EAX_REG_0_ <= n7186;
    P1_P2_EAX_REG_1_ <= n7191;
    P1_P2_EAX_REG_2_ <= n7196;
    P1_P2_EAX_REG_3_ <= n7201;
    P1_P2_EAX_REG_4_ <= n7206;
    P1_P2_EAX_REG_5_ <= n7211;
    P1_P2_EAX_REG_6_ <= n7216;
    P1_P2_EAX_REG_7_ <= n7221;
    P1_P2_EAX_REG_8_ <= n7226;
    P1_P2_EAX_REG_9_ <= n7231;
    P1_P2_EAX_REG_10_ <= n7236;
    P1_P2_EAX_REG_11_ <= n7241;
    P1_P2_EAX_REG_12_ <= n7246;
    P1_P2_EAX_REG_13_ <= n7251;
    P1_P2_EAX_REG_14_ <= n7256;
    P1_P2_EAX_REG_15_ <= n7261;
    P1_P2_EAX_REG_16_ <= n7266;
    P1_P2_EAX_REG_17_ <= n7271;
    P1_P2_EAX_REG_18_ <= n7276;
    P1_P2_EAX_REG_19_ <= n7281;
    P1_P2_EAX_REG_20_ <= n7286;
    P1_P2_EAX_REG_21_ <= n7291;
    P1_P2_EAX_REG_22_ <= n7296;
    P1_P2_EAX_REG_23_ <= n7301;
    P1_P2_EAX_REG_24_ <= n7306;
    P1_P2_EAX_REG_25_ <= n7311;
    P1_P2_EAX_REG_26_ <= n7316;
    P1_P2_EAX_REG_27_ <= n7321;
    P1_P2_EAX_REG_28_ <= n7326;
    P1_P2_EAX_REG_29_ <= n7331;
    P1_P2_EAX_REG_30_ <= n7336;
    P1_P2_EAX_REG_31_ <= n7341;
    P1_P2_EBX_REG_0_ <= n7346;
    P1_P2_EBX_REG_1_ <= n7351;
    P1_P2_EBX_REG_2_ <= n7356;
    P1_P2_EBX_REG_3_ <= n7361;
    P1_P2_EBX_REG_4_ <= n7366;
    P1_P2_EBX_REG_5_ <= n7371;
    P1_P2_EBX_REG_6_ <= n7376;
    P1_P2_EBX_REG_7_ <= n7381;
    P1_P2_EBX_REG_8_ <= n7386;
    P1_P2_EBX_REG_9_ <= n7391;
    P1_P2_EBX_REG_10_ <= n7396;
    P1_P2_EBX_REG_11_ <= n7401;
    P1_P2_EBX_REG_12_ <= n7406;
    P1_P2_EBX_REG_13_ <= n7411;
    P1_P2_EBX_REG_14_ <= n7416;
    P1_P2_EBX_REG_15_ <= n7421;
    P1_P2_EBX_REG_16_ <= n7426;
    P1_P2_EBX_REG_17_ <= n7431;
    P1_P2_EBX_REG_18_ <= n7436;
    P1_P2_EBX_REG_19_ <= n7441;
    P1_P2_EBX_REG_20_ <= n7446;
    P1_P2_EBX_REG_21_ <= n7451;
    P1_P2_EBX_REG_22_ <= n7456;
    P1_P2_EBX_REG_23_ <= n7461;
    P1_P2_EBX_REG_24_ <= n7466;
    P1_P2_EBX_REG_25_ <= n7471;
    P1_P2_EBX_REG_26_ <= n7476;
    P1_P2_EBX_REG_27_ <= n7481;
    P1_P2_EBX_REG_28_ <= n7486;
    P1_P2_EBX_REG_29_ <= n7491;
    P1_P2_EBX_REG_30_ <= n7496;
    P1_P2_EBX_REG_31_ <= n7501;
    P1_P2_REIP_REG_0_ <= n7506;
    P1_P2_REIP_REG_1_ <= n7511;
    P1_P2_REIP_REG_2_ <= n7516;
    P1_P2_REIP_REG_3_ <= n7521;
    P1_P2_REIP_REG_4_ <= n7526;
    P1_P2_REIP_REG_5_ <= n7531;
    P1_P2_REIP_REG_6_ <= n7536;
    P1_P2_REIP_REG_7_ <= n7541;
    P1_P2_REIP_REG_8_ <= n7546;
    P1_P2_REIP_REG_9_ <= n7551;
    P1_P2_REIP_REG_10_ <= n7556;
    P1_P2_REIP_REG_11_ <= n7561;
    P1_P2_REIP_REG_12_ <= n7566;
    P1_P2_REIP_REG_13_ <= n7571;
    P1_P2_REIP_REG_14_ <= n7576;
    P1_P2_REIP_REG_15_ <= n7581;
    P1_P2_REIP_REG_16_ <= n7586;
    P1_P2_REIP_REG_17_ <= n7591;
    P1_P2_REIP_REG_18_ <= n7596;
    P1_P2_REIP_REG_19_ <= n7601;
    P1_P2_REIP_REG_20_ <= n7606;
    P1_P2_REIP_REG_21_ <= n7611;
    P1_P2_REIP_REG_22_ <= n7616;
    P1_P2_REIP_REG_23_ <= n7621;
    P1_P2_REIP_REG_24_ <= n7626;
    P1_P2_REIP_REG_25_ <= n7631;
    P1_P2_REIP_REG_26_ <= n7636;
    P1_P2_REIP_REG_27_ <= n7641;
    P1_P2_REIP_REG_28_ <= n7646;
    P1_P2_REIP_REG_29_ <= n7651;
    P1_P2_REIP_REG_30_ <= n7656;
    P1_P2_REIP_REG_31_ <= n7661;
    P1_P2_BYTEENABLE_REG_3_ <= n7666;
    P1_P2_BYTEENABLE_REG_2_ <= n7671;
    P1_P2_BYTEENABLE_REG_1_ <= n7676;
    P1_P2_BYTEENABLE_REG_0_ <= n7681;
    P1_P2_W_R_N_REG <= n7686;
    P1_P2_FLUSH_REG <= n7691;
    P1_P2_MORE_REG <= n7696;
    P1_P2_STATEBS16_REG <= n7701;
    P1_P2_REQUESTPENDING_REG <= n7706;
    P1_P2_D_C_N_REG <= n7711;
    P1_P2_M_IO_N_REG <= n7716;
    P1_P2_CODEFETCH_REG <= n7721;
    P1_P2_ADS_N_REG <= n7726;
    P1_P2_READREQUEST_REG <= n7731;
    P1_P2_MEMORYFETCH_REG <= n7736;
    P1_P1_BE_N_REG_3_ <= n7741;
    P1_P1_BE_N_REG_2_ <= n7746;
    P1_P1_BE_N_REG_1_ <= n7751;
    P1_P1_BE_N_REG_0_ <= n7756;
    P1_P1_ADDRESS_REG_29_ <= n7761;
    P1_P1_ADDRESS_REG_28_ <= n7766;
    P1_P1_ADDRESS_REG_27_ <= n7771;
    P1_P1_ADDRESS_REG_26_ <= n7776;
    P1_P1_ADDRESS_REG_25_ <= n7781;
    P1_P1_ADDRESS_REG_24_ <= n7786;
    P1_P1_ADDRESS_REG_23_ <= n7791;
    P1_P1_ADDRESS_REG_22_ <= n7796;
    P1_P1_ADDRESS_REG_21_ <= n7801;
    P1_P1_ADDRESS_REG_20_ <= n7806;
    P1_P1_ADDRESS_REG_19_ <= n7811;
    P1_P1_ADDRESS_REG_18_ <= n7816;
    P1_P1_ADDRESS_REG_17_ <= n7821;
    P1_P1_ADDRESS_REG_16_ <= n7826;
    P1_P1_ADDRESS_REG_15_ <= n7831;
    P1_P1_ADDRESS_REG_14_ <= n7836;
    P1_P1_ADDRESS_REG_13_ <= n7841;
    P1_P1_ADDRESS_REG_12_ <= n7846;
    P1_P1_ADDRESS_REG_11_ <= n7851;
    P1_P1_ADDRESS_REG_10_ <= n7856;
    P1_P1_ADDRESS_REG_9_ <= n7861;
    P1_P1_ADDRESS_REG_8_ <= n7866;
    P1_P1_ADDRESS_REG_7_ <= n7871;
    P1_P1_ADDRESS_REG_6_ <= n7876;
    P1_P1_ADDRESS_REG_5_ <= n7881;
    P1_P1_ADDRESS_REG_4_ <= n7886;
    P1_P1_ADDRESS_REG_3_ <= n7891;
    P1_P1_ADDRESS_REG_2_ <= n7896;
    P1_P1_ADDRESS_REG_1_ <= n7901;
    P1_P1_ADDRESS_REG_0_ <= n7906;
    P1_P1_STATE_REG_2_ <= n7911;
    P1_P1_STATE_REG_1_ <= n7916;
    P1_P1_STATE_REG_0_ <= n7921;
    P1_P1_DATAWIDTH_REG_0_ <= n7926;
    P1_P1_DATAWIDTH_REG_1_ <= n7931;
    P1_P1_DATAWIDTH_REG_2_ <= n7936;
    P1_P1_DATAWIDTH_REG_3_ <= n7941;
    P1_P1_DATAWIDTH_REG_4_ <= n7946;
    P1_P1_DATAWIDTH_REG_5_ <= n7951;
    P1_P1_DATAWIDTH_REG_6_ <= n7956;
    P1_P1_DATAWIDTH_REG_7_ <= n7961;
    P1_P1_DATAWIDTH_REG_8_ <= n7966;
    P1_P1_DATAWIDTH_REG_9_ <= n7971;
    P1_P1_DATAWIDTH_REG_10_ <= n7976;
    P1_P1_DATAWIDTH_REG_11_ <= n7981;
    P1_P1_DATAWIDTH_REG_12_ <= n7986;
    P1_P1_DATAWIDTH_REG_13_ <= n7991;
    P1_P1_DATAWIDTH_REG_14_ <= n7996;
    P1_P1_DATAWIDTH_REG_15_ <= n8001;
    P1_P1_DATAWIDTH_REG_16_ <= n8006;
    P1_P1_DATAWIDTH_REG_17_ <= n8011;
    P1_P1_DATAWIDTH_REG_18_ <= n8016;
    P1_P1_DATAWIDTH_REG_19_ <= n8021;
    P1_P1_DATAWIDTH_REG_20_ <= n8026;
    P1_P1_DATAWIDTH_REG_21_ <= n8031;
    P1_P1_DATAWIDTH_REG_22_ <= n8036;
    P1_P1_DATAWIDTH_REG_23_ <= n8041;
    P1_P1_DATAWIDTH_REG_24_ <= n8046;
    P1_P1_DATAWIDTH_REG_25_ <= n8051;
    P1_P1_DATAWIDTH_REG_26_ <= n8056;
    P1_P1_DATAWIDTH_REG_27_ <= n8061;
    P1_P1_DATAWIDTH_REG_28_ <= n8066;
    P1_P1_DATAWIDTH_REG_29_ <= n8071;
    P1_P1_DATAWIDTH_REG_30_ <= n8076;
    P1_P1_DATAWIDTH_REG_31_ <= n8081;
    P1_P1_STATE2_REG_3_ <= n8086;
    P1_P1_STATE2_REG_2_ <= n8091;
    P1_P1_STATE2_REG_1_ <= n8096;
    P1_P1_STATE2_REG_0_ <= n8101;
    P1_P1_INSTQUEUE_REG_15__7_ <= n8106;
    P1_P1_INSTQUEUE_REG_15__6_ <= n8111;
    P1_P1_INSTQUEUE_REG_15__5_ <= n8116;
    P1_P1_INSTQUEUE_REG_15__4_ <= n8121;
    P1_P1_INSTQUEUE_REG_15__3_ <= n8126;
    P1_P1_INSTQUEUE_REG_15__2_ <= n8131;
    P1_P1_INSTQUEUE_REG_15__1_ <= n8136;
    P1_P1_INSTQUEUE_REG_15__0_ <= n8141;
    P1_P1_INSTQUEUE_REG_14__7_ <= n8146;
    P1_P1_INSTQUEUE_REG_14__6_ <= n8151;
    P1_P1_INSTQUEUE_REG_14__5_ <= n8156;
    P1_P1_INSTQUEUE_REG_14__4_ <= n8161;
    P1_P1_INSTQUEUE_REG_14__3_ <= n8166;
    P1_P1_INSTQUEUE_REG_14__2_ <= n8171;
    P1_P1_INSTQUEUE_REG_14__1_ <= n8176;
    P1_P1_INSTQUEUE_REG_14__0_ <= n8181;
    P1_P1_INSTQUEUE_REG_13__7_ <= n8186;
    P1_P1_INSTQUEUE_REG_13__6_ <= n8191;
    P1_P1_INSTQUEUE_REG_13__5_ <= n8196;
    P1_P1_INSTQUEUE_REG_13__4_ <= n8201;
    P1_P1_INSTQUEUE_REG_13__3_ <= n8206;
    P1_P1_INSTQUEUE_REG_13__2_ <= n8211;
    P1_P1_INSTQUEUE_REG_13__1_ <= n8216;
    P1_P1_INSTQUEUE_REG_13__0_ <= n8221;
    P1_P1_INSTQUEUE_REG_12__7_ <= n8226;
    P1_P1_INSTQUEUE_REG_12__6_ <= n8231;
    P1_P1_INSTQUEUE_REG_12__5_ <= n8236;
    P1_P1_INSTQUEUE_REG_12__4_ <= n8241;
    P1_P1_INSTQUEUE_REG_12__3_ <= n8246;
    P1_P1_INSTQUEUE_REG_12__2_ <= n8251;
    P1_P1_INSTQUEUE_REG_12__1_ <= n8256;
    P1_P1_INSTQUEUE_REG_12__0_ <= n8261;
    P1_P1_INSTQUEUE_REG_11__7_ <= n8266;
    P1_P1_INSTQUEUE_REG_11__6_ <= n8271;
    P1_P1_INSTQUEUE_REG_11__5_ <= n8276;
    P1_P1_INSTQUEUE_REG_11__4_ <= n8281;
    P1_P1_INSTQUEUE_REG_11__3_ <= n8286;
    P1_P1_INSTQUEUE_REG_11__2_ <= n8291;
    P1_P1_INSTQUEUE_REG_11__1_ <= n8296;
    P1_P1_INSTQUEUE_REG_11__0_ <= n8301;
    P1_P1_INSTQUEUE_REG_10__7_ <= n8306;
    P1_P1_INSTQUEUE_REG_10__6_ <= n8311;
    P1_P1_INSTQUEUE_REG_10__5_ <= n8316;
    P1_P1_INSTQUEUE_REG_10__4_ <= n8321;
    P1_P1_INSTQUEUE_REG_10__3_ <= n8326;
    P1_P1_INSTQUEUE_REG_10__2_ <= n8331;
    P1_P1_INSTQUEUE_REG_10__1_ <= n8336;
    P1_P1_INSTQUEUE_REG_10__0_ <= n8341;
    P1_P1_INSTQUEUE_REG_9__7_ <= n8346;
    P1_P1_INSTQUEUE_REG_9__6_ <= n8351;
    P1_P1_INSTQUEUE_REG_9__5_ <= n8356;
    P1_P1_INSTQUEUE_REG_9__4_ <= n8361;
    P1_P1_INSTQUEUE_REG_9__3_ <= n8366;
    P1_P1_INSTQUEUE_REG_9__2_ <= n8371;
    P1_P1_INSTQUEUE_REG_9__1_ <= n8376;
    P1_P1_INSTQUEUE_REG_9__0_ <= n8381;
    P1_P1_INSTQUEUE_REG_8__7_ <= n8386;
    P1_P1_INSTQUEUE_REG_8__6_ <= n8391;
    P1_P1_INSTQUEUE_REG_8__5_ <= n8396;
    P1_P1_INSTQUEUE_REG_8__4_ <= n8401;
    P1_P1_INSTQUEUE_REG_8__3_ <= n8406;
    P1_P1_INSTQUEUE_REG_8__2_ <= n8411;
    P1_P1_INSTQUEUE_REG_8__1_ <= n8416;
    P1_P1_INSTQUEUE_REG_8__0_ <= n8421;
    P1_P1_INSTQUEUE_REG_7__7_ <= n8426;
    P1_P1_INSTQUEUE_REG_7__6_ <= n8431;
    P1_P1_INSTQUEUE_REG_7__5_ <= n8436;
    P1_P1_INSTQUEUE_REG_7__4_ <= n8441;
    P1_P1_INSTQUEUE_REG_7__3_ <= n8446;
    P1_P1_INSTQUEUE_REG_7__2_ <= n8451;
    P1_P1_INSTQUEUE_REG_7__1_ <= n8456;
    P1_P1_INSTQUEUE_REG_7__0_ <= n8461;
    P1_P1_INSTQUEUE_REG_6__7_ <= n8466;
    P1_P1_INSTQUEUE_REG_6__6_ <= n8471;
    P1_P1_INSTQUEUE_REG_6__5_ <= n8476;
    P1_P1_INSTQUEUE_REG_6__4_ <= n8481;
    P1_P1_INSTQUEUE_REG_6__3_ <= n8486;
    P1_P1_INSTQUEUE_REG_6__2_ <= n8491;
    P1_P1_INSTQUEUE_REG_6__1_ <= n8496;
    P1_P1_INSTQUEUE_REG_6__0_ <= n8501;
    P1_P1_INSTQUEUE_REG_5__7_ <= n8506;
    P1_P1_INSTQUEUE_REG_5__6_ <= n8511;
    P1_P1_INSTQUEUE_REG_5__5_ <= n8516;
    P1_P1_INSTQUEUE_REG_5__4_ <= n8521;
    P1_P1_INSTQUEUE_REG_5__3_ <= n8526;
    P1_P1_INSTQUEUE_REG_5__2_ <= n8531;
    P1_P1_INSTQUEUE_REG_5__1_ <= n8536;
    P1_P1_INSTQUEUE_REG_5__0_ <= n8541;
    P1_P1_INSTQUEUE_REG_4__7_ <= n8546;
    P1_P1_INSTQUEUE_REG_4__6_ <= n8551;
    P1_P1_INSTQUEUE_REG_4__5_ <= n8556;
    P1_P1_INSTQUEUE_REG_4__4_ <= n8561;
    P1_P1_INSTQUEUE_REG_4__3_ <= n8566;
    P1_P1_INSTQUEUE_REG_4__2_ <= n8571;
    P1_P1_INSTQUEUE_REG_4__1_ <= n8576;
    P1_P1_INSTQUEUE_REG_4__0_ <= n8581;
    P1_P1_INSTQUEUE_REG_3__7_ <= n8586;
    P1_P1_INSTQUEUE_REG_3__6_ <= n8591;
    P1_P1_INSTQUEUE_REG_3__5_ <= n8596;
    P1_P1_INSTQUEUE_REG_3__4_ <= n8601;
    P1_P1_INSTQUEUE_REG_3__3_ <= n8606;
    P1_P1_INSTQUEUE_REG_3__2_ <= n8611;
    P1_P1_INSTQUEUE_REG_3__1_ <= n8616;
    P1_P1_INSTQUEUE_REG_3__0_ <= n8621;
    P1_P1_INSTQUEUE_REG_2__7_ <= n8626;
    P1_P1_INSTQUEUE_REG_2__6_ <= n8631;
    P1_P1_INSTQUEUE_REG_2__5_ <= n8636;
    P1_P1_INSTQUEUE_REG_2__4_ <= n8641;
    P1_P1_INSTQUEUE_REG_2__3_ <= n8646;
    P1_P1_INSTQUEUE_REG_2__2_ <= n8651;
    P1_P1_INSTQUEUE_REG_2__1_ <= n8656;
    P1_P1_INSTQUEUE_REG_2__0_ <= n8661;
    P1_P1_INSTQUEUE_REG_1__7_ <= n8666;
    P1_P1_INSTQUEUE_REG_1__6_ <= n8671;
    P1_P1_INSTQUEUE_REG_1__5_ <= n8676;
    P1_P1_INSTQUEUE_REG_1__4_ <= n8681;
    P1_P1_INSTQUEUE_REG_1__3_ <= n8686;
    P1_P1_INSTQUEUE_REG_1__2_ <= n8691;
    P1_P1_INSTQUEUE_REG_1__1_ <= n8696;
    P1_P1_INSTQUEUE_REG_1__0_ <= n8701;
    P1_P1_INSTQUEUE_REG_0__7_ <= n8706;
    P1_P1_INSTQUEUE_REG_0__6_ <= n8711;
    P1_P1_INSTQUEUE_REG_0__5_ <= n8716;
    P1_P1_INSTQUEUE_REG_0__4_ <= n8721;
    P1_P1_INSTQUEUE_REG_0__3_ <= n8726;
    P1_P1_INSTQUEUE_REG_0__2_ <= n8731;
    P1_P1_INSTQUEUE_REG_0__1_ <= n8736;
    P1_P1_INSTQUEUE_REG_0__0_ <= n8741;
    P1_P1_INSTQUEUERD_ADDR_REG_4_ <= n8746;
    P1_P1_INSTQUEUERD_ADDR_REG_3_ <= n8751;
    P1_P1_INSTQUEUERD_ADDR_REG_2_ <= n8756;
    P1_P1_INSTQUEUERD_ADDR_REG_1_ <= n8761;
    P1_P1_INSTQUEUERD_ADDR_REG_0_ <= n8766;
    P1_P1_INSTQUEUEWR_ADDR_REG_4_ <= n8771;
    P1_P1_INSTQUEUEWR_ADDR_REG_3_ <= n8776;
    P1_P1_INSTQUEUEWR_ADDR_REG_2_ <= n8781;
    P1_P1_INSTQUEUEWR_ADDR_REG_1_ <= n8786;
    P1_P1_INSTQUEUEWR_ADDR_REG_0_ <= n8791;
    P1_P1_INSTADDRPOINTER_REG_0_ <= n8796;
    P1_P1_INSTADDRPOINTER_REG_1_ <= n8801;
    P1_P1_INSTADDRPOINTER_REG_2_ <= n8806;
    P1_P1_INSTADDRPOINTER_REG_3_ <= n8811;
    P1_P1_INSTADDRPOINTER_REG_4_ <= n8816;
    P1_P1_INSTADDRPOINTER_REG_5_ <= n8821;
    P1_P1_INSTADDRPOINTER_REG_6_ <= n8826;
    P1_P1_INSTADDRPOINTER_REG_7_ <= n8831;
    P1_P1_INSTADDRPOINTER_REG_8_ <= n8836;
    P1_P1_INSTADDRPOINTER_REG_9_ <= n8841;
    P1_P1_INSTADDRPOINTER_REG_10_ <= n8846;
    P1_P1_INSTADDRPOINTER_REG_11_ <= n8851;
    P1_P1_INSTADDRPOINTER_REG_12_ <= n8856;
    P1_P1_INSTADDRPOINTER_REG_13_ <= n8861;
    P1_P1_INSTADDRPOINTER_REG_14_ <= n8866;
    P1_P1_INSTADDRPOINTER_REG_15_ <= n8871;
    P1_P1_INSTADDRPOINTER_REG_16_ <= n8876;
    P1_P1_INSTADDRPOINTER_REG_17_ <= n8881;
    P1_P1_INSTADDRPOINTER_REG_18_ <= n8886;
    P1_P1_INSTADDRPOINTER_REG_19_ <= n8891;
    P1_P1_INSTADDRPOINTER_REG_20_ <= n8896;
    P1_P1_INSTADDRPOINTER_REG_21_ <= n8901;
    P1_P1_INSTADDRPOINTER_REG_22_ <= n8906;
    P1_P1_INSTADDRPOINTER_REG_23_ <= n8911;
    P1_P1_INSTADDRPOINTER_REG_24_ <= n8916;
    P1_P1_INSTADDRPOINTER_REG_25_ <= n8921;
    P1_P1_INSTADDRPOINTER_REG_26_ <= n8926;
    P1_P1_INSTADDRPOINTER_REG_27_ <= n8931;
    P1_P1_INSTADDRPOINTER_REG_28_ <= n8936;
    P1_P1_INSTADDRPOINTER_REG_29_ <= n8941;
    P1_P1_INSTADDRPOINTER_REG_30_ <= n8946;
    P1_P1_INSTADDRPOINTER_REG_31_ <= n8951;
    P1_P1_PHYADDRPOINTER_REG_0_ <= n8956;
    P1_P1_PHYADDRPOINTER_REG_1_ <= n8961;
    P1_P1_PHYADDRPOINTER_REG_2_ <= n8966;
    P1_P1_PHYADDRPOINTER_REG_3_ <= n8971;
    P1_P1_PHYADDRPOINTER_REG_4_ <= n8976;
    P1_P1_PHYADDRPOINTER_REG_5_ <= n8981;
    P1_P1_PHYADDRPOINTER_REG_6_ <= n8986;
    P1_P1_PHYADDRPOINTER_REG_7_ <= n8991;
    P1_P1_PHYADDRPOINTER_REG_8_ <= n8996;
    P1_P1_PHYADDRPOINTER_REG_9_ <= n9001;
    P1_P1_PHYADDRPOINTER_REG_10_ <= n9006;
    P1_P1_PHYADDRPOINTER_REG_11_ <= n9011;
    P1_P1_PHYADDRPOINTER_REG_12_ <= n9016;
    P1_P1_PHYADDRPOINTER_REG_13_ <= n9021;
    P1_P1_PHYADDRPOINTER_REG_14_ <= n9026;
    P1_P1_PHYADDRPOINTER_REG_15_ <= n9031;
    P1_P1_PHYADDRPOINTER_REG_16_ <= n9036;
    P1_P1_PHYADDRPOINTER_REG_17_ <= n9041;
    P1_P1_PHYADDRPOINTER_REG_18_ <= n9046;
    P1_P1_PHYADDRPOINTER_REG_19_ <= n9051;
    P1_P1_PHYADDRPOINTER_REG_20_ <= n9056;
    P1_P1_PHYADDRPOINTER_REG_21_ <= n9061;
    P1_P1_PHYADDRPOINTER_REG_22_ <= n9066;
    P1_P1_PHYADDRPOINTER_REG_23_ <= n9071;
    P1_P1_PHYADDRPOINTER_REG_24_ <= n9076;
    P1_P1_PHYADDRPOINTER_REG_25_ <= n9081;
    P1_P1_PHYADDRPOINTER_REG_26_ <= n9086;
    P1_P1_PHYADDRPOINTER_REG_27_ <= n9091;
    P1_P1_PHYADDRPOINTER_REG_28_ <= n9096;
    P1_P1_PHYADDRPOINTER_REG_29_ <= n9101;
    P1_P1_PHYADDRPOINTER_REG_30_ <= n9106;
    P1_P1_PHYADDRPOINTER_REG_31_ <= n9111;
    P1_P1_LWORD_REG_15_ <= n9116;
    P1_P1_LWORD_REG_14_ <= n9121;
    P1_P1_LWORD_REG_13_ <= n9126;
    P1_P1_LWORD_REG_12_ <= n9131;
    P1_P1_LWORD_REG_11_ <= n9136;
    P1_P1_LWORD_REG_10_ <= n9141;
    P1_P1_LWORD_REG_9_ <= n9146;
    P1_P1_LWORD_REG_8_ <= n9151;
    P1_P1_LWORD_REG_7_ <= n9156;
    P1_P1_LWORD_REG_6_ <= n9161;
    P1_P1_LWORD_REG_5_ <= n9166;
    P1_P1_LWORD_REG_4_ <= n9171;
    P1_P1_LWORD_REG_3_ <= n9176;
    P1_P1_LWORD_REG_2_ <= n9181;
    P1_P1_LWORD_REG_1_ <= n9186;
    P1_P1_LWORD_REG_0_ <= n9191;
    P1_P1_UWORD_REG_14_ <= n9196;
    P1_P1_UWORD_REG_13_ <= n9201;
    P1_P1_UWORD_REG_12_ <= n9206;
    P1_P1_UWORD_REG_11_ <= n9211;
    P1_P1_UWORD_REG_10_ <= n9216;
    P1_P1_UWORD_REG_9_ <= n9221;
    P1_P1_UWORD_REG_8_ <= n9226;
    P1_P1_UWORD_REG_7_ <= n9231;
    P1_P1_UWORD_REG_6_ <= n9236;
    P1_P1_UWORD_REG_5_ <= n9241;
    P1_P1_UWORD_REG_4_ <= n9246;
    P1_P1_UWORD_REG_3_ <= n9251;
    P1_P1_UWORD_REG_2_ <= n9256;
    P1_P1_UWORD_REG_1_ <= n9261;
    P1_P1_UWORD_REG_0_ <= n9266;
    P1_P1_DATAO_REG_0_ <= n9271;
    P1_P1_DATAO_REG_1_ <= n9276;
    P1_P1_DATAO_REG_2_ <= n9281;
    P1_P1_DATAO_REG_3_ <= n9286;
    P1_P1_DATAO_REG_4_ <= n9291;
    P1_P1_DATAO_REG_5_ <= n9296;
    P1_P1_DATAO_REG_6_ <= n9301;
    P1_P1_DATAO_REG_7_ <= n9306;
    P1_P1_DATAO_REG_8_ <= n9311;
    P1_P1_DATAO_REG_9_ <= n9316;
    P1_P1_DATAO_REG_10_ <= n9321;
    P1_P1_DATAO_REG_11_ <= n9326;
    P1_P1_DATAO_REG_12_ <= n9331;
    P1_P1_DATAO_REG_13_ <= n9336;
    P1_P1_DATAO_REG_14_ <= n9341;
    P1_P1_DATAO_REG_15_ <= n9346;
    P1_P1_DATAO_REG_16_ <= n9351;
    P1_P1_DATAO_REG_17_ <= n9356;
    P1_P1_DATAO_REG_18_ <= n9361;
    P1_P1_DATAO_REG_19_ <= n9366;
    P1_P1_DATAO_REG_20_ <= n9371;
    P1_P1_DATAO_REG_21_ <= n9376;
    P1_P1_DATAO_REG_22_ <= n9381;
    P1_P1_DATAO_REG_23_ <= n9386;
    P1_P1_DATAO_REG_24_ <= n9391;
    P1_P1_DATAO_REG_25_ <= n9396;
    P1_P1_DATAO_REG_26_ <= n9401;
    P1_P1_DATAO_REG_27_ <= n9406;
    P1_P1_DATAO_REG_28_ <= n9411;
    P1_P1_DATAO_REG_29_ <= n9416;
    P1_P1_DATAO_REG_30_ <= n9421;
    P1_P1_DATAO_REG_31_ <= n9426;
    P1_P1_EAX_REG_0_ <= n9431;
    P1_P1_EAX_REG_1_ <= n9436;
    P1_P1_EAX_REG_2_ <= n9441;
    P1_P1_EAX_REG_3_ <= n9446;
    P1_P1_EAX_REG_4_ <= n9451;
    P1_P1_EAX_REG_5_ <= n9456;
    P1_P1_EAX_REG_6_ <= n9461;
    P1_P1_EAX_REG_7_ <= n9466;
    P1_P1_EAX_REG_8_ <= n9471;
    P1_P1_EAX_REG_9_ <= n9476;
    P1_P1_EAX_REG_10_ <= n9481;
    P1_P1_EAX_REG_11_ <= n9486;
    P1_P1_EAX_REG_12_ <= n9491;
    P1_P1_EAX_REG_13_ <= n9496;
    P1_P1_EAX_REG_14_ <= n9501;
    P1_P1_EAX_REG_15_ <= n9506;
    P1_P1_EAX_REG_16_ <= n9511;
    P1_P1_EAX_REG_17_ <= n9516;
    P1_P1_EAX_REG_18_ <= n9521;
    P1_P1_EAX_REG_19_ <= n9526;
    P1_P1_EAX_REG_20_ <= n9531;
    P1_P1_EAX_REG_21_ <= n9536;
    P1_P1_EAX_REG_22_ <= n9541;
    P1_P1_EAX_REG_23_ <= n9546;
    P1_P1_EAX_REG_24_ <= n9551;
    P1_P1_EAX_REG_25_ <= n9556;
    P1_P1_EAX_REG_26_ <= n9561;
    P1_P1_EAX_REG_27_ <= n9566;
    P1_P1_EAX_REG_28_ <= n9571;
    P1_P1_EAX_REG_29_ <= n9576;
    P1_P1_EAX_REG_30_ <= n9581;
    P1_P1_EAX_REG_31_ <= n9586;
    P1_P1_EBX_REG_0_ <= n9591;
    P1_P1_EBX_REG_1_ <= n9596;
    P1_P1_EBX_REG_2_ <= n9601;
    P1_P1_EBX_REG_3_ <= n9606;
    P1_P1_EBX_REG_4_ <= n9611;
    P1_P1_EBX_REG_5_ <= n9616;
    P1_P1_EBX_REG_6_ <= n9621;
    P1_P1_EBX_REG_7_ <= n9626;
    P1_P1_EBX_REG_8_ <= n9631;
    P1_P1_EBX_REG_9_ <= n9636;
    P1_P1_EBX_REG_10_ <= n9641;
    P1_P1_EBX_REG_11_ <= n9646;
    P1_P1_EBX_REG_12_ <= n9651;
    P1_P1_EBX_REG_13_ <= n9656;
    P1_P1_EBX_REG_14_ <= n9661;
    P1_P1_EBX_REG_15_ <= n9666;
    P1_P1_EBX_REG_16_ <= n9671;
    P1_P1_EBX_REG_17_ <= n9676;
    P1_P1_EBX_REG_18_ <= n9681;
    P1_P1_EBX_REG_19_ <= n9686;
    P1_P1_EBX_REG_20_ <= n9691;
    P1_P1_EBX_REG_21_ <= n9696;
    P1_P1_EBX_REG_22_ <= n9701;
    P1_P1_EBX_REG_23_ <= n9706;
    P1_P1_EBX_REG_24_ <= n9711;
    P1_P1_EBX_REG_25_ <= n9716;
    P1_P1_EBX_REG_26_ <= n9721;
    P1_P1_EBX_REG_27_ <= n9726;
    P1_P1_EBX_REG_28_ <= n9731;
    P1_P1_EBX_REG_29_ <= n9736;
    P1_P1_EBX_REG_30_ <= n9741;
    P1_P1_EBX_REG_31_ <= n9746;
    P1_P1_REIP_REG_0_ <= n9751;
    P1_P1_REIP_REG_1_ <= n9756;
    P1_P1_REIP_REG_2_ <= n9761;
    P1_P1_REIP_REG_3_ <= n9766;
    P1_P1_REIP_REG_4_ <= n9771;
    P1_P1_REIP_REG_5_ <= n9776;
    P1_P1_REIP_REG_6_ <= n9781;
    P1_P1_REIP_REG_7_ <= n9786;
    P1_P1_REIP_REG_8_ <= n9791;
    P1_P1_REIP_REG_9_ <= n9796;
    P1_P1_REIP_REG_10_ <= n9801;
    P1_P1_REIP_REG_11_ <= n9806;
    P1_P1_REIP_REG_12_ <= n9811;
    P1_P1_REIP_REG_13_ <= n9816;
    P1_P1_REIP_REG_14_ <= n9821;
    P1_P1_REIP_REG_15_ <= n9826;
    P1_P1_REIP_REG_16_ <= n9831;
    P1_P1_REIP_REG_17_ <= n9836;
    P1_P1_REIP_REG_18_ <= n9841;
    P1_P1_REIP_REG_19_ <= n9846;
    P1_P1_REIP_REG_20_ <= n9851;
    P1_P1_REIP_REG_21_ <= n9856;
    P1_P1_REIP_REG_22_ <= n9861;
    P1_P1_REIP_REG_23_ <= n9866;
    P1_P1_REIP_REG_24_ <= n9871;
    P1_P1_REIP_REG_25_ <= n9876;
    P1_P1_REIP_REG_26_ <= n9881;
    P1_P1_REIP_REG_27_ <= n9886;
    P1_P1_REIP_REG_28_ <= n9891;
    P1_P1_REIP_REG_29_ <= n9896;
    P1_P1_REIP_REG_30_ <= n9901;
    P1_P1_REIP_REG_31_ <= n9906;
    P1_P1_BYTEENABLE_REG_3_ <= n9911;
    P1_P1_BYTEENABLE_REG_2_ <= n9916;
    P1_P1_BYTEENABLE_REG_1_ <= n9921;
    P1_P1_BYTEENABLE_REG_0_ <= n9926;
    P1_P1_W_R_N_REG <= n9931;
    P1_P1_FLUSH_REG <= n9936;
    P1_P1_MORE_REG <= n9941;
    P1_P1_STATEBS16_REG <= n9946;
    P1_P1_REQUESTPENDING_REG <= n9951;
    P1_P1_D_C_N_REG <= n9956;
    P1_P1_M_IO_N_REG <= n9961;
    P1_P1_CODEFETCH_REG <= n9966;
    P1_P1_ADS_N_REG <= n9971;
    P1_P1_READREQUEST_REG <= n9976;
    P1_P1_MEMORYFETCH_REG <= n9981;
    P2_P3_BE_N_REG_3_ <= n9986;
    P2_P3_BE_N_REG_2_ <= n9991;
    P2_P3_BE_N_REG_1_ <= n9996;
    P2_P3_BE_N_REG_0_ <= n10001;
    P2_P3_ADDRESS_REG_29_ <= n10006;
    P2_P3_ADDRESS_REG_28_ <= n10011;
    P2_P3_ADDRESS_REG_27_ <= n10016;
    P2_P3_ADDRESS_REG_26_ <= n10021;
    P2_P3_ADDRESS_REG_25_ <= n10026;
    P2_P3_ADDRESS_REG_24_ <= n10031;
    P2_P3_ADDRESS_REG_23_ <= n10036;
    P2_P3_ADDRESS_REG_22_ <= n10041;
    P2_P3_ADDRESS_REG_21_ <= n10046;
    P2_P3_ADDRESS_REG_20_ <= n10051;
    P2_P3_ADDRESS_REG_19_ <= n10056;
    P2_P3_ADDRESS_REG_18_ <= n10061;
    P2_P3_ADDRESS_REG_17_ <= n10066;
    P2_P3_ADDRESS_REG_16_ <= n10071;
    P2_P3_ADDRESS_REG_15_ <= n10076;
    P2_P3_ADDRESS_REG_14_ <= n10081;
    P2_P3_ADDRESS_REG_13_ <= n10086;
    P2_P3_ADDRESS_REG_12_ <= n10091;
    P2_P3_ADDRESS_REG_11_ <= n10096;
    P2_P3_ADDRESS_REG_10_ <= n10101;
    P2_P3_ADDRESS_REG_9_ <= n10106;
    P2_P3_ADDRESS_REG_8_ <= n10111;
    P2_P3_ADDRESS_REG_7_ <= n10116;
    P2_P3_ADDRESS_REG_6_ <= n10121;
    P2_P3_ADDRESS_REG_5_ <= n10126;
    P2_P3_ADDRESS_REG_4_ <= n10131;
    P2_P3_ADDRESS_REG_3_ <= n10136;
    P2_P3_ADDRESS_REG_2_ <= n10141;
    P2_P3_ADDRESS_REG_1_ <= n10146;
    P2_P3_ADDRESS_REG_0_ <= n10151;
    P2_P3_STATE_REG_2_ <= n10156;
    P2_P3_STATE_REG_1_ <= n10161;
    P2_P3_STATE_REG_0_ <= n10166;
    P2_P3_DATAWIDTH_REG_0_ <= n10171;
    P2_P3_DATAWIDTH_REG_1_ <= n10176;
    P2_P3_DATAWIDTH_REG_2_ <= n10181;
    P2_P3_DATAWIDTH_REG_3_ <= n10186;
    P2_P3_DATAWIDTH_REG_4_ <= n10191;
    P2_P3_DATAWIDTH_REG_5_ <= n10196;
    P2_P3_DATAWIDTH_REG_6_ <= n10201;
    P2_P3_DATAWIDTH_REG_7_ <= n10206;
    P2_P3_DATAWIDTH_REG_8_ <= n10211;
    P2_P3_DATAWIDTH_REG_9_ <= n10216;
    P2_P3_DATAWIDTH_REG_10_ <= n10221;
    P2_P3_DATAWIDTH_REG_11_ <= n10226;
    P2_P3_DATAWIDTH_REG_12_ <= n10231;
    P2_P3_DATAWIDTH_REG_13_ <= n10236;
    P2_P3_DATAWIDTH_REG_14_ <= n10241;
    P2_P3_DATAWIDTH_REG_15_ <= n10246;
    P2_P3_DATAWIDTH_REG_16_ <= n10251;
    P2_P3_DATAWIDTH_REG_17_ <= n10256;
    P2_P3_DATAWIDTH_REG_18_ <= n10261;
    P2_P3_DATAWIDTH_REG_19_ <= n10266;
    P2_P3_DATAWIDTH_REG_20_ <= n10271;
    P2_P3_DATAWIDTH_REG_21_ <= n10276;
    P2_P3_DATAWIDTH_REG_22_ <= n10281;
    P2_P3_DATAWIDTH_REG_23_ <= n10286;
    P2_P3_DATAWIDTH_REG_24_ <= n10291;
    P2_P3_DATAWIDTH_REG_25_ <= n10296;
    P2_P3_DATAWIDTH_REG_26_ <= n10301;
    P2_P3_DATAWIDTH_REG_27_ <= n10306;
    P2_P3_DATAWIDTH_REG_28_ <= n10311;
    P2_P3_DATAWIDTH_REG_29_ <= n10316;
    P2_P3_DATAWIDTH_REG_30_ <= n10321;
    P2_P3_DATAWIDTH_REG_31_ <= n10326;
    P2_P3_STATE2_REG_3_ <= n10331;
    P2_P3_STATE2_REG_2_ <= n10336;
    P2_P3_STATE2_REG_1_ <= n10341;
    P2_P3_STATE2_REG_0_ <= n10346;
    P2_P3_INSTQUEUE_REG_15__7_ <= n10351;
    P2_P3_INSTQUEUE_REG_15__6_ <= n10356;
    P2_P3_INSTQUEUE_REG_15__5_ <= n10361;
    P2_P3_INSTQUEUE_REG_15__4_ <= n10366;
    P2_P3_INSTQUEUE_REG_15__3_ <= n10371;
    P2_P3_INSTQUEUE_REG_15__2_ <= n10376;
    P2_P3_INSTQUEUE_REG_15__1_ <= n10381;
    P2_P3_INSTQUEUE_REG_15__0_ <= n10386;
    P2_P3_INSTQUEUE_REG_14__7_ <= n10391;
    P2_P3_INSTQUEUE_REG_14__6_ <= n10396;
    P2_P3_INSTQUEUE_REG_14__5_ <= n10401;
    P2_P3_INSTQUEUE_REG_14__4_ <= n10406;
    P2_P3_INSTQUEUE_REG_14__3_ <= n10411;
    P2_P3_INSTQUEUE_REG_14__2_ <= n10416;
    P2_P3_INSTQUEUE_REG_14__1_ <= n10421;
    P2_P3_INSTQUEUE_REG_14__0_ <= n10426;
    P2_P3_INSTQUEUE_REG_13__7_ <= n10431;
    P2_P3_INSTQUEUE_REG_13__6_ <= n10436;
    P2_P3_INSTQUEUE_REG_13__5_ <= n10441;
    P2_P3_INSTQUEUE_REG_13__4_ <= n10446;
    P2_P3_INSTQUEUE_REG_13__3_ <= n10451;
    P2_P3_INSTQUEUE_REG_13__2_ <= n10456;
    P2_P3_INSTQUEUE_REG_13__1_ <= n10461;
    P2_P3_INSTQUEUE_REG_13__0_ <= n10466;
    P2_P3_INSTQUEUE_REG_12__7_ <= n10471;
    P2_P3_INSTQUEUE_REG_12__6_ <= n10476;
    P2_P3_INSTQUEUE_REG_12__5_ <= n10481;
    P2_P3_INSTQUEUE_REG_12__4_ <= n10486;
    P2_P3_INSTQUEUE_REG_12__3_ <= n10491;
    P2_P3_INSTQUEUE_REG_12__2_ <= n10496;
    P2_P3_INSTQUEUE_REG_12__1_ <= n10501;
    P2_P3_INSTQUEUE_REG_12__0_ <= n10506;
    P2_P3_INSTQUEUE_REG_11__7_ <= n10511;
    P2_P3_INSTQUEUE_REG_11__6_ <= n10516;
    P2_P3_INSTQUEUE_REG_11__5_ <= n10521;
    P2_P3_INSTQUEUE_REG_11__4_ <= n10526;
    P2_P3_INSTQUEUE_REG_11__3_ <= n10531;
    P2_P3_INSTQUEUE_REG_11__2_ <= n10536;
    P2_P3_INSTQUEUE_REG_11__1_ <= n10541;
    P2_P3_INSTQUEUE_REG_11__0_ <= n10546;
    P2_P3_INSTQUEUE_REG_10__7_ <= n10551;
    P2_P3_INSTQUEUE_REG_10__6_ <= n10556;
    P2_P3_INSTQUEUE_REG_10__5_ <= n10561;
    P2_P3_INSTQUEUE_REG_10__4_ <= n10566;
    P2_P3_INSTQUEUE_REG_10__3_ <= n10571;
    P2_P3_INSTQUEUE_REG_10__2_ <= n10576;
    P2_P3_INSTQUEUE_REG_10__1_ <= n10581;
    P2_P3_INSTQUEUE_REG_10__0_ <= n10586;
    P2_P3_INSTQUEUE_REG_9__7_ <= n10591;
    P2_P3_INSTQUEUE_REG_9__6_ <= n10596;
    P2_P3_INSTQUEUE_REG_9__5_ <= n10601;
    P2_P3_INSTQUEUE_REG_9__4_ <= n10606;
    P2_P3_INSTQUEUE_REG_9__3_ <= n10611;
    P2_P3_INSTQUEUE_REG_9__2_ <= n10616;
    P2_P3_INSTQUEUE_REG_9__1_ <= n10621;
    P2_P3_INSTQUEUE_REG_9__0_ <= n10626;
    P2_P3_INSTQUEUE_REG_8__7_ <= n10631;
    P2_P3_INSTQUEUE_REG_8__6_ <= n10636;
    P2_P3_INSTQUEUE_REG_8__5_ <= n10641;
    P2_P3_INSTQUEUE_REG_8__4_ <= n10646;
    P2_P3_INSTQUEUE_REG_8__3_ <= n10651;
    P2_P3_INSTQUEUE_REG_8__2_ <= n10656;
    P2_P3_INSTQUEUE_REG_8__1_ <= n10661;
    P2_P3_INSTQUEUE_REG_8__0_ <= n10666;
    P2_P3_INSTQUEUE_REG_7__7_ <= n10671;
    P2_P3_INSTQUEUE_REG_7__6_ <= n10676;
    P2_P3_INSTQUEUE_REG_7__5_ <= n10681;
    P2_P3_INSTQUEUE_REG_7__4_ <= n10686;
    P2_P3_INSTQUEUE_REG_7__3_ <= n10691;
    P2_P3_INSTQUEUE_REG_7__2_ <= n10696;
    P2_P3_INSTQUEUE_REG_7__1_ <= n10701;
    P2_P3_INSTQUEUE_REG_7__0_ <= n10706;
    P2_P3_INSTQUEUE_REG_6__7_ <= n10711;
    P2_P3_INSTQUEUE_REG_6__6_ <= n10716;
    P2_P3_INSTQUEUE_REG_6__5_ <= n10721;
    P2_P3_INSTQUEUE_REG_6__4_ <= n10726;
    P2_P3_INSTQUEUE_REG_6__3_ <= n10731;
    P2_P3_INSTQUEUE_REG_6__2_ <= n10736;
    P2_P3_INSTQUEUE_REG_6__1_ <= n10741;
    P2_P3_INSTQUEUE_REG_6__0_ <= n10746;
    P2_P3_INSTQUEUE_REG_5__7_ <= n10751;
    P2_P3_INSTQUEUE_REG_5__6_ <= n10756;
    P2_P3_INSTQUEUE_REG_5__5_ <= n10761;
    P2_P3_INSTQUEUE_REG_5__4_ <= n10766;
    P2_P3_INSTQUEUE_REG_5__3_ <= n10771;
    P2_P3_INSTQUEUE_REG_5__2_ <= n10776;
    P2_P3_INSTQUEUE_REG_5__1_ <= n10781;
    P2_P3_INSTQUEUE_REG_5__0_ <= n10786;
    P2_P3_INSTQUEUE_REG_4__7_ <= n10791;
    P2_P3_INSTQUEUE_REG_4__6_ <= n10796;
    P2_P3_INSTQUEUE_REG_4__5_ <= n10801;
    P2_P3_INSTQUEUE_REG_4__4_ <= n10806;
    P2_P3_INSTQUEUE_REG_4__3_ <= n10811;
    P2_P3_INSTQUEUE_REG_4__2_ <= n10816;
    P2_P3_INSTQUEUE_REG_4__1_ <= n10821;
    P2_P3_INSTQUEUE_REG_4__0_ <= n10826;
    P2_P3_INSTQUEUE_REG_3__7_ <= n10831;
    P2_P3_INSTQUEUE_REG_3__6_ <= n10836;
    P2_P3_INSTQUEUE_REG_3__5_ <= n10841;
    P2_P3_INSTQUEUE_REG_3__4_ <= n10846;
    P2_P3_INSTQUEUE_REG_3__3_ <= n10851;
    P2_P3_INSTQUEUE_REG_3__2_ <= n10856;
    P2_P3_INSTQUEUE_REG_3__1_ <= n10861;
    P2_P3_INSTQUEUE_REG_3__0_ <= n10866;
    P2_P3_INSTQUEUE_REG_2__7_ <= n10871;
    P2_P3_INSTQUEUE_REG_2__6_ <= n10876;
    P2_P3_INSTQUEUE_REG_2__5_ <= n10881;
    P2_P3_INSTQUEUE_REG_2__4_ <= n10886;
    P2_P3_INSTQUEUE_REG_2__3_ <= n10891;
    P2_P3_INSTQUEUE_REG_2__2_ <= n10896;
    P2_P3_INSTQUEUE_REG_2__1_ <= n10901;
    P2_P3_INSTQUEUE_REG_2__0_ <= n10906;
    P2_P3_INSTQUEUE_REG_1__7_ <= n10911;
    P2_P3_INSTQUEUE_REG_1__6_ <= n10916;
    P2_P3_INSTQUEUE_REG_1__5_ <= n10921;
    P2_P3_INSTQUEUE_REG_1__4_ <= n10926;
    P2_P3_INSTQUEUE_REG_1__3_ <= n10931;
    P2_P3_INSTQUEUE_REG_1__2_ <= n10936;
    P2_P3_INSTQUEUE_REG_1__1_ <= n10941;
    P2_P3_INSTQUEUE_REG_1__0_ <= n10946;
    P2_P3_INSTQUEUE_REG_0__7_ <= n10951;
    P2_P3_INSTQUEUE_REG_0__6_ <= n10956;
    P2_P3_INSTQUEUE_REG_0__5_ <= n10961;
    P2_P3_INSTQUEUE_REG_0__4_ <= n10966;
    P2_P3_INSTQUEUE_REG_0__3_ <= n10971;
    P2_P3_INSTQUEUE_REG_0__2_ <= n10976;
    P2_P3_INSTQUEUE_REG_0__1_ <= n10981;
    P2_P3_INSTQUEUE_REG_0__0_ <= n10986;
    P2_P3_INSTQUEUERD_ADDR_REG_4_ <= n10991;
    P2_P3_INSTQUEUERD_ADDR_REG_3_ <= n10996;
    P2_P3_INSTQUEUERD_ADDR_REG_2_ <= n11001;
    P2_P3_INSTQUEUERD_ADDR_REG_1_ <= n11006;
    P2_P3_INSTQUEUERD_ADDR_REG_0_ <= n11011;
    P2_P3_INSTQUEUEWR_ADDR_REG_4_ <= n11016;
    P2_P3_INSTQUEUEWR_ADDR_REG_3_ <= n11021;
    P2_P3_INSTQUEUEWR_ADDR_REG_2_ <= n11026;
    P2_P3_INSTQUEUEWR_ADDR_REG_1_ <= n11031;
    P2_P3_INSTQUEUEWR_ADDR_REG_0_ <= n11036;
    P2_P3_INSTADDRPOINTER_REG_0_ <= n11041;
    P2_P3_INSTADDRPOINTER_REG_1_ <= n11046;
    P2_P3_INSTADDRPOINTER_REG_2_ <= n11051;
    P2_P3_INSTADDRPOINTER_REG_3_ <= n11056;
    P2_P3_INSTADDRPOINTER_REG_4_ <= n11061;
    P2_P3_INSTADDRPOINTER_REG_5_ <= n11066;
    P2_P3_INSTADDRPOINTER_REG_6_ <= n11071;
    P2_P3_INSTADDRPOINTER_REG_7_ <= n11076;
    P2_P3_INSTADDRPOINTER_REG_8_ <= n11081;
    P2_P3_INSTADDRPOINTER_REG_9_ <= n11086;
    P2_P3_INSTADDRPOINTER_REG_10_ <= n11091;
    P2_P3_INSTADDRPOINTER_REG_11_ <= n11096;
    P2_P3_INSTADDRPOINTER_REG_12_ <= n11101;
    P2_P3_INSTADDRPOINTER_REG_13_ <= n11106;
    P2_P3_INSTADDRPOINTER_REG_14_ <= n11111;
    P2_P3_INSTADDRPOINTER_REG_15_ <= n11116;
    P2_P3_INSTADDRPOINTER_REG_16_ <= n11121;
    P2_P3_INSTADDRPOINTER_REG_17_ <= n11126;
    P2_P3_INSTADDRPOINTER_REG_18_ <= n11131;
    P2_P3_INSTADDRPOINTER_REG_19_ <= n11136;
    P2_P3_INSTADDRPOINTER_REG_20_ <= n11141;
    P2_P3_INSTADDRPOINTER_REG_21_ <= n11146;
    P2_P3_INSTADDRPOINTER_REG_22_ <= n11151;
    P2_P3_INSTADDRPOINTER_REG_23_ <= n11156;
    P2_P3_INSTADDRPOINTER_REG_24_ <= n11161;
    P2_P3_INSTADDRPOINTER_REG_25_ <= n11166;
    P2_P3_INSTADDRPOINTER_REG_26_ <= n11171;
    P2_P3_INSTADDRPOINTER_REG_27_ <= n11176;
    P2_P3_INSTADDRPOINTER_REG_28_ <= n11181;
    P2_P3_INSTADDRPOINTER_REG_29_ <= n11186;
    P2_P3_INSTADDRPOINTER_REG_30_ <= n11191;
    P2_P3_INSTADDRPOINTER_REG_31_ <= n11196;
    P2_P3_PHYADDRPOINTER_REG_0_ <= n11201;
    P2_P3_PHYADDRPOINTER_REG_1_ <= n11206;
    P2_P3_PHYADDRPOINTER_REG_2_ <= n11211;
    P2_P3_PHYADDRPOINTER_REG_3_ <= n11216;
    P2_P3_PHYADDRPOINTER_REG_4_ <= n11221;
    P2_P3_PHYADDRPOINTER_REG_5_ <= n11226;
    P2_P3_PHYADDRPOINTER_REG_6_ <= n11231;
    P2_P3_PHYADDRPOINTER_REG_7_ <= n11236;
    P2_P3_PHYADDRPOINTER_REG_8_ <= n11241;
    P2_P3_PHYADDRPOINTER_REG_9_ <= n11246;
    P2_P3_PHYADDRPOINTER_REG_10_ <= n11251;
    P2_P3_PHYADDRPOINTER_REG_11_ <= n11256;
    P2_P3_PHYADDRPOINTER_REG_12_ <= n11261;
    P2_P3_PHYADDRPOINTER_REG_13_ <= n11266;
    P2_P3_PHYADDRPOINTER_REG_14_ <= n11271;
    P2_P3_PHYADDRPOINTER_REG_15_ <= n11276;
    P2_P3_PHYADDRPOINTER_REG_16_ <= n11281;
    P2_P3_PHYADDRPOINTER_REG_17_ <= n11286;
    P2_P3_PHYADDRPOINTER_REG_18_ <= n11291;
    P2_P3_PHYADDRPOINTER_REG_19_ <= n11296;
    P2_P3_PHYADDRPOINTER_REG_20_ <= n11301;
    P2_P3_PHYADDRPOINTER_REG_21_ <= n11306;
    P2_P3_PHYADDRPOINTER_REG_22_ <= n11311;
    P2_P3_PHYADDRPOINTER_REG_23_ <= n11316;
    P2_P3_PHYADDRPOINTER_REG_24_ <= n11321;
    P2_P3_PHYADDRPOINTER_REG_25_ <= n11326;
    P2_P3_PHYADDRPOINTER_REG_26_ <= n11331;
    P2_P3_PHYADDRPOINTER_REG_27_ <= n11336;
    P2_P3_PHYADDRPOINTER_REG_28_ <= n11341;
    P2_P3_PHYADDRPOINTER_REG_29_ <= n11346;
    P2_P3_PHYADDRPOINTER_REG_30_ <= n11351;
    P2_P3_PHYADDRPOINTER_REG_31_ <= n11356;
    P2_P3_LWORD_REG_15_ <= n11361;
    P2_P3_LWORD_REG_14_ <= n11366;
    P2_P3_LWORD_REG_13_ <= n11371;
    P2_P3_LWORD_REG_12_ <= n11376;
    P2_P3_LWORD_REG_11_ <= n11381;
    P2_P3_LWORD_REG_10_ <= n11386;
    P2_P3_LWORD_REG_9_ <= n11391;
    P2_P3_LWORD_REG_8_ <= n11396;
    P2_P3_LWORD_REG_7_ <= n11401;
    P2_P3_LWORD_REG_6_ <= n11406;
    P2_P3_LWORD_REG_5_ <= n11411;
    P2_P3_LWORD_REG_4_ <= n11416;
    P2_P3_LWORD_REG_3_ <= n11421;
    P2_P3_LWORD_REG_2_ <= n11426;
    P2_P3_LWORD_REG_1_ <= n11431;
    P2_P3_LWORD_REG_0_ <= n11436;
    P2_P3_UWORD_REG_14_ <= n11441;
    P2_P3_UWORD_REG_13_ <= n11446;
    P2_P3_UWORD_REG_12_ <= n11451;
    P2_P3_UWORD_REG_11_ <= n11456;
    P2_P3_UWORD_REG_10_ <= n11461;
    P2_P3_UWORD_REG_9_ <= n11466;
    P2_P3_UWORD_REG_8_ <= n11471;
    P2_P3_UWORD_REG_7_ <= n11476;
    P2_P3_UWORD_REG_6_ <= n11481;
    P2_P3_UWORD_REG_5_ <= n11486;
    P2_P3_UWORD_REG_4_ <= n11491;
    P2_P3_UWORD_REG_3_ <= n11496;
    P2_P3_UWORD_REG_2_ <= n11501;
    P2_P3_UWORD_REG_1_ <= n11506;
    P2_P3_UWORD_REG_0_ <= n11511;
    P2_P3_DATAO_REG_0_ <= n11516;
    P2_P3_DATAO_REG_1_ <= n11521;
    P2_P3_DATAO_REG_2_ <= n11526;
    P2_P3_DATAO_REG_3_ <= n11531;
    P2_P3_DATAO_REG_4_ <= n11536;
    P2_P3_DATAO_REG_5_ <= n11541;
    P2_P3_DATAO_REG_6_ <= n11546;
    P2_P3_DATAO_REG_7_ <= n11551;
    P2_P3_DATAO_REG_8_ <= n11556;
    P2_P3_DATAO_REG_9_ <= n11561;
    P2_P3_DATAO_REG_10_ <= n11566;
    P2_P3_DATAO_REG_11_ <= n11571;
    P2_P3_DATAO_REG_12_ <= n11576;
    P2_P3_DATAO_REG_13_ <= n11581;
    P2_P3_DATAO_REG_14_ <= n11586;
    P2_P3_DATAO_REG_15_ <= n11591;
    P2_P3_DATAO_REG_16_ <= n11596;
    P2_P3_DATAO_REG_17_ <= n11601;
    P2_P3_DATAO_REG_18_ <= n11606;
    P2_P3_DATAO_REG_19_ <= n11611;
    P2_P3_DATAO_REG_20_ <= n11616;
    P2_P3_DATAO_REG_21_ <= n11621;
    P2_P3_DATAO_REG_22_ <= n11626;
    P2_P3_DATAO_REG_23_ <= n11631;
    P2_P3_DATAO_REG_24_ <= n11636;
    P2_P3_DATAO_REG_25_ <= n11641;
    P2_P3_DATAO_REG_26_ <= n11646;
    P2_P3_DATAO_REG_27_ <= n11651;
    P2_P3_DATAO_REG_28_ <= n11656;
    P2_P3_DATAO_REG_29_ <= n11661;
    P2_P3_DATAO_REG_30_ <= n11666;
    P2_P3_DATAO_REG_31_ <= n11671;
    P2_P3_EAX_REG_0_ <= n11676;
    P2_P3_EAX_REG_1_ <= n11681;
    P2_P3_EAX_REG_2_ <= n11686;
    P2_P3_EAX_REG_3_ <= n11691;
    P2_P3_EAX_REG_4_ <= n11696;
    P2_P3_EAX_REG_5_ <= n11701;
    P2_P3_EAX_REG_6_ <= n11706;
    P2_P3_EAX_REG_7_ <= n11711;
    P2_P3_EAX_REG_8_ <= n11716;
    P2_P3_EAX_REG_9_ <= n11721;
    P2_P3_EAX_REG_10_ <= n11726;
    P2_P3_EAX_REG_11_ <= n11731;
    P2_P3_EAX_REG_12_ <= n11736;
    P2_P3_EAX_REG_13_ <= n11741;
    P2_P3_EAX_REG_14_ <= n11746;
    P2_P3_EAX_REG_15_ <= n11751;
    P2_P3_EAX_REG_16_ <= n11756;
    P2_P3_EAX_REG_17_ <= n11761;
    P2_P3_EAX_REG_18_ <= n11766;
    P2_P3_EAX_REG_19_ <= n11771;
    P2_P3_EAX_REG_20_ <= n11776;
    P2_P3_EAX_REG_21_ <= n11781;
    P2_P3_EAX_REG_22_ <= n11786;
    P2_P3_EAX_REG_23_ <= n11791;
    P2_P3_EAX_REG_24_ <= n11796;
    P2_P3_EAX_REG_25_ <= n11801;
    P2_P3_EAX_REG_26_ <= n11806;
    P2_P3_EAX_REG_27_ <= n11811;
    P2_P3_EAX_REG_28_ <= n11816;
    P2_P3_EAX_REG_29_ <= n11821;
    P2_P3_EAX_REG_30_ <= n11826;
    P2_P3_EAX_REG_31_ <= n11831;
    P2_P3_EBX_REG_0_ <= n11836;
    P2_P3_EBX_REG_1_ <= n11841;
    P2_P3_EBX_REG_2_ <= n11846;
    P2_P3_EBX_REG_3_ <= n11851;
    P2_P3_EBX_REG_4_ <= n11856;
    P2_P3_EBX_REG_5_ <= n11861;
    P2_P3_EBX_REG_6_ <= n11866;
    P2_P3_EBX_REG_7_ <= n11871;
    P2_P3_EBX_REG_8_ <= n11876;
    P2_P3_EBX_REG_9_ <= n11881;
    P2_P3_EBX_REG_10_ <= n11886;
    P2_P3_EBX_REG_11_ <= n11891;
    P2_P3_EBX_REG_12_ <= n11896;
    P2_P3_EBX_REG_13_ <= n11901;
    P2_P3_EBX_REG_14_ <= n11906;
    P2_P3_EBX_REG_15_ <= n11911;
    P2_P3_EBX_REG_16_ <= n11916;
    P2_P3_EBX_REG_17_ <= n11921;
    P2_P3_EBX_REG_18_ <= n11926;
    P2_P3_EBX_REG_19_ <= n11931;
    P2_P3_EBX_REG_20_ <= n11936;
    P2_P3_EBX_REG_21_ <= n11941;
    P2_P3_EBX_REG_22_ <= n11946;
    P2_P3_EBX_REG_23_ <= n11951;
    P2_P3_EBX_REG_24_ <= n11956;
    P2_P3_EBX_REG_25_ <= n11961;
    P2_P3_EBX_REG_26_ <= n11966;
    P2_P3_EBX_REG_27_ <= n11971;
    P2_P3_EBX_REG_28_ <= n11976;
    P2_P3_EBX_REG_29_ <= n11981;
    P2_P3_EBX_REG_30_ <= n11986;
    P2_P3_EBX_REG_31_ <= n11991;
    P2_P3_REIP_REG_0_ <= n11996;
    P2_P3_REIP_REG_1_ <= n12001;
    P2_P3_REIP_REG_2_ <= n12006;
    P2_P3_REIP_REG_3_ <= n12011;
    P2_P3_REIP_REG_4_ <= n12016;
    P2_P3_REIP_REG_5_ <= n12021;
    P2_P3_REIP_REG_6_ <= n12026;
    P2_P3_REIP_REG_7_ <= n12031;
    P2_P3_REIP_REG_8_ <= n12036;
    P2_P3_REIP_REG_9_ <= n12041;
    P2_P3_REIP_REG_10_ <= n12046;
    P2_P3_REIP_REG_11_ <= n12051;
    P2_P3_REIP_REG_12_ <= n12056;
    P2_P3_REIP_REG_13_ <= n12061;
    P2_P3_REIP_REG_14_ <= n12066;
    P2_P3_REIP_REG_15_ <= n12071;
    P2_P3_REIP_REG_16_ <= n12076;
    P2_P3_REIP_REG_17_ <= n12081;
    P2_P3_REIP_REG_18_ <= n12086;
    P2_P3_REIP_REG_19_ <= n12091;
    P2_P3_REIP_REG_20_ <= n12096;
    P2_P3_REIP_REG_21_ <= n12101;
    P2_P3_REIP_REG_22_ <= n12106;
    P2_P3_REIP_REG_23_ <= n12111;
    P2_P3_REIP_REG_24_ <= n12116;
    P2_P3_REIP_REG_25_ <= n12121;
    P2_P3_REIP_REG_26_ <= n12126;
    P2_P3_REIP_REG_27_ <= n12131;
    P2_P3_REIP_REG_28_ <= n12136;
    P2_P3_REIP_REG_29_ <= n12141;
    P2_P3_REIP_REG_30_ <= n12146;
    P2_P3_REIP_REG_31_ <= n12151;
    P2_P3_BYTEENABLE_REG_3_ <= n12156;
    P2_P3_BYTEENABLE_REG_2_ <= n12161;
    P2_P3_BYTEENABLE_REG_1_ <= n12166;
    P2_P3_BYTEENABLE_REG_0_ <= n12171;
    P2_P3_W_R_N_REG <= n12176;
    P2_P3_FLUSH_REG <= n12181;
    P2_P3_MORE_REG <= n12186;
    P2_P3_STATEBS16_REG <= n12191;
    P2_P3_REQUESTPENDING_REG <= n12196;
    P2_P3_D_C_N_REG <= n12201;
    P2_P3_M_IO_N_REG <= n12206;
    P2_P3_CODEFETCH_REG <= n12211;
    P2_P3_ADS_N_REG <= n12216;
    P2_P3_READREQUEST_REG <= n12221;
    P2_P3_MEMORYFETCH_REG <= n12226;
    P2_P2_BE_N_REG_3_ <= n12231;
    P2_P2_BE_N_REG_2_ <= n12236;
    P2_P2_BE_N_REG_1_ <= n12241;
    P2_P2_BE_N_REG_0_ <= n12246;
    P2_P2_ADDRESS_REG_29_ <= n12251;
    P2_P2_ADDRESS_REG_28_ <= n12256;
    P2_P2_ADDRESS_REG_27_ <= n12261;
    P2_P2_ADDRESS_REG_26_ <= n12266;
    P2_P2_ADDRESS_REG_25_ <= n12271;
    P2_P2_ADDRESS_REG_24_ <= n12276;
    P2_P2_ADDRESS_REG_23_ <= n12281;
    P2_P2_ADDRESS_REG_22_ <= n12286;
    P2_P2_ADDRESS_REG_21_ <= n12291;
    P2_P2_ADDRESS_REG_20_ <= n12296;
    P2_P2_ADDRESS_REG_19_ <= n12301;
    P2_P2_ADDRESS_REG_18_ <= n12306;
    P2_P2_ADDRESS_REG_17_ <= n12311;
    P2_P2_ADDRESS_REG_16_ <= n12316;
    P2_P2_ADDRESS_REG_15_ <= n12321;
    P2_P2_ADDRESS_REG_14_ <= n12326;
    P2_P2_ADDRESS_REG_13_ <= n12331;
    P2_P2_ADDRESS_REG_12_ <= n12336;
    P2_P2_ADDRESS_REG_11_ <= n12341;
    P2_P2_ADDRESS_REG_10_ <= n12346;
    P2_P2_ADDRESS_REG_9_ <= n12351;
    P2_P2_ADDRESS_REG_8_ <= n12356;
    P2_P2_ADDRESS_REG_7_ <= n12361;
    P2_P2_ADDRESS_REG_6_ <= n12366;
    P2_P2_ADDRESS_REG_5_ <= n12371;
    P2_P2_ADDRESS_REG_4_ <= n12376;
    P2_P2_ADDRESS_REG_3_ <= n12381;
    P2_P2_ADDRESS_REG_2_ <= n12386;
    P2_P2_ADDRESS_REG_1_ <= n12391;
    P2_P2_ADDRESS_REG_0_ <= n12396;
    P2_P2_STATE_REG_2_ <= n12401;
    P2_P2_STATE_REG_1_ <= n12406;
    P2_P2_STATE_REG_0_ <= n12411;
    P2_P2_DATAWIDTH_REG_0_ <= n12416;
    P2_P2_DATAWIDTH_REG_1_ <= n12421;
    P2_P2_DATAWIDTH_REG_2_ <= n12426;
    P2_P2_DATAWIDTH_REG_3_ <= n12431;
    P2_P2_DATAWIDTH_REG_4_ <= n12436;
    P2_P2_DATAWIDTH_REG_5_ <= n12441;
    P2_P2_DATAWIDTH_REG_6_ <= n12446;
    P2_P2_DATAWIDTH_REG_7_ <= n12451;
    P2_P2_DATAWIDTH_REG_8_ <= n12456;
    P2_P2_DATAWIDTH_REG_9_ <= n12461;
    P2_P2_DATAWIDTH_REG_10_ <= n12466;
    P2_P2_DATAWIDTH_REG_11_ <= n12471;
    P2_P2_DATAWIDTH_REG_12_ <= n12476;
    P2_P2_DATAWIDTH_REG_13_ <= n12481;
    P2_P2_DATAWIDTH_REG_14_ <= n12486;
    P2_P2_DATAWIDTH_REG_15_ <= n12491;
    P2_P2_DATAWIDTH_REG_16_ <= n12496;
    P2_P2_DATAWIDTH_REG_17_ <= n12501;
    P2_P2_DATAWIDTH_REG_18_ <= n12506;
    P2_P2_DATAWIDTH_REG_19_ <= n12511;
    P2_P2_DATAWIDTH_REG_20_ <= n12516;
    P2_P2_DATAWIDTH_REG_21_ <= n12521;
    P2_P2_DATAWIDTH_REG_22_ <= n12526;
    P2_P2_DATAWIDTH_REG_23_ <= n12531;
    P2_P2_DATAWIDTH_REG_24_ <= n12536;
    P2_P2_DATAWIDTH_REG_25_ <= n12541;
    P2_P2_DATAWIDTH_REG_26_ <= n12546;
    P2_P2_DATAWIDTH_REG_27_ <= n12551;
    P2_P2_DATAWIDTH_REG_28_ <= n12556;
    P2_P2_DATAWIDTH_REG_29_ <= n12561;
    P2_P2_DATAWIDTH_REG_30_ <= n12566;
    P2_P2_DATAWIDTH_REG_31_ <= n12571;
    P2_P2_STATE2_REG_3_ <= n12576;
    P2_P2_STATE2_REG_2_ <= n12581;
    P2_P2_STATE2_REG_1_ <= n12586;
    P2_P2_STATE2_REG_0_ <= n12591;
    P2_P2_INSTQUEUE_REG_15__7_ <= n12596;
    P2_P2_INSTQUEUE_REG_15__6_ <= n12601;
    P2_P2_INSTQUEUE_REG_15__5_ <= n12606;
    P2_P2_INSTQUEUE_REG_15__4_ <= n12611;
    P2_P2_INSTQUEUE_REG_15__3_ <= n12616;
    P2_P2_INSTQUEUE_REG_15__2_ <= n12621;
    P2_P2_INSTQUEUE_REG_15__1_ <= n12626;
    P2_P2_INSTQUEUE_REG_15__0_ <= n12631;
    P2_P2_INSTQUEUE_REG_14__7_ <= n12636;
    P2_P2_INSTQUEUE_REG_14__6_ <= n12641;
    P2_P2_INSTQUEUE_REG_14__5_ <= n12646;
    P2_P2_INSTQUEUE_REG_14__4_ <= n12651;
    P2_P2_INSTQUEUE_REG_14__3_ <= n12656;
    P2_P2_INSTQUEUE_REG_14__2_ <= n12661;
    P2_P2_INSTQUEUE_REG_14__1_ <= n12666;
    P2_P2_INSTQUEUE_REG_14__0_ <= n12671;
    P2_P2_INSTQUEUE_REG_13__7_ <= n12676;
    P2_P2_INSTQUEUE_REG_13__6_ <= n12681;
    P2_P2_INSTQUEUE_REG_13__5_ <= n12686;
    P2_P2_INSTQUEUE_REG_13__4_ <= n12691;
    P2_P2_INSTQUEUE_REG_13__3_ <= n12696;
    P2_P2_INSTQUEUE_REG_13__2_ <= n12701;
    P2_P2_INSTQUEUE_REG_13__1_ <= n12706;
    P2_P2_INSTQUEUE_REG_13__0_ <= n12711;
    P2_P2_INSTQUEUE_REG_12__7_ <= n12716;
    P2_P2_INSTQUEUE_REG_12__6_ <= n12721;
    P2_P2_INSTQUEUE_REG_12__5_ <= n12726;
    P2_P2_INSTQUEUE_REG_12__4_ <= n12731;
    P2_P2_INSTQUEUE_REG_12__3_ <= n12736;
    P2_P2_INSTQUEUE_REG_12__2_ <= n12741;
    P2_P2_INSTQUEUE_REG_12__1_ <= n12746;
    P2_P2_INSTQUEUE_REG_12__0_ <= n12751;
    P2_P2_INSTQUEUE_REG_11__7_ <= n12756;
    P2_P2_INSTQUEUE_REG_11__6_ <= n12761;
    P2_P2_INSTQUEUE_REG_11__5_ <= n12766;
    P2_P2_INSTQUEUE_REG_11__4_ <= n12771;
    P2_P2_INSTQUEUE_REG_11__3_ <= n12776;
    P2_P2_INSTQUEUE_REG_11__2_ <= n12781;
    P2_P2_INSTQUEUE_REG_11__1_ <= n12786;
    P2_P2_INSTQUEUE_REG_11__0_ <= n12791;
    P2_P2_INSTQUEUE_REG_10__7_ <= n12796;
    P2_P2_INSTQUEUE_REG_10__6_ <= n12801;
    P2_P2_INSTQUEUE_REG_10__5_ <= n12806;
    P2_P2_INSTQUEUE_REG_10__4_ <= n12811;
    P2_P2_INSTQUEUE_REG_10__3_ <= n12816;
    P2_P2_INSTQUEUE_REG_10__2_ <= n12821;
    P2_P2_INSTQUEUE_REG_10__1_ <= n12826;
    P2_P2_INSTQUEUE_REG_10__0_ <= n12831;
    P2_P2_INSTQUEUE_REG_9__7_ <= n12836;
    P2_P2_INSTQUEUE_REG_9__6_ <= n12841;
    P2_P2_INSTQUEUE_REG_9__5_ <= n12846;
    P2_P2_INSTQUEUE_REG_9__4_ <= n12851;
    P2_P2_INSTQUEUE_REG_9__3_ <= n12856;
    P2_P2_INSTQUEUE_REG_9__2_ <= n12861;
    P2_P2_INSTQUEUE_REG_9__1_ <= n12866;
    P2_P2_INSTQUEUE_REG_9__0_ <= n12871;
    P2_P2_INSTQUEUE_REG_8__7_ <= n12876;
    P2_P2_INSTQUEUE_REG_8__6_ <= n12881;
    P2_P2_INSTQUEUE_REG_8__5_ <= n12886;
    P2_P2_INSTQUEUE_REG_8__4_ <= n12891;
    P2_P2_INSTQUEUE_REG_8__3_ <= n12896;
    P2_P2_INSTQUEUE_REG_8__2_ <= n12901;
    P2_P2_INSTQUEUE_REG_8__1_ <= n12906;
    P2_P2_INSTQUEUE_REG_8__0_ <= n12911;
    P2_P2_INSTQUEUE_REG_7__7_ <= n12916;
    P2_P2_INSTQUEUE_REG_7__6_ <= n12921;
    P2_P2_INSTQUEUE_REG_7__5_ <= n12926;
    P2_P2_INSTQUEUE_REG_7__4_ <= n12931;
    P2_P2_INSTQUEUE_REG_7__3_ <= n12936;
    P2_P2_INSTQUEUE_REG_7__2_ <= n12941;
    P2_P2_INSTQUEUE_REG_7__1_ <= n12946;
    P2_P2_INSTQUEUE_REG_7__0_ <= n12951;
    P2_P2_INSTQUEUE_REG_6__7_ <= n12956;
    P2_P2_INSTQUEUE_REG_6__6_ <= n12961;
    P2_P2_INSTQUEUE_REG_6__5_ <= n12966;
    P2_P2_INSTQUEUE_REG_6__4_ <= n12971;
    P2_P2_INSTQUEUE_REG_6__3_ <= n12976;
    P2_P2_INSTQUEUE_REG_6__2_ <= n12981;
    P2_P2_INSTQUEUE_REG_6__1_ <= n12986;
    P2_P2_INSTQUEUE_REG_6__0_ <= n12991;
    P2_P2_INSTQUEUE_REG_5__7_ <= n12996;
    P2_P2_INSTQUEUE_REG_5__6_ <= n13001;
    P2_P2_INSTQUEUE_REG_5__5_ <= n13006;
    P2_P2_INSTQUEUE_REG_5__4_ <= n13011;
    P2_P2_INSTQUEUE_REG_5__3_ <= n13016;
    P2_P2_INSTQUEUE_REG_5__2_ <= n13021;
    P2_P2_INSTQUEUE_REG_5__1_ <= n13026;
    P2_P2_INSTQUEUE_REG_5__0_ <= n13031;
    P2_P2_INSTQUEUE_REG_4__7_ <= n13036;
    P2_P2_INSTQUEUE_REG_4__6_ <= n13041;
    P2_P2_INSTQUEUE_REG_4__5_ <= n13046;
    P2_P2_INSTQUEUE_REG_4__4_ <= n13051;
    P2_P2_INSTQUEUE_REG_4__3_ <= n13056;
    P2_P2_INSTQUEUE_REG_4__2_ <= n13061;
    P2_P2_INSTQUEUE_REG_4__1_ <= n13066;
    P2_P2_INSTQUEUE_REG_4__0_ <= n13071;
    P2_P2_INSTQUEUE_REG_3__7_ <= n13076;
    P2_P2_INSTQUEUE_REG_3__6_ <= n13081;
    P2_P2_INSTQUEUE_REG_3__5_ <= n13086;
    P2_P2_INSTQUEUE_REG_3__4_ <= n13091;
    P2_P2_INSTQUEUE_REG_3__3_ <= n13096;
    P2_P2_INSTQUEUE_REG_3__2_ <= n13101;
    P2_P2_INSTQUEUE_REG_3__1_ <= n13106;
    P2_P2_INSTQUEUE_REG_3__0_ <= n13111;
    P2_P2_INSTQUEUE_REG_2__7_ <= n13116;
    P2_P2_INSTQUEUE_REG_2__6_ <= n13121;
    P2_P2_INSTQUEUE_REG_2__5_ <= n13126;
    P2_P2_INSTQUEUE_REG_2__4_ <= n13131;
    P2_P2_INSTQUEUE_REG_2__3_ <= n13136;
    P2_P2_INSTQUEUE_REG_2__2_ <= n13141;
    P2_P2_INSTQUEUE_REG_2__1_ <= n13146;
    P2_P2_INSTQUEUE_REG_2__0_ <= n13151;
    P2_P2_INSTQUEUE_REG_1__7_ <= n13156;
    P2_P2_INSTQUEUE_REG_1__6_ <= n13161;
    P2_P2_INSTQUEUE_REG_1__5_ <= n13166;
    P2_P2_INSTQUEUE_REG_1__4_ <= n13171;
    P2_P2_INSTQUEUE_REG_1__3_ <= n13176;
    P2_P2_INSTQUEUE_REG_1__2_ <= n13181;
    P2_P2_INSTQUEUE_REG_1__1_ <= n13186;
    P2_P2_INSTQUEUE_REG_1__0_ <= n13191;
    P2_P2_INSTQUEUE_REG_0__7_ <= n13196;
    P2_P2_INSTQUEUE_REG_0__6_ <= n13201;
    P2_P2_INSTQUEUE_REG_0__5_ <= n13206;
    P2_P2_INSTQUEUE_REG_0__4_ <= n13211;
    P2_P2_INSTQUEUE_REG_0__3_ <= n13216;
    P2_P2_INSTQUEUE_REG_0__2_ <= n13221;
    P2_P2_INSTQUEUE_REG_0__1_ <= n13226;
    P2_P2_INSTQUEUE_REG_0__0_ <= n13231;
    P2_P2_INSTQUEUERD_ADDR_REG_4_ <= n13236;
    P2_P2_INSTQUEUERD_ADDR_REG_3_ <= n13241;
    P2_P2_INSTQUEUERD_ADDR_REG_2_ <= n13246;
    P2_P2_INSTQUEUERD_ADDR_REG_1_ <= n13251;
    P2_P2_INSTQUEUERD_ADDR_REG_0_ <= n13256;
    P2_P2_INSTQUEUEWR_ADDR_REG_4_ <= n13261;
    P2_P2_INSTQUEUEWR_ADDR_REG_3_ <= n13266;
    P2_P2_INSTQUEUEWR_ADDR_REG_2_ <= n13271;
    P2_P2_INSTQUEUEWR_ADDR_REG_1_ <= n13276;
    P2_P2_INSTQUEUEWR_ADDR_REG_0_ <= n13281;
    P2_P2_INSTADDRPOINTER_REG_0_ <= n13286;
    P2_P2_INSTADDRPOINTER_REG_1_ <= n13291;
    P2_P2_INSTADDRPOINTER_REG_2_ <= n13296;
    P2_P2_INSTADDRPOINTER_REG_3_ <= n13301;
    P2_P2_INSTADDRPOINTER_REG_4_ <= n13306;
    P2_P2_INSTADDRPOINTER_REG_5_ <= n13311;
    P2_P2_INSTADDRPOINTER_REG_6_ <= n13316;
    P2_P2_INSTADDRPOINTER_REG_7_ <= n13321;
    P2_P2_INSTADDRPOINTER_REG_8_ <= n13326;
    P2_P2_INSTADDRPOINTER_REG_9_ <= n13331;
    P2_P2_INSTADDRPOINTER_REG_10_ <= n13336;
    P2_P2_INSTADDRPOINTER_REG_11_ <= n13341;
    P2_P2_INSTADDRPOINTER_REG_12_ <= n13346;
    P2_P2_INSTADDRPOINTER_REG_13_ <= n13351;
    P2_P2_INSTADDRPOINTER_REG_14_ <= n13356;
    P2_P2_INSTADDRPOINTER_REG_15_ <= n13361;
    P2_P2_INSTADDRPOINTER_REG_16_ <= n13366;
    P2_P2_INSTADDRPOINTER_REG_17_ <= n13371;
    P2_P2_INSTADDRPOINTER_REG_18_ <= n13376;
    P2_P2_INSTADDRPOINTER_REG_19_ <= n13381;
    P2_P2_INSTADDRPOINTER_REG_20_ <= n13386;
    P2_P2_INSTADDRPOINTER_REG_21_ <= n13391;
    P2_P2_INSTADDRPOINTER_REG_22_ <= n13396;
    P2_P2_INSTADDRPOINTER_REG_23_ <= n13401;
    P2_P2_INSTADDRPOINTER_REG_24_ <= n13406;
    P2_P2_INSTADDRPOINTER_REG_25_ <= n13411;
    P2_P2_INSTADDRPOINTER_REG_26_ <= n13416;
    P2_P2_INSTADDRPOINTER_REG_27_ <= n13421;
    P2_P2_INSTADDRPOINTER_REG_28_ <= n13426;
    P2_P2_INSTADDRPOINTER_REG_29_ <= n13431;
    P2_P2_INSTADDRPOINTER_REG_30_ <= n13436;
    P2_P2_INSTADDRPOINTER_REG_31_ <= n13441;
    P2_P2_PHYADDRPOINTER_REG_0_ <= n13446;
    P2_P2_PHYADDRPOINTER_REG_1_ <= n13451;
    P2_P2_PHYADDRPOINTER_REG_2_ <= n13456;
    P2_P2_PHYADDRPOINTER_REG_3_ <= n13461;
    P2_P2_PHYADDRPOINTER_REG_4_ <= n13466;
    P2_P2_PHYADDRPOINTER_REG_5_ <= n13471;
    P2_P2_PHYADDRPOINTER_REG_6_ <= n13476;
    P2_P2_PHYADDRPOINTER_REG_7_ <= n13481;
    P2_P2_PHYADDRPOINTER_REG_8_ <= n13486;
    P2_P2_PHYADDRPOINTER_REG_9_ <= n13491;
    P2_P2_PHYADDRPOINTER_REG_10_ <= n13496;
    P2_P2_PHYADDRPOINTER_REG_11_ <= n13501;
    P2_P2_PHYADDRPOINTER_REG_12_ <= n13506;
    P2_P2_PHYADDRPOINTER_REG_13_ <= n13511;
    P2_P2_PHYADDRPOINTER_REG_14_ <= n13516;
    P2_P2_PHYADDRPOINTER_REG_15_ <= n13521;
    P2_P2_PHYADDRPOINTER_REG_16_ <= n13526;
    P2_P2_PHYADDRPOINTER_REG_17_ <= n13531;
    P2_P2_PHYADDRPOINTER_REG_18_ <= n13536;
    P2_P2_PHYADDRPOINTER_REG_19_ <= n13541;
    P2_P2_PHYADDRPOINTER_REG_20_ <= n13546;
    P2_P2_PHYADDRPOINTER_REG_21_ <= n13551;
    P2_P2_PHYADDRPOINTER_REG_22_ <= n13556;
    P2_P2_PHYADDRPOINTER_REG_23_ <= n13561;
    P2_P2_PHYADDRPOINTER_REG_24_ <= n13566;
    P2_P2_PHYADDRPOINTER_REG_25_ <= n13571;
    P2_P2_PHYADDRPOINTER_REG_26_ <= n13576;
    P2_P2_PHYADDRPOINTER_REG_27_ <= n13581;
    P2_P2_PHYADDRPOINTER_REG_28_ <= n13586;
    P2_P2_PHYADDRPOINTER_REG_29_ <= n13591;
    P2_P2_PHYADDRPOINTER_REG_30_ <= n13596;
    P2_P2_PHYADDRPOINTER_REG_31_ <= n13601;
    P2_P2_LWORD_REG_15_ <= n13606;
    P2_P2_LWORD_REG_14_ <= n13611;
    P2_P2_LWORD_REG_13_ <= n13616;
    P2_P2_LWORD_REG_12_ <= n13621;
    P2_P2_LWORD_REG_11_ <= n13626;
    P2_P2_LWORD_REG_10_ <= n13631;
    P2_P2_LWORD_REG_9_ <= n13636;
    P2_P2_LWORD_REG_8_ <= n13641;
    P2_P2_LWORD_REG_7_ <= n13646;
    P2_P2_LWORD_REG_6_ <= n13651;
    P2_P2_LWORD_REG_5_ <= n13656;
    P2_P2_LWORD_REG_4_ <= n13661;
    P2_P2_LWORD_REG_3_ <= n13666;
    P2_P2_LWORD_REG_2_ <= n13671;
    P2_P2_LWORD_REG_1_ <= n13676;
    P2_P2_LWORD_REG_0_ <= n13681;
    P2_P2_UWORD_REG_14_ <= n13686;
    P2_P2_UWORD_REG_13_ <= n13691;
    P2_P2_UWORD_REG_12_ <= n13696;
    P2_P2_UWORD_REG_11_ <= n13701;
    P2_P2_UWORD_REG_10_ <= n13706;
    P2_P2_UWORD_REG_9_ <= n13711;
    P2_P2_UWORD_REG_8_ <= n13716;
    P2_P2_UWORD_REG_7_ <= n13721;
    P2_P2_UWORD_REG_6_ <= n13726;
    P2_P2_UWORD_REG_5_ <= n13731;
    P2_P2_UWORD_REG_4_ <= n13736;
    P2_P2_UWORD_REG_3_ <= n13741;
    P2_P2_UWORD_REG_2_ <= n13746;
    P2_P2_UWORD_REG_1_ <= n13751;
    P2_P2_UWORD_REG_0_ <= n13756;
    P2_P2_DATAO_REG_0_ <= n13761;
    P2_P2_DATAO_REG_1_ <= n13766;
    P2_P2_DATAO_REG_2_ <= n13771;
    P2_P2_DATAO_REG_3_ <= n13776;
    P2_P2_DATAO_REG_4_ <= n13781;
    P2_P2_DATAO_REG_5_ <= n13786;
    P2_P2_DATAO_REG_6_ <= n13791;
    P2_P2_DATAO_REG_7_ <= n13796;
    P2_P2_DATAO_REG_8_ <= n13801;
    P2_P2_DATAO_REG_9_ <= n13806;
    P2_P2_DATAO_REG_10_ <= n13811;
    P2_P2_DATAO_REG_11_ <= n13816;
    P2_P2_DATAO_REG_12_ <= n13821;
    P2_P2_DATAO_REG_13_ <= n13826;
    P2_P2_DATAO_REG_14_ <= n13831;
    P2_P2_DATAO_REG_15_ <= n13836;
    P2_P2_DATAO_REG_16_ <= n13841;
    P2_P2_DATAO_REG_17_ <= n13846;
    P2_P2_DATAO_REG_18_ <= n13851;
    P2_P2_DATAO_REG_19_ <= n13856;
    P2_P2_DATAO_REG_20_ <= n13861;
    P2_P2_DATAO_REG_21_ <= n13866;
    P2_P2_DATAO_REG_22_ <= n13871;
    P2_P2_DATAO_REG_23_ <= n13876;
    P2_P2_DATAO_REG_24_ <= n13881;
    P2_P2_DATAO_REG_25_ <= n13886;
    P2_P2_DATAO_REG_26_ <= n13891;
    P2_P2_DATAO_REG_27_ <= n13896;
    P2_P2_DATAO_REG_28_ <= n13901;
    P2_P2_DATAO_REG_29_ <= n13906;
    P2_P2_DATAO_REG_30_ <= n13911;
    P2_P2_DATAO_REG_31_ <= n13916;
    P2_P2_EAX_REG_0_ <= n13921;
    P2_P2_EAX_REG_1_ <= n13926;
    P2_P2_EAX_REG_2_ <= n13931;
    P2_P2_EAX_REG_3_ <= n13936;
    P2_P2_EAX_REG_4_ <= n13941;
    P2_P2_EAX_REG_5_ <= n13946;
    P2_P2_EAX_REG_6_ <= n13951;
    P2_P2_EAX_REG_7_ <= n13956;
    P2_P2_EAX_REG_8_ <= n13961;
    P2_P2_EAX_REG_9_ <= n13966;
    P2_P2_EAX_REG_10_ <= n13971;
    P2_P2_EAX_REG_11_ <= n13976;
    P2_P2_EAX_REG_12_ <= n13981;
    P2_P2_EAX_REG_13_ <= n13986;
    P2_P2_EAX_REG_14_ <= n13991;
    P2_P2_EAX_REG_15_ <= n13996;
    P2_P2_EAX_REG_16_ <= n14001;
    P2_P2_EAX_REG_17_ <= n14006;
    P2_P2_EAX_REG_18_ <= n14011;
    P2_P2_EAX_REG_19_ <= n14016;
    P2_P2_EAX_REG_20_ <= n14021;
    P2_P2_EAX_REG_21_ <= n14026;
    P2_P2_EAX_REG_22_ <= n14031;
    P2_P2_EAX_REG_23_ <= n14036;
    P2_P2_EAX_REG_24_ <= n14041;
    P2_P2_EAX_REG_25_ <= n14046;
    P2_P2_EAX_REG_26_ <= n14051;
    P2_P2_EAX_REG_27_ <= n14056;
    P2_P2_EAX_REG_28_ <= n14061;
    P2_P2_EAX_REG_29_ <= n14066;
    P2_P2_EAX_REG_30_ <= n14071;
    P2_P2_EAX_REG_31_ <= n14076;
    P2_P2_EBX_REG_0_ <= n14081;
    P2_P2_EBX_REG_1_ <= n14086;
    P2_P2_EBX_REG_2_ <= n14091;
    P2_P2_EBX_REG_3_ <= n14096;
    P2_P2_EBX_REG_4_ <= n14101;
    P2_P2_EBX_REG_5_ <= n14106;
    P2_P2_EBX_REG_6_ <= n14111;
    P2_P2_EBX_REG_7_ <= n14116;
    P2_P2_EBX_REG_8_ <= n14121;
    P2_P2_EBX_REG_9_ <= n14126;
    P2_P2_EBX_REG_10_ <= n14131;
    P2_P2_EBX_REG_11_ <= n14136;
    P2_P2_EBX_REG_12_ <= n14141;
    P2_P2_EBX_REG_13_ <= n14146;
    P2_P2_EBX_REG_14_ <= n14151;
    P2_P2_EBX_REG_15_ <= n14156;
    P2_P2_EBX_REG_16_ <= n14161;
    P2_P2_EBX_REG_17_ <= n14166;
    P2_P2_EBX_REG_18_ <= n14171;
    P2_P2_EBX_REG_19_ <= n14176;
    P2_P2_EBX_REG_20_ <= n14181;
    P2_P2_EBX_REG_21_ <= n14186;
    P2_P2_EBX_REG_22_ <= n14191;
    P2_P2_EBX_REG_23_ <= n14196;
    P2_P2_EBX_REG_24_ <= n14201;
    P2_P2_EBX_REG_25_ <= n14206;
    P2_P2_EBX_REG_26_ <= n14211;
    P2_P2_EBX_REG_27_ <= n14216;
    P2_P2_EBX_REG_28_ <= n14221;
    P2_P2_EBX_REG_29_ <= n14226;
    P2_P2_EBX_REG_30_ <= n14231;
    P2_P2_EBX_REG_31_ <= n14236;
    P2_P2_REIP_REG_0_ <= n14241;
    P2_P2_REIP_REG_1_ <= n14246;
    P2_P2_REIP_REG_2_ <= n14251;
    P2_P2_REIP_REG_3_ <= n14256;
    P2_P2_REIP_REG_4_ <= n14261;
    P2_P2_REIP_REG_5_ <= n14266;
    P2_P2_REIP_REG_6_ <= n14271;
    P2_P2_REIP_REG_7_ <= n14276;
    P2_P2_REIP_REG_8_ <= n14281;
    P2_P2_REIP_REG_9_ <= n14286;
    P2_P2_REIP_REG_10_ <= n14291;
    P2_P2_REIP_REG_11_ <= n14296;
    P2_P2_REIP_REG_12_ <= n14301;
    P2_P2_REIP_REG_13_ <= n14306;
    P2_P2_REIP_REG_14_ <= n14311;
    P2_P2_REIP_REG_15_ <= n14316;
    P2_P2_REIP_REG_16_ <= n14321;
    P2_P2_REIP_REG_17_ <= n14326;
    P2_P2_REIP_REG_18_ <= n14331;
    P2_P2_REIP_REG_19_ <= n14336;
    P2_P2_REIP_REG_20_ <= n14341;
    P2_P2_REIP_REG_21_ <= n14346;
    P2_P2_REIP_REG_22_ <= n14351;
    P2_P2_REIP_REG_23_ <= n14356;
    P2_P2_REIP_REG_24_ <= n14361;
    P2_P2_REIP_REG_25_ <= n14366;
    P2_P2_REIP_REG_26_ <= n14371;
    P2_P2_REIP_REG_27_ <= n14376;
    P2_P2_REIP_REG_28_ <= n14381;
    P2_P2_REIP_REG_29_ <= n14386;
    P2_P2_REIP_REG_30_ <= n14391;
    P2_P2_REIP_REG_31_ <= n14396;
    P2_P2_BYTEENABLE_REG_3_ <= n14401;
    P2_P2_BYTEENABLE_REG_2_ <= n14406;
    P2_P2_BYTEENABLE_REG_1_ <= n14411;
    P2_P2_BYTEENABLE_REG_0_ <= n14416;
    P2_P2_W_R_N_REG <= n14421;
    P2_P2_FLUSH_REG <= n14426;
    P2_P2_MORE_REG <= n14431;
    P2_P2_STATEBS16_REG <= n14436;
    P2_P2_REQUESTPENDING_REG <= n14441;
    P2_P2_D_C_N_REG <= n14446;
    P2_P2_M_IO_N_REG <= n14451;
    P2_P2_CODEFETCH_REG <= n14456;
    P2_P2_ADS_N_REG <= n14461;
    P2_P2_READREQUEST_REG <= n14466;
    P2_P2_MEMORYFETCH_REG <= n14471;
    P2_P1_BE_N_REG_3_ <= n14476;
    P2_P1_BE_N_REG_2_ <= n14481;
    P2_P1_BE_N_REG_1_ <= n14486;
    P2_P1_BE_N_REG_0_ <= n14491;
    P2_P1_ADDRESS_REG_29_ <= n14496;
    P2_P1_ADDRESS_REG_28_ <= n14501;
    P2_P1_ADDRESS_REG_27_ <= n14506;
    P2_P1_ADDRESS_REG_26_ <= n14511;
    P2_P1_ADDRESS_REG_25_ <= n14516;
    P2_P1_ADDRESS_REG_24_ <= n14521;
    P2_P1_ADDRESS_REG_23_ <= n14526;
    P2_P1_ADDRESS_REG_22_ <= n14531;
    P2_P1_ADDRESS_REG_21_ <= n14536;
    P2_P1_ADDRESS_REG_20_ <= n14541;
    P2_P1_ADDRESS_REG_19_ <= n14546;
    P2_P1_ADDRESS_REG_18_ <= n14551;
    P2_P1_ADDRESS_REG_17_ <= n14556;
    P2_P1_ADDRESS_REG_16_ <= n14561;
    P2_P1_ADDRESS_REG_15_ <= n14566;
    P2_P1_ADDRESS_REG_14_ <= n14571;
    P2_P1_ADDRESS_REG_13_ <= n14576;
    P2_P1_ADDRESS_REG_12_ <= n14581;
    P2_P1_ADDRESS_REG_11_ <= n14586;
    P2_P1_ADDRESS_REG_10_ <= n14591;
    P2_P1_ADDRESS_REG_9_ <= n14596;
    P2_P1_ADDRESS_REG_8_ <= n14601;
    P2_P1_ADDRESS_REG_7_ <= n14606;
    P2_P1_ADDRESS_REG_6_ <= n14611;
    P2_P1_ADDRESS_REG_5_ <= n14616;
    P2_P1_ADDRESS_REG_4_ <= n14621;
    P2_P1_ADDRESS_REG_3_ <= n14626;
    P2_P1_ADDRESS_REG_2_ <= n14631;
    P2_P1_ADDRESS_REG_1_ <= n14636;
    P2_P1_ADDRESS_REG_0_ <= n14641;
    P2_P1_STATE_REG_2_ <= n14646;
    P2_P1_STATE_REG_1_ <= n14651;
    P2_P1_STATE_REG_0_ <= n14656;
    P2_P1_DATAWIDTH_REG_0_ <= n14661;
    P2_P1_DATAWIDTH_REG_1_ <= n14666;
    P2_P1_DATAWIDTH_REG_2_ <= n14671;
    P2_P1_DATAWIDTH_REG_3_ <= n14676;
    P2_P1_DATAWIDTH_REG_4_ <= n14681;
    P2_P1_DATAWIDTH_REG_5_ <= n14686;
    P2_P1_DATAWIDTH_REG_6_ <= n14691;
    P2_P1_DATAWIDTH_REG_7_ <= n14696;
    P2_P1_DATAWIDTH_REG_8_ <= n14701;
    P2_P1_DATAWIDTH_REG_9_ <= n14706;
    P2_P1_DATAWIDTH_REG_10_ <= n14711;
    P2_P1_DATAWIDTH_REG_11_ <= n14716;
    P2_P1_DATAWIDTH_REG_12_ <= n14721;
    P2_P1_DATAWIDTH_REG_13_ <= n14726;
    P2_P1_DATAWIDTH_REG_14_ <= n14731;
    P2_P1_DATAWIDTH_REG_15_ <= n14736;
    P2_P1_DATAWIDTH_REG_16_ <= n14741;
    P2_P1_DATAWIDTH_REG_17_ <= n14746;
    P2_P1_DATAWIDTH_REG_18_ <= n14751;
    P2_P1_DATAWIDTH_REG_19_ <= n14756;
    P2_P1_DATAWIDTH_REG_20_ <= n14761;
    P2_P1_DATAWIDTH_REG_21_ <= n14766;
    P2_P1_DATAWIDTH_REG_22_ <= n14771;
    P2_P1_DATAWIDTH_REG_23_ <= n14776;
    P2_P1_DATAWIDTH_REG_24_ <= n14781;
    P2_P1_DATAWIDTH_REG_25_ <= n14786;
    P2_P1_DATAWIDTH_REG_26_ <= n14791;
    P2_P1_DATAWIDTH_REG_27_ <= n14796;
    P2_P1_DATAWIDTH_REG_28_ <= n14801;
    P2_P1_DATAWIDTH_REG_29_ <= n14806;
    P2_P1_DATAWIDTH_REG_30_ <= n14811;
    P2_P1_DATAWIDTH_REG_31_ <= n14816;
    P2_P1_STATE2_REG_3_ <= n14821;
    P2_P1_STATE2_REG_2_ <= n14826;
    P2_P1_STATE2_REG_1_ <= n14831;
    P2_P1_STATE2_REG_0_ <= n14836;
    P2_P1_INSTQUEUE_REG_15__7_ <= n14841;
    P2_P1_INSTQUEUE_REG_15__6_ <= n14846;
    P2_P1_INSTQUEUE_REG_15__5_ <= n14851;
    P2_P1_INSTQUEUE_REG_15__4_ <= n14856;
    P2_P1_INSTQUEUE_REG_15__3_ <= n14861;
    P2_P1_INSTQUEUE_REG_15__2_ <= n14866;
    P2_P1_INSTQUEUE_REG_15__1_ <= n14871;
    P2_P1_INSTQUEUE_REG_15__0_ <= n14876;
    P2_P1_INSTQUEUE_REG_14__7_ <= n14881;
    P2_P1_INSTQUEUE_REG_14__6_ <= n14886;
    P2_P1_INSTQUEUE_REG_14__5_ <= n14891;
    P2_P1_INSTQUEUE_REG_14__4_ <= n14896;
    P2_P1_INSTQUEUE_REG_14__3_ <= n14901;
    P2_P1_INSTQUEUE_REG_14__2_ <= n14906;
    P2_P1_INSTQUEUE_REG_14__1_ <= n14911;
    P2_P1_INSTQUEUE_REG_14__0_ <= n14916;
    P2_P1_INSTQUEUE_REG_13__7_ <= n14921;
    P2_P1_INSTQUEUE_REG_13__6_ <= n14926;
    P2_P1_INSTQUEUE_REG_13__5_ <= n14931;
    P2_P1_INSTQUEUE_REG_13__4_ <= n14936;
    P2_P1_INSTQUEUE_REG_13__3_ <= n14941;
    P2_P1_INSTQUEUE_REG_13__2_ <= n14946;
    P2_P1_INSTQUEUE_REG_13__1_ <= n14951;
    P2_P1_INSTQUEUE_REG_13__0_ <= n14956;
    P2_P1_INSTQUEUE_REG_12__7_ <= n14961;
    P2_P1_INSTQUEUE_REG_12__6_ <= n14966;
    P2_P1_INSTQUEUE_REG_12__5_ <= n14971;
    P2_P1_INSTQUEUE_REG_12__4_ <= n14976;
    P2_P1_INSTQUEUE_REG_12__3_ <= n14981;
    P2_P1_INSTQUEUE_REG_12__2_ <= n14986;
    P2_P1_INSTQUEUE_REG_12__1_ <= n14991;
    P2_P1_INSTQUEUE_REG_12__0_ <= n14996;
    P2_P1_INSTQUEUE_REG_11__7_ <= n15001;
    P2_P1_INSTQUEUE_REG_11__6_ <= n15006;
    P2_P1_INSTQUEUE_REG_11__5_ <= n15011;
    P2_P1_INSTQUEUE_REG_11__4_ <= n15016;
    P2_P1_INSTQUEUE_REG_11__3_ <= n15021;
    P2_P1_INSTQUEUE_REG_11__2_ <= n15026;
    P2_P1_INSTQUEUE_REG_11__1_ <= n15031;
    P2_P1_INSTQUEUE_REG_11__0_ <= n15036;
    P2_P1_INSTQUEUE_REG_10__7_ <= n15041;
    P2_P1_INSTQUEUE_REG_10__6_ <= n15046;
    P2_P1_INSTQUEUE_REG_10__5_ <= n15051;
    P2_P1_INSTQUEUE_REG_10__4_ <= n15056;
    P2_P1_INSTQUEUE_REG_10__3_ <= n15061;
    P2_P1_INSTQUEUE_REG_10__2_ <= n15066;
    P2_P1_INSTQUEUE_REG_10__1_ <= n15071;
    P2_P1_INSTQUEUE_REG_10__0_ <= n15076;
    P2_P1_INSTQUEUE_REG_9__7_ <= n15081;
    P2_P1_INSTQUEUE_REG_9__6_ <= n15086;
    P2_P1_INSTQUEUE_REG_9__5_ <= n15091;
    P2_P1_INSTQUEUE_REG_9__4_ <= n15096;
    P2_P1_INSTQUEUE_REG_9__3_ <= n15101;
    P2_P1_INSTQUEUE_REG_9__2_ <= n15106;
    P2_P1_INSTQUEUE_REG_9__1_ <= n15111;
    P2_P1_INSTQUEUE_REG_9__0_ <= n15116;
    P2_P1_INSTQUEUE_REG_8__7_ <= n15121;
    P2_P1_INSTQUEUE_REG_8__6_ <= n15126;
    P2_P1_INSTQUEUE_REG_8__5_ <= n15131;
    P2_P1_INSTQUEUE_REG_8__4_ <= n15136;
    P2_P1_INSTQUEUE_REG_8__3_ <= n15141;
    P2_P1_INSTQUEUE_REG_8__2_ <= n15146;
    P2_P1_INSTQUEUE_REG_8__1_ <= n15151;
    P2_P1_INSTQUEUE_REG_8__0_ <= n15156;
    P2_P1_INSTQUEUE_REG_7__7_ <= n15161;
    P2_P1_INSTQUEUE_REG_7__6_ <= n15166;
    P2_P1_INSTQUEUE_REG_7__5_ <= n15171;
    P2_P1_INSTQUEUE_REG_7__4_ <= n15176;
    P2_P1_INSTQUEUE_REG_7__3_ <= n15181;
    P2_P1_INSTQUEUE_REG_7__2_ <= n15186;
    P2_P1_INSTQUEUE_REG_7__1_ <= n15191;
    P2_P1_INSTQUEUE_REG_7__0_ <= n15196;
    P2_P1_INSTQUEUE_REG_6__7_ <= n15201;
    P2_P1_INSTQUEUE_REG_6__6_ <= n15206;
    P2_P1_INSTQUEUE_REG_6__5_ <= n15211;
    P2_P1_INSTQUEUE_REG_6__4_ <= n15216;
    P2_P1_INSTQUEUE_REG_6__3_ <= n15221;
    P2_P1_INSTQUEUE_REG_6__2_ <= n15226;
    P2_P1_INSTQUEUE_REG_6__1_ <= n15231;
    P2_P1_INSTQUEUE_REG_6__0_ <= n15236;
    P2_P1_INSTQUEUE_REG_5__7_ <= n15241;
    P2_P1_INSTQUEUE_REG_5__6_ <= n15246;
    P2_P1_INSTQUEUE_REG_5__5_ <= n15251;
    P2_P1_INSTQUEUE_REG_5__4_ <= n15256;
    P2_P1_INSTQUEUE_REG_5__3_ <= n15261;
    P2_P1_INSTQUEUE_REG_5__2_ <= n15266;
    P2_P1_INSTQUEUE_REG_5__1_ <= n15271;
    P2_P1_INSTQUEUE_REG_5__0_ <= n15276;
    P2_P1_INSTQUEUE_REG_4__7_ <= n15281;
    P2_P1_INSTQUEUE_REG_4__6_ <= n15286;
    P2_P1_INSTQUEUE_REG_4__5_ <= n15291;
    P2_P1_INSTQUEUE_REG_4__4_ <= n15296;
    P2_P1_INSTQUEUE_REG_4__3_ <= n15301;
    P2_P1_INSTQUEUE_REG_4__2_ <= n15306;
    P2_P1_INSTQUEUE_REG_4__1_ <= n15311;
    P2_P1_INSTQUEUE_REG_4__0_ <= n15316;
    P2_P1_INSTQUEUE_REG_3__7_ <= n15321;
    P2_P1_INSTQUEUE_REG_3__6_ <= n15326;
    P2_P1_INSTQUEUE_REG_3__5_ <= n15331;
    P2_P1_INSTQUEUE_REG_3__4_ <= n15336;
    P2_P1_INSTQUEUE_REG_3__3_ <= n15341;
    P2_P1_INSTQUEUE_REG_3__2_ <= n15346;
    P2_P1_INSTQUEUE_REG_3__1_ <= n15351;
    P2_P1_INSTQUEUE_REG_3__0_ <= n15356;
    P2_P1_INSTQUEUE_REG_2__7_ <= n15361;
    P2_P1_INSTQUEUE_REG_2__6_ <= n15366;
    P2_P1_INSTQUEUE_REG_2__5_ <= n15371;
    P2_P1_INSTQUEUE_REG_2__4_ <= n15376;
    P2_P1_INSTQUEUE_REG_2__3_ <= n15381;
    P2_P1_INSTQUEUE_REG_2__2_ <= n15386;
    P2_P1_INSTQUEUE_REG_2__1_ <= n15391;
    P2_P1_INSTQUEUE_REG_2__0_ <= n15396;
    P2_P1_INSTQUEUE_REG_1__7_ <= n15401;
    P2_P1_INSTQUEUE_REG_1__6_ <= n15406;
    P2_P1_INSTQUEUE_REG_1__5_ <= n15411;
    P2_P1_INSTQUEUE_REG_1__4_ <= n15416;
    P2_P1_INSTQUEUE_REG_1__3_ <= n15421;
    P2_P1_INSTQUEUE_REG_1__2_ <= n15426;
    P2_P1_INSTQUEUE_REG_1__1_ <= n15431;
    P2_P1_INSTQUEUE_REG_1__0_ <= n15436;
    P2_P1_INSTQUEUE_REG_0__7_ <= n15441;
    P2_P1_INSTQUEUE_REG_0__6_ <= n15446;
    P2_P1_INSTQUEUE_REG_0__5_ <= n15451;
    P2_P1_INSTQUEUE_REG_0__4_ <= n15456;
    P2_P1_INSTQUEUE_REG_0__3_ <= n15461;
    P2_P1_INSTQUEUE_REG_0__2_ <= n15466;
    P2_P1_INSTQUEUE_REG_0__1_ <= n15471;
    P2_P1_INSTQUEUE_REG_0__0_ <= n15476;
    P2_P1_INSTQUEUERD_ADDR_REG_4_ <= n15481;
    P2_P1_INSTQUEUERD_ADDR_REG_3_ <= n15486;
    P2_P1_INSTQUEUERD_ADDR_REG_2_ <= n15491;
    P2_P1_INSTQUEUERD_ADDR_REG_1_ <= n15496;
    P2_P1_INSTQUEUERD_ADDR_REG_0_ <= n15501;
    P2_P1_INSTQUEUEWR_ADDR_REG_4_ <= n15506;
    P2_P1_INSTQUEUEWR_ADDR_REG_3_ <= n15511;
    P2_P1_INSTQUEUEWR_ADDR_REG_2_ <= n15516;
    P2_P1_INSTQUEUEWR_ADDR_REG_1_ <= n15521;
    P2_P1_INSTQUEUEWR_ADDR_REG_0_ <= n15526;
    P2_P1_INSTADDRPOINTER_REG_0_ <= n15531;
    P2_P1_INSTADDRPOINTER_REG_1_ <= n15536;
    P2_P1_INSTADDRPOINTER_REG_2_ <= n15541;
    P2_P1_INSTADDRPOINTER_REG_3_ <= n15546;
    P2_P1_INSTADDRPOINTER_REG_4_ <= n15551;
    P2_P1_INSTADDRPOINTER_REG_5_ <= n15556;
    P2_P1_INSTADDRPOINTER_REG_6_ <= n15561;
    P2_P1_INSTADDRPOINTER_REG_7_ <= n15566;
    P2_P1_INSTADDRPOINTER_REG_8_ <= n15571;
    P2_P1_INSTADDRPOINTER_REG_9_ <= n15576;
    P2_P1_INSTADDRPOINTER_REG_10_ <= n15581;
    P2_P1_INSTADDRPOINTER_REG_11_ <= n15586;
    P2_P1_INSTADDRPOINTER_REG_12_ <= n15591;
    P2_P1_INSTADDRPOINTER_REG_13_ <= n15596;
    P2_P1_INSTADDRPOINTER_REG_14_ <= n15601;
    P2_P1_INSTADDRPOINTER_REG_15_ <= n15606;
    P2_P1_INSTADDRPOINTER_REG_16_ <= n15611;
    P2_P1_INSTADDRPOINTER_REG_17_ <= n15616;
    P2_P1_INSTADDRPOINTER_REG_18_ <= n15621;
    P2_P1_INSTADDRPOINTER_REG_19_ <= n15626;
    P2_P1_INSTADDRPOINTER_REG_20_ <= n15631;
    P2_P1_INSTADDRPOINTER_REG_21_ <= n15636;
    P2_P1_INSTADDRPOINTER_REG_22_ <= n15641;
    P2_P1_INSTADDRPOINTER_REG_23_ <= n15646;
    P2_P1_INSTADDRPOINTER_REG_24_ <= n15651;
    P2_P1_INSTADDRPOINTER_REG_25_ <= n15656;
    P2_P1_INSTADDRPOINTER_REG_26_ <= n15661;
    P2_P1_INSTADDRPOINTER_REG_27_ <= n15666;
    P2_P1_INSTADDRPOINTER_REG_28_ <= n15671;
    P2_P1_INSTADDRPOINTER_REG_29_ <= n15676;
    P2_P1_INSTADDRPOINTER_REG_30_ <= n15681;
    P2_P1_INSTADDRPOINTER_REG_31_ <= n15686;
    P2_P1_PHYADDRPOINTER_REG_0_ <= n15691;
    P2_P1_PHYADDRPOINTER_REG_1_ <= n15696;
    P2_P1_PHYADDRPOINTER_REG_2_ <= n15701;
    P2_P1_PHYADDRPOINTER_REG_3_ <= n15706;
    P2_P1_PHYADDRPOINTER_REG_4_ <= n15711;
    P2_P1_PHYADDRPOINTER_REG_5_ <= n15716;
    P2_P1_PHYADDRPOINTER_REG_6_ <= n15721;
    P2_P1_PHYADDRPOINTER_REG_7_ <= n15726;
    P2_P1_PHYADDRPOINTER_REG_8_ <= n15731;
    P2_P1_PHYADDRPOINTER_REG_9_ <= n15736;
    P2_P1_PHYADDRPOINTER_REG_10_ <= n15741;
    P2_P1_PHYADDRPOINTER_REG_11_ <= n15746;
    P2_P1_PHYADDRPOINTER_REG_12_ <= n15751;
    P2_P1_PHYADDRPOINTER_REG_13_ <= n15756;
    P2_P1_PHYADDRPOINTER_REG_14_ <= n15761;
    P2_P1_PHYADDRPOINTER_REG_15_ <= n15766;
    P2_P1_PHYADDRPOINTER_REG_16_ <= n15771;
    P2_P1_PHYADDRPOINTER_REG_17_ <= n15776;
    P2_P1_PHYADDRPOINTER_REG_18_ <= n15781;
    P2_P1_PHYADDRPOINTER_REG_19_ <= n15786;
    P2_P1_PHYADDRPOINTER_REG_20_ <= n15791;
    P2_P1_PHYADDRPOINTER_REG_21_ <= n15796;
    P2_P1_PHYADDRPOINTER_REG_22_ <= n15801;
    P2_P1_PHYADDRPOINTER_REG_23_ <= n15806;
    P2_P1_PHYADDRPOINTER_REG_24_ <= n15811;
    P2_P1_PHYADDRPOINTER_REG_25_ <= n15816;
    P2_P1_PHYADDRPOINTER_REG_26_ <= n15821;
    P2_P1_PHYADDRPOINTER_REG_27_ <= n15826;
    P2_P1_PHYADDRPOINTER_REG_28_ <= n15831;
    P2_P1_PHYADDRPOINTER_REG_29_ <= n15836;
    P2_P1_PHYADDRPOINTER_REG_30_ <= n15841;
    P2_P1_PHYADDRPOINTER_REG_31_ <= n15846;
    P2_P1_LWORD_REG_15_ <= n15851;
    P2_P1_LWORD_REG_14_ <= n15856;
    P2_P1_LWORD_REG_13_ <= n15861;
    P2_P1_LWORD_REG_12_ <= n15866;
    P2_P1_LWORD_REG_11_ <= n15871;
    P2_P1_LWORD_REG_10_ <= n15876;
    P2_P1_LWORD_REG_9_ <= n15881;
    P2_P1_LWORD_REG_8_ <= n15886;
    P2_P1_LWORD_REG_7_ <= n15891;
    P2_P1_LWORD_REG_6_ <= n15896;
    P2_P1_LWORD_REG_5_ <= n15901;
    P2_P1_LWORD_REG_4_ <= n15906;
    P2_P1_LWORD_REG_3_ <= n15911;
    P2_P1_LWORD_REG_2_ <= n15916;
    P2_P1_LWORD_REG_1_ <= n15921;
    P2_P1_LWORD_REG_0_ <= n15926;
    P2_P1_UWORD_REG_14_ <= n15931;
    P2_P1_UWORD_REG_13_ <= n15936;
    P2_P1_UWORD_REG_12_ <= n15941;
    P2_P1_UWORD_REG_11_ <= n15946;
    P2_P1_UWORD_REG_10_ <= n15951;
    P2_P1_UWORD_REG_9_ <= n15956;
    P2_P1_UWORD_REG_8_ <= n15961;
    P2_P1_UWORD_REG_7_ <= n15966;
    P2_P1_UWORD_REG_6_ <= n15971;
    P2_P1_UWORD_REG_5_ <= n15976;
    P2_P1_UWORD_REG_4_ <= n15981;
    P2_P1_UWORD_REG_3_ <= n15986;
    P2_P1_UWORD_REG_2_ <= n15991;
    P2_P1_UWORD_REG_1_ <= n15996;
    P2_P1_UWORD_REG_0_ <= n16001;
    P2_P1_DATAO_REG_0_ <= n16006;
    P2_P1_DATAO_REG_1_ <= n16011;
    P2_P1_DATAO_REG_2_ <= n16016;
    P2_P1_DATAO_REG_3_ <= n16021;
    P2_P1_DATAO_REG_4_ <= n16026;
    P2_P1_DATAO_REG_5_ <= n16031;
    P2_P1_DATAO_REG_6_ <= n16036;
    P2_P1_DATAO_REG_7_ <= n16041;
    P2_P1_DATAO_REG_8_ <= n16046;
    P2_P1_DATAO_REG_9_ <= n16051;
    P2_P1_DATAO_REG_10_ <= n16056;
    P2_P1_DATAO_REG_11_ <= n16061;
    P2_P1_DATAO_REG_12_ <= n16066;
    P2_P1_DATAO_REG_13_ <= n16071;
    P2_P1_DATAO_REG_14_ <= n16076;
    P2_P1_DATAO_REG_15_ <= n16081;
    P2_P1_DATAO_REG_16_ <= n16086;
    P2_P1_DATAO_REG_17_ <= n16091;
    P2_P1_DATAO_REG_18_ <= n16096;
    P2_P1_DATAO_REG_19_ <= n16101;
    P2_P1_DATAO_REG_20_ <= n16106;
    P2_P1_DATAO_REG_21_ <= n16111;
    P2_P1_DATAO_REG_22_ <= n16116;
    P2_P1_DATAO_REG_23_ <= n16121;
    P2_P1_DATAO_REG_24_ <= n16126;
    P2_P1_DATAO_REG_25_ <= n16131;
    P2_P1_DATAO_REG_26_ <= n16136;
    P2_P1_DATAO_REG_27_ <= n16141;
    P2_P1_DATAO_REG_28_ <= n16146;
    P2_P1_DATAO_REG_29_ <= n16151;
    P2_P1_DATAO_REG_30_ <= n16156;
    P2_P1_DATAO_REG_31_ <= n16161;
    P2_P1_EAX_REG_0_ <= n16166;
    P2_P1_EAX_REG_1_ <= n16171;
    P2_P1_EAX_REG_2_ <= n16176;
    P2_P1_EAX_REG_3_ <= n16181;
    P2_P1_EAX_REG_4_ <= n16186;
    P2_P1_EAX_REG_5_ <= n16191;
    P2_P1_EAX_REG_6_ <= n16196;
    P2_P1_EAX_REG_7_ <= n16201;
    P2_P1_EAX_REG_8_ <= n16206;
    P2_P1_EAX_REG_9_ <= n16211;
    P2_P1_EAX_REG_10_ <= n16216;
    P2_P1_EAX_REG_11_ <= n16221;
    P2_P1_EAX_REG_12_ <= n16226;
    P2_P1_EAX_REG_13_ <= n16231;
    P2_P1_EAX_REG_14_ <= n16236;
    P2_P1_EAX_REG_15_ <= n16241;
    P2_P1_EAX_REG_16_ <= n16246;
    P2_P1_EAX_REG_17_ <= n16251;
    P2_P1_EAX_REG_18_ <= n16256;
    P2_P1_EAX_REG_19_ <= n16261;
    P2_P1_EAX_REG_20_ <= n16266;
    P2_P1_EAX_REG_21_ <= n16271;
    P2_P1_EAX_REG_22_ <= n16276;
    P2_P1_EAX_REG_23_ <= n16281;
    P2_P1_EAX_REG_24_ <= n16286;
    P2_P1_EAX_REG_25_ <= n16291;
    P2_P1_EAX_REG_26_ <= n16296;
    P2_P1_EAX_REG_27_ <= n16301;
    P2_P1_EAX_REG_28_ <= n16306;
    P2_P1_EAX_REG_29_ <= n16311;
    P2_P1_EAX_REG_30_ <= n16316;
    P2_P1_EAX_REG_31_ <= n16321;
    P2_P1_EBX_REG_0_ <= n16326;
    P2_P1_EBX_REG_1_ <= n16331;
    P2_P1_EBX_REG_2_ <= n16336;
    P2_P1_EBX_REG_3_ <= n16341;
    P2_P1_EBX_REG_4_ <= n16346;
    P2_P1_EBX_REG_5_ <= n16351;
    P2_P1_EBX_REG_6_ <= n16356;
    P2_P1_EBX_REG_7_ <= n16361;
    P2_P1_EBX_REG_8_ <= n16366;
    P2_P1_EBX_REG_9_ <= n16371;
    P2_P1_EBX_REG_10_ <= n16376;
    P2_P1_EBX_REG_11_ <= n16381;
    P2_P1_EBX_REG_12_ <= n16386;
    P2_P1_EBX_REG_13_ <= n16391;
    P2_P1_EBX_REG_14_ <= n16396;
    P2_P1_EBX_REG_15_ <= n16401;
    P2_P1_EBX_REG_16_ <= n16406;
    P2_P1_EBX_REG_17_ <= n16411;
    P2_P1_EBX_REG_18_ <= n16416;
    P2_P1_EBX_REG_19_ <= n16421;
    P2_P1_EBX_REG_20_ <= n16426;
    P2_P1_EBX_REG_21_ <= n16431;
    P2_P1_EBX_REG_22_ <= n16436;
    P2_P1_EBX_REG_23_ <= n16441;
    P2_P1_EBX_REG_24_ <= n16446;
    P2_P1_EBX_REG_25_ <= n16451;
    P2_P1_EBX_REG_26_ <= n16456;
    P2_P1_EBX_REG_27_ <= n16461;
    P2_P1_EBX_REG_28_ <= n16466;
    P2_P1_EBX_REG_29_ <= n16471;
    P2_P1_EBX_REG_30_ <= n16476;
    P2_P1_EBX_REG_31_ <= n16481;
    P2_P1_REIP_REG_0_ <= n16486;
    P2_P1_REIP_REG_1_ <= n16491;
    P2_P1_REIP_REG_2_ <= n16496;
    P2_P1_REIP_REG_3_ <= n16501;
    P2_P1_REIP_REG_4_ <= n16506;
    P2_P1_REIP_REG_5_ <= n16511;
    P2_P1_REIP_REG_6_ <= n16516;
    P2_P1_REIP_REG_7_ <= n16521;
    P2_P1_REIP_REG_8_ <= n16526;
    P2_P1_REIP_REG_9_ <= n16531;
    P2_P1_REIP_REG_10_ <= n16536;
    P2_P1_REIP_REG_11_ <= n16541;
    P2_P1_REIP_REG_12_ <= n16546;
    P2_P1_REIP_REG_13_ <= n16551;
    P2_P1_REIP_REG_14_ <= n16556;
    P2_P1_REIP_REG_15_ <= n16561;
    P2_P1_REIP_REG_16_ <= n16566;
    P2_P1_REIP_REG_17_ <= n16571;
    P2_P1_REIP_REG_18_ <= n16576;
    P2_P1_REIP_REG_19_ <= n16581;
    P2_P1_REIP_REG_20_ <= n16586;
    P2_P1_REIP_REG_21_ <= n16591;
    P2_P1_REIP_REG_22_ <= n16596;
    P2_P1_REIP_REG_23_ <= n16601;
    P2_P1_REIP_REG_24_ <= n16606;
    P2_P1_REIP_REG_25_ <= n16611;
    P2_P1_REIP_REG_26_ <= n16616;
    P2_P1_REIP_REG_27_ <= n16621;
    P2_P1_REIP_REG_28_ <= n16626;
    P2_P1_REIP_REG_29_ <= n16631;
    P2_P1_REIP_REG_30_ <= n16636;
    P2_P1_REIP_REG_31_ <= n16641;
    P2_P1_BYTEENABLE_REG_3_ <= n16646;
    P2_P1_BYTEENABLE_REG_2_ <= n16651;
    P2_P1_BYTEENABLE_REG_1_ <= n16656;
    P2_P1_BYTEENABLE_REG_0_ <= n16661;
    P2_P1_W_R_N_REG <= n16666;
    P2_P1_FLUSH_REG <= n16671;
    P2_P1_MORE_REG <= n16676;
    P2_P1_STATEBS16_REG <= n16681;
    P2_P1_REQUESTPENDING_REG <= n16686;
    P2_P1_D_C_N_REG <= n16691;
    P2_P1_M_IO_N_REG <= n16696;
    P2_P1_CODEFETCH_REG <= n16701;
    P2_P1_ADS_N_REG <= n16706;
    P2_P1_READREQUEST_REG <= n16711;
    P2_P1_MEMORYFETCH_REG <= n16716;
  end
endmodule


