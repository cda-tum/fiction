// Benchmark "top" written by ABC on Mon Feb 19 11:52:43 2024

module top ( 
    pcount_3_, pdata_22_, pdata_35_, pdata_48_, pinreg_1_, poutreg_51_,
    pcount_2_, pdata_10_, pdata_21_, pdata_36_, pdata_47_, pinreg_0_,
    poutreg_52_, poutreg_63_, pcount_1_, pdata_8_, pdata_24_, pdata_37_,
    pdata_46_, pdata_59_, poutreg_40_, poutreg_53_, poutreg_62_, pcount_0_,
    pdata_9_, pdata_23_, pdata_38_, pdata_45_, poutreg_54_, poutreg_61_,
    pdata_6_, pdata_26_, pdata_31_, pdata_44_, pinreg_5_, poutreg_55_,
    pdata_7_, pdata_25_, pdata_32_, pdata_43_, pinreg_4_, poutreg_30_,
    poutreg_56_, pdata_4_, pdata_28_, pdata_33_, pdata_42_, pinreg_3_,
    poutreg_57_, pdata_5_, pdata_27_, pdata_34_, pdata_41_, pinreg_2_,
    poutreg_58_, pd_20_, pdata_17_, pdata_40_, pinreg_9_, poutreg_0_,
    poutreg_33_, poutreg_46_, pc_20_, pd_10_, pdata_18_, pinreg_8_,
    poutreg_1_, poutreg_34_, poutreg_45_, preset_0_, pc_21_, pd_11_,
    pd_22_, pdata_15_, pinreg_7_, poutreg_31_, poutreg_48_, pc_22_, pd_12_,
    pd_21_, pdata_16_, pdata_30_, pinreg_6_, poutreg_32_, poutreg_47_,
    pc_12_, pdata_13_, poutreg_19_, poutreg_37_, poutreg_42_, poutreg_60_,
    pc_11_, pdata_14_, poutreg_38_, poutreg_41_, pc_10_, pdata_11_,
    pdata_20_, poutreg_35_, poutreg_44_, pdata_12_, poutreg_29_,
    poutreg_36_, poutreg_43_, poutreg_50_, pc_9_, pc_16_, pc_27_, pd_8_,
    pd_17_, pdata_in_4_, pinreg_30_, pinreg_41_, pinreg_52_, poutreg_8_,
    poutreg_15_, poutreg_28_, pc_15_, pd_9_, pd_18_, pd_27_, pdata_in_3_,
    pinreg_31_, pinreg_40_, pinreg_53_, poutreg_9_, poutreg_16_,
    poutreg_27_, pc_14_, pd_19_, pdata_60_, pdata_in_6_, pinreg_32_,
    pinreg_43_, pinreg_50_, poutreg_6_, poutreg_17_, poutreg_26_,
    poutreg_39_, pc_13_, pdata_in_5_, pinreg_33_, pinreg_42_, pinreg_51_,
    poutreg_7_, poutreg_18_, poutreg_25_, pc_5_, pc_23_, pd_4_, pd_13_,
    pd_24_, pinreg_12_, pinreg_23_, poutreg_4_, poutreg_11_, poutreg_24_,
    pc_6_, pc_19_, pc_24_, pd_5_, pd_14_, pd_23_, pdata_50_, pdata_in_7_,
    pencrypt_0_, pinreg_13_, pinreg_22_, poutreg_5_, poutreg_12_,
    poutreg_23_, poutreg_49_, pc_7_, pc_18_, pc_25_, pd_6_, pd_15_, pd_26_,
    pdata_19_, pinreg_10_, pinreg_21_, pload_key_0_, poutreg_2_,
    poutreg_13_, poutreg_22_, pc_8_, pc_17_, pc_26_, pd_7_, pd_16_, pd_25_,
    pinreg_11_, pinreg_20_, poutreg_3_, poutreg_14_, poutreg_21_, pc_1_,
    pd_0_, pdata_2_, pdata_53_, pinreg_16_, pinreg_27_, pinreg_38_,
    pinreg_49_, poutreg_20_, poutreg_59_, pc_2_, pd_1_, pdata_3_,
    pdata_29_, pdata_54_, pinreg_17_, pinreg_26_, pinreg_39_, pinreg_48_,
    pc_3_, pd_2_, pdata_0_, pdata_51_, pinreg_14_, pinreg_25_, pc_4_,
    pd_3_, pdata_1_, pdata_52_, pencrypt_mode_0_, pinreg_15_, pinreg_24_,
    poutreg_10_, pdata_39_, pdata_57_, pdata_62_, pdata_in_0_, pinreg_34_,
    pinreg_45_, pdata_58_, pdata_61_, pinreg_35_, pinreg_44_, pdata_55_,
    pdata_in_2_, pinreg_18_, pinreg_29_, pinreg_36_, pinreg_47_,
    pinreg_54_, pc_0_, pdata_49_, pdata_56_, pdata_63_, pdata_in_1_,
    pinreg_19_, pinreg_28_, pinreg_37_, pinreg_46_, pinreg_55_,
    pc_new_6_, pc_new_19_, pd_new_5_, pdata_new_14_, pdata_new_27_,
    pinreg_new_6_, pinreg_new_19_, poutreg_new_9_, pc_new_7_, pd_new_6_,
    pd_new_19_, pdata_new_13_, pdata_new_28_, pdata_new_39_, pinreg_new_5_,
    pinreg_new_18_, poutreg_new_19_, pc_new_4_, pd_new_3_, pdata_new_9_,
    pdata_new_12_, pdata_new_25_, pinreg_new_8_, pinreg_new_17_,
    poutreg_new_7_, pc_new_5_, pd_new_4_, pdata_new_11_, pdata_new_26_,
    pinreg_new_7_, pinreg_new_16_, poutreg_new_8_, pc_new_2_, pd_new_1_,
    pdata_new_10_, pdata_new_36_, pinreg_new_2_, pinreg_new_15_,
    poutreg_new_16_, pc_new_3_, pd_new_2_, pdata_new_35_, pinreg_new_1_,
    pinreg_new_14_, poutreg_new_15_, pc_new_0_, pdata_new_29_,
    pdata_new_38_, pinreg_new_4_, pinreg_new_13_, poutreg_new_18_,
    pc_new_1_, pd_new_0_, pdata_new_37_, pinreg_new_3_, pinreg_new_12_,
    poutreg_new_17_, pc_new_11_, pc_new_22_, pd_new_12_, pd_new_23_,
    pcount_new_0_, pdata_new_3_, pdata_new_45_, pdata_new_58_,
    pinreg_new_22_, pinreg_new_33_, pinreg_new_44_, pinreg_new_55_,
    poutreg_new_1_, poutreg_new_25_, poutreg_new_38_, poutreg_new_61_,
    pc_new_12_, pc_new_21_, pd_new_11_, pd_new_24_, pdata_new_4_,
    pdata_new_46_, pdata_new_57_, pinreg_new_23_, pinreg_new_32_,
    pinreg_new_45_, pinreg_new_54_, poutreg_new_2_, poutreg_new_26_,
    poutreg_new_37_, poutreg_new_62_, pc_new_13_, pc_new_24_, pd_new_14_,
    pd_new_21_, pcount_new_2_, pdata_new_1_, pdata_new_47_, pdata_new_56_,
    pinreg_new_0_, pinreg_new_24_, pinreg_new_35_, pinreg_new_42_,
    pinreg_new_53_, poutreg_new_27_, poutreg_new_36_, poutreg_new_49_,
    poutreg_new_50_, poutreg_new_63_, pc_new_14_, pc_new_23_, pd_new_13_,
    pd_new_22_, pcount_new_1_, pdata_new_2_, pdata_new_48_, pdata_new_55_,
    pinreg_new_25_, pinreg_new_34_, pinreg_new_43_, pinreg_new_52_,
    poutreg_new_0_, poutreg_new_28_, poutreg_new_35_, pc_new_15_,
    pc_new_26_, pd_new_16_, pd_new_27_, pdata_new_7_, pdata_new_49_,
    pinreg_new_26_, pinreg_new_37_, pinreg_new_48_, poutreg_new_5_,
    poutreg_new_29_, poutreg_new_47_, poutreg_new_52_, pc_new_16_,
    pc_new_25_, pd_new_15_, pcount_new_3_, pdata_new_8_, pinreg_new_27_,
    pinreg_new_36_, pinreg_new_49_, poutreg_new_6_, poutreg_new_48_,
    poutreg_new_51_, pc_new_17_, pd_new_18_, pd_new_25_, pdata_new_5_,
    pinreg_new_28_, pinreg_new_39_, pinreg_new_46_, poutreg_new_3_,
    poutreg_new_45_, poutreg_new_54_, pc_new_18_, pc_new_27_, pd_new_17_,
    pd_new_26_, pdata_new_6_, pdata_new_59_, pinreg_new_29_,
    pinreg_new_38_, pinreg_new_47_, poutreg_new_4_, poutreg_new_39_,
    poutreg_new_46_, poutreg_new_53_, poutreg_new_60_, pdata_new_50_,
    pdata_new_63_, poutreg_new_30_, poutreg_new_43_, poutreg_new_56_,
    poutreg_new_44_, poutreg_new_55_, pdata_new_61_, pencrypt_mode_new_0_,
    poutreg_new_41_, poutreg_new_58_, pdata_new_40_, pdata_new_62_,
    poutreg_new_20_, poutreg_new_42_, poutreg_new_57_, pdata_new_41_,
    pdata_new_54_, pinreg_new_40_, pinreg_new_51_, poutreg_new_21_,
    poutreg_new_34_, pd_new_20_, pdata_new_0_, pdata_new_42_,
    pdata_new_53_, pdata_new_60_, pinreg_new_41_, pinreg_new_50_,
    poutreg_new_22_, poutreg_new_33_, poutreg_new_40_, poutreg_new_59_,
    pc_new_20_, pd_new_10_, pdata_new_43_, pdata_new_52_, pinreg_new_20_,
    pinreg_new_31_, poutreg_new_23_, poutreg_new_32_, pc_new_10_,
    pdata_new_44_, pdata_new_51_, pinreg_new_21_, pinreg_new_30_,
    poutreg_new_24_, poutreg_new_31_, pdata_new_32_, pinreg_new_11_,
    poutreg_new_12_, pdata_new_20_, pdata_new_31_, pinreg_new_10_,
    poutreg_new_11_, pdata_new_34_, poutreg_new_14_, pdata_new_19_,
    pdata_new_33_, poutreg_new_13_, pd_new_9_, pdata_new_18_,
    pdata_new_23_, pdata_new_17_, pdata_new_24_, pinreg_new_9_, pc_new_8_,
    pd_new_7_, pdata_new_16_, pdata_new_21_, pdata_new_30_,
    poutreg_new_10_, pc_new_9_, pd_new_8_, pdata_new_15_, pdata_new_22_  );
  input  pcount_3_, pdata_22_, pdata_35_, pdata_48_, pinreg_1_,
    poutreg_51_, pcount_2_, pdata_10_, pdata_21_, pdata_36_, pdata_47_,
    pinreg_0_, poutreg_52_, poutreg_63_, pcount_1_, pdata_8_, pdata_24_,
    pdata_37_, pdata_46_, pdata_59_, poutreg_40_, poutreg_53_, poutreg_62_,
    pcount_0_, pdata_9_, pdata_23_, pdata_38_, pdata_45_, poutreg_54_,
    poutreg_61_, pdata_6_, pdata_26_, pdata_31_, pdata_44_, pinreg_5_,
    poutreg_55_, pdata_7_, pdata_25_, pdata_32_, pdata_43_, pinreg_4_,
    poutreg_30_, poutreg_56_, pdata_4_, pdata_28_, pdata_33_, pdata_42_,
    pinreg_3_, poutreg_57_, pdata_5_, pdata_27_, pdata_34_, pdata_41_,
    pinreg_2_, poutreg_58_, pd_20_, pdata_17_, pdata_40_, pinreg_9_,
    poutreg_0_, poutreg_33_, poutreg_46_, pc_20_, pd_10_, pdata_18_,
    pinreg_8_, poutreg_1_, poutreg_34_, poutreg_45_, preset_0_, pc_21_,
    pd_11_, pd_22_, pdata_15_, pinreg_7_, poutreg_31_, poutreg_48_, pc_22_,
    pd_12_, pd_21_, pdata_16_, pdata_30_, pinreg_6_, poutreg_32_,
    poutreg_47_, pc_12_, pdata_13_, poutreg_19_, poutreg_37_, poutreg_42_,
    poutreg_60_, pc_11_, pdata_14_, poutreg_38_, poutreg_41_, pc_10_,
    pdata_11_, pdata_20_, poutreg_35_, poutreg_44_, pdata_12_, poutreg_29_,
    poutreg_36_, poutreg_43_, poutreg_50_, pc_9_, pc_16_, pc_27_, pd_8_,
    pd_17_, pdata_in_4_, pinreg_30_, pinreg_41_, pinreg_52_, poutreg_8_,
    poutreg_15_, poutreg_28_, pc_15_, pd_9_, pd_18_, pd_27_, pdata_in_3_,
    pinreg_31_, pinreg_40_, pinreg_53_, poutreg_9_, poutreg_16_,
    poutreg_27_, pc_14_, pd_19_, pdata_60_, pdata_in_6_, pinreg_32_,
    pinreg_43_, pinreg_50_, poutreg_6_, poutreg_17_, poutreg_26_,
    poutreg_39_, pc_13_, pdata_in_5_, pinreg_33_, pinreg_42_, pinreg_51_,
    poutreg_7_, poutreg_18_, poutreg_25_, pc_5_, pc_23_, pd_4_, pd_13_,
    pd_24_, pinreg_12_, pinreg_23_, poutreg_4_, poutreg_11_, poutreg_24_,
    pc_6_, pc_19_, pc_24_, pd_5_, pd_14_, pd_23_, pdata_50_, pdata_in_7_,
    pencrypt_0_, pinreg_13_, pinreg_22_, poutreg_5_, poutreg_12_,
    poutreg_23_, poutreg_49_, pc_7_, pc_18_, pc_25_, pd_6_, pd_15_, pd_26_,
    pdata_19_, pinreg_10_, pinreg_21_, pload_key_0_, poutreg_2_,
    poutreg_13_, poutreg_22_, pc_8_, pc_17_, pc_26_, pd_7_, pd_16_, pd_25_,
    pinreg_11_, pinreg_20_, poutreg_3_, poutreg_14_, poutreg_21_, pc_1_,
    pd_0_, pdata_2_, pdata_53_, pinreg_16_, pinreg_27_, pinreg_38_,
    pinreg_49_, poutreg_20_, poutreg_59_, pc_2_, pd_1_, pdata_3_,
    pdata_29_, pdata_54_, pinreg_17_, pinreg_26_, pinreg_39_, pinreg_48_,
    pc_3_, pd_2_, pdata_0_, pdata_51_, pinreg_14_, pinreg_25_, pc_4_,
    pd_3_, pdata_1_, pdata_52_, pencrypt_mode_0_, pinreg_15_, pinreg_24_,
    poutreg_10_, pdata_39_, pdata_57_, pdata_62_, pdata_in_0_, pinreg_34_,
    pinreg_45_, pdata_58_, pdata_61_, pinreg_35_, pinreg_44_, pdata_55_,
    pdata_in_2_, pinreg_18_, pinreg_29_, pinreg_36_, pinreg_47_,
    pinreg_54_, pc_0_, pdata_49_, pdata_56_, pdata_63_, pdata_in_1_,
    pinreg_19_, pinreg_28_, pinreg_37_, pinreg_46_, pinreg_55_;
  output pc_new_6_, pc_new_19_, pd_new_5_, pdata_new_14_, pdata_new_27_,
    pinreg_new_6_, pinreg_new_19_, poutreg_new_9_, pc_new_7_, pd_new_6_,
    pd_new_19_, pdata_new_13_, pdata_new_28_, pdata_new_39_, pinreg_new_5_,
    pinreg_new_18_, poutreg_new_19_, pc_new_4_, pd_new_3_, pdata_new_9_,
    pdata_new_12_, pdata_new_25_, pinreg_new_8_, pinreg_new_17_,
    poutreg_new_7_, pc_new_5_, pd_new_4_, pdata_new_11_, pdata_new_26_,
    pinreg_new_7_, pinreg_new_16_, poutreg_new_8_, pc_new_2_, pd_new_1_,
    pdata_new_10_, pdata_new_36_, pinreg_new_2_, pinreg_new_15_,
    poutreg_new_16_, pc_new_3_, pd_new_2_, pdata_new_35_, pinreg_new_1_,
    pinreg_new_14_, poutreg_new_15_, pc_new_0_, pdata_new_29_,
    pdata_new_38_, pinreg_new_4_, pinreg_new_13_, poutreg_new_18_,
    pc_new_1_, pd_new_0_, pdata_new_37_, pinreg_new_3_, pinreg_new_12_,
    poutreg_new_17_, pc_new_11_, pc_new_22_, pd_new_12_, pd_new_23_,
    pcount_new_0_, pdata_new_3_, pdata_new_45_, pdata_new_58_,
    pinreg_new_22_, pinreg_new_33_, pinreg_new_44_, pinreg_new_55_,
    poutreg_new_1_, poutreg_new_25_, poutreg_new_38_, poutreg_new_61_,
    pc_new_12_, pc_new_21_, pd_new_11_, pd_new_24_, pdata_new_4_,
    pdata_new_46_, pdata_new_57_, pinreg_new_23_, pinreg_new_32_,
    pinreg_new_45_, pinreg_new_54_, poutreg_new_2_, poutreg_new_26_,
    poutreg_new_37_, poutreg_new_62_, pc_new_13_, pc_new_24_, pd_new_14_,
    pd_new_21_, pcount_new_2_, pdata_new_1_, pdata_new_47_, pdata_new_56_,
    pinreg_new_0_, pinreg_new_24_, pinreg_new_35_, pinreg_new_42_,
    pinreg_new_53_, poutreg_new_27_, poutreg_new_36_, poutreg_new_49_,
    poutreg_new_50_, poutreg_new_63_, pc_new_14_, pc_new_23_, pd_new_13_,
    pd_new_22_, pcount_new_1_, pdata_new_2_, pdata_new_48_, pdata_new_55_,
    pinreg_new_25_, pinreg_new_34_, pinreg_new_43_, pinreg_new_52_,
    poutreg_new_0_, poutreg_new_28_, poutreg_new_35_, pc_new_15_,
    pc_new_26_, pd_new_16_, pd_new_27_, pdata_new_7_, pdata_new_49_,
    pinreg_new_26_, pinreg_new_37_, pinreg_new_48_, poutreg_new_5_,
    poutreg_new_29_, poutreg_new_47_, poutreg_new_52_, pc_new_16_,
    pc_new_25_, pd_new_15_, pcount_new_3_, pdata_new_8_, pinreg_new_27_,
    pinreg_new_36_, pinreg_new_49_, poutreg_new_6_, poutreg_new_48_,
    poutreg_new_51_, pc_new_17_, pd_new_18_, pd_new_25_, pdata_new_5_,
    pinreg_new_28_, pinreg_new_39_, pinreg_new_46_, poutreg_new_3_,
    poutreg_new_45_, poutreg_new_54_, pc_new_18_, pc_new_27_, pd_new_17_,
    pd_new_26_, pdata_new_6_, pdata_new_59_, pinreg_new_29_,
    pinreg_new_38_, pinreg_new_47_, poutreg_new_4_, poutreg_new_39_,
    poutreg_new_46_, poutreg_new_53_, poutreg_new_60_, pdata_new_50_,
    pdata_new_63_, poutreg_new_30_, poutreg_new_43_, poutreg_new_56_,
    poutreg_new_44_, poutreg_new_55_, pdata_new_61_, pencrypt_mode_new_0_,
    poutreg_new_41_, poutreg_new_58_, pdata_new_40_, pdata_new_62_,
    poutreg_new_20_, poutreg_new_42_, poutreg_new_57_, pdata_new_41_,
    pdata_new_54_, pinreg_new_40_, pinreg_new_51_, poutreg_new_21_,
    poutreg_new_34_, pd_new_20_, pdata_new_0_, pdata_new_42_,
    pdata_new_53_, pdata_new_60_, pinreg_new_41_, pinreg_new_50_,
    poutreg_new_22_, poutreg_new_33_, poutreg_new_40_, poutreg_new_59_,
    pc_new_20_, pd_new_10_, pdata_new_43_, pdata_new_52_, pinreg_new_20_,
    pinreg_new_31_, poutreg_new_23_, poutreg_new_32_, pc_new_10_,
    pdata_new_44_, pdata_new_51_, pinreg_new_21_, pinreg_new_30_,
    poutreg_new_24_, poutreg_new_31_, pdata_new_32_, pinreg_new_11_,
    poutreg_new_12_, pdata_new_20_, pdata_new_31_, pinreg_new_10_,
    poutreg_new_11_, pdata_new_34_, poutreg_new_14_, pdata_new_19_,
    pdata_new_33_, poutreg_new_13_, pd_new_9_, pdata_new_18_,
    pdata_new_23_, pdata_new_17_, pdata_new_24_, pinreg_new_9_, pc_new_8_,
    pd_new_7_, pdata_new_16_, pdata_new_21_, pdata_new_30_,
    poutreg_new_10_, pc_new_9_, pd_new_8_, pdata_new_15_, pdata_new_22_;
  wire new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n625, new_n626, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1095, new_n1096, new_n1097,
    new_n1098, new_n1099, new_n1100, new_n1101, new_n1102, new_n1103,
    new_n1104, new_n1105, new_n1106, new_n1107, new_n1108, new_n1109,
    new_n1110, new_n1111, new_n1112, new_n1113, new_n1114, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1151, new_n1152, new_n1154,
    new_n1155, new_n1157, new_n1158, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1165, new_n1166, new_n1167, new_n1168, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1288,
    new_n1289, new_n1291, new_n1292, new_n1293, new_n1294, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1362, new_n1363, new_n1365, new_n1366, new_n1367,
    new_n1368, new_n1369, new_n1370, new_n1371, new_n1372, new_n1373,
    new_n1374, new_n1375, new_n1376, new_n1377, new_n1378, new_n1379,
    new_n1380, new_n1381, new_n1382, new_n1383, new_n1384, new_n1385,
    new_n1386, new_n1387, new_n1388, new_n1389, new_n1390, new_n1391,
    new_n1392, new_n1393, new_n1394, new_n1395, new_n1396, new_n1397,
    new_n1398, new_n1399, new_n1400, new_n1401, new_n1402, new_n1403,
    new_n1404, new_n1405, new_n1406, new_n1407, new_n1408, new_n1409,
    new_n1410, new_n1411, new_n1412, new_n1413, new_n1414, new_n1415,
    new_n1416, new_n1417, new_n1418, new_n1419, new_n1420, new_n1421,
    new_n1422, new_n1423, new_n1424, new_n1425, new_n1426, new_n1427,
    new_n1428, new_n1429, new_n1430, new_n1431, new_n1432, new_n1433,
    new_n1434, new_n1435, new_n1436, new_n1437, new_n1438, new_n1439,
    new_n1440, new_n1441, new_n1442, new_n1443, new_n1444, new_n1445,
    new_n1446, new_n1447, new_n1448, new_n1449, new_n1450, new_n1451,
    new_n1452, new_n1453, new_n1454, new_n1455, new_n1456, new_n1457,
    new_n1458, new_n1459, new_n1460, new_n1461, new_n1462, new_n1463,
    new_n1464, new_n1465, new_n1466, new_n1467, new_n1468, new_n1469,
    new_n1470, new_n1471, new_n1472, new_n1473, new_n1474, new_n1475,
    new_n1476, new_n1477, new_n1478, new_n1479, new_n1480, new_n1481,
    new_n1482, new_n1483, new_n1484, new_n1485, new_n1486, new_n1487,
    new_n1488, new_n1489, new_n1490, new_n1491, new_n1492, new_n1493,
    new_n1494, new_n1495, new_n1496, new_n1497, new_n1498, new_n1499,
    new_n1500, new_n1501, new_n1502, new_n1503, new_n1505, new_n1506,
    new_n1507, new_n1508, new_n1510, new_n1511, new_n1512, new_n1513,
    new_n1515, new_n1516, new_n1517, new_n1518, new_n1519, new_n1520,
    new_n1522, new_n1523, new_n1524, new_n1525, new_n1526, new_n1527,
    new_n1528, new_n1529, new_n1530, new_n1531, new_n1532, new_n1533,
    new_n1534, new_n1535, new_n1536, new_n1537, new_n1538, new_n1539,
    new_n1540, new_n1541, new_n1542, new_n1543, new_n1544, new_n1545,
    new_n1546, new_n1547, new_n1549, new_n1550, new_n1551, new_n1552,
    new_n1553, new_n1554, new_n1555, new_n1556, new_n1557, new_n1558,
    new_n1559, new_n1560, new_n1561, new_n1562, new_n1563, new_n1564,
    new_n1565, new_n1566, new_n1567, new_n1568, new_n1569, new_n1570,
    new_n1571, new_n1572, new_n1573, new_n1574, new_n1576, new_n1577,
    new_n1578, new_n1579, new_n1580, new_n1581, new_n1582, new_n1583,
    new_n1584, new_n1585, new_n1586, new_n1587, new_n1588, new_n1589,
    new_n1590, new_n1591, new_n1592, new_n1593, new_n1594, new_n1595,
    new_n1596, new_n1597, new_n1598, new_n1599, new_n1600, new_n1601,
    new_n1602, new_n1603, new_n1604, new_n1605, new_n1606, new_n1607,
    new_n1608, new_n1609, new_n1610, new_n1611, new_n1612, new_n1613,
    new_n1614, new_n1615, new_n1616, new_n1617, new_n1618, new_n1619,
    new_n1620, new_n1621, new_n1622, new_n1623, new_n1624, new_n1625,
    new_n1626, new_n1627, new_n1628, new_n1629, new_n1630, new_n1631,
    new_n1632, new_n1633, new_n1634, new_n1635, new_n1636, new_n1637,
    new_n1638, new_n1639, new_n1640, new_n1641, new_n1642, new_n1643,
    new_n1644, new_n1645, new_n1646, new_n1647, new_n1648, new_n1649,
    new_n1650, new_n1651, new_n1652, new_n1653, new_n1654, new_n1655,
    new_n1656, new_n1657, new_n1658, new_n1659, new_n1660, new_n1661,
    new_n1662, new_n1663, new_n1664, new_n1665, new_n1666, new_n1667,
    new_n1668, new_n1669, new_n1670, new_n1671, new_n1672, new_n1673,
    new_n1674, new_n1675, new_n1676, new_n1677, new_n1678, new_n1679,
    new_n1680, new_n1681, new_n1682, new_n1683, new_n1684, new_n1685,
    new_n1686, new_n1687, new_n1688, new_n1689, new_n1690, new_n1691,
    new_n1692, new_n1693, new_n1694, new_n1695, new_n1696, new_n1697,
    new_n1698, new_n1699, new_n1700, new_n1701, new_n1702, new_n1703,
    new_n1704, new_n1705, new_n1706, new_n1707, new_n1708, new_n1709,
    new_n1710, new_n1711, new_n1712, new_n1713, new_n1714, new_n1715,
    new_n1716, new_n1717, new_n1718, new_n1720, new_n1721, new_n1722,
    new_n1723, new_n1725, new_n1726, new_n1727, new_n1728, new_n1730,
    new_n1731, new_n1732, new_n1733, new_n1734, new_n1735, new_n1736,
    new_n1737, new_n1738, new_n1739, new_n1740, new_n1741, new_n1742,
    new_n1743, new_n1744, new_n1745, new_n1746, new_n1747, new_n1748,
    new_n1749, new_n1750, new_n1751, new_n1752, new_n1753, new_n1754,
    new_n1755, new_n1756, new_n1757, new_n1758, new_n1759, new_n1760,
    new_n1761, new_n1762, new_n1763, new_n1764, new_n1765, new_n1766,
    new_n1767, new_n1768, new_n1769, new_n1770, new_n1771, new_n1772,
    new_n1773, new_n1774, new_n1775, new_n1776, new_n1777, new_n1778,
    new_n1779, new_n1780, new_n1781, new_n1782, new_n1783, new_n1784,
    new_n1785, new_n1786, new_n1787, new_n1788, new_n1789, new_n1790,
    new_n1791, new_n1792, new_n1793, new_n1794, new_n1795, new_n1796,
    new_n1797, new_n1798, new_n1799, new_n1800, new_n1801, new_n1802,
    new_n1803, new_n1804, new_n1805, new_n1806, new_n1807, new_n1808,
    new_n1809, new_n1810, new_n1811, new_n1812, new_n1813, new_n1814,
    new_n1815, new_n1816, new_n1817, new_n1818, new_n1819, new_n1820,
    new_n1821, new_n1822, new_n1823, new_n1824, new_n1825, new_n1826,
    new_n1827, new_n1828, new_n1829, new_n1830, new_n1831, new_n1832,
    new_n1833, new_n1834, new_n1835, new_n1836, new_n1837, new_n1838,
    new_n1839, new_n1840, new_n1841, new_n1842, new_n1843, new_n1844,
    new_n1845, new_n1846, new_n1847, new_n1848, new_n1849, new_n1850,
    new_n1851, new_n1852, new_n1853, new_n1854, new_n1855, new_n1856,
    new_n1857, new_n1858, new_n1859, new_n1860, new_n1861, new_n1862,
    new_n1863, new_n1864, new_n1865, new_n1866, new_n1867, new_n1868,
    new_n1869, new_n1870, new_n1871, new_n1872, new_n1873, new_n1875,
    new_n1876, new_n1877, new_n1878, new_n1879, new_n1880, new_n1881,
    new_n1882, new_n1883, new_n1884, new_n1885, new_n1886, new_n1887,
    new_n1888, new_n1889, new_n1890, new_n1891, new_n1892, new_n1893,
    new_n1894, new_n1895, new_n1896, new_n1897, new_n1898, new_n1899,
    new_n1900, new_n1902, new_n1903, new_n1905, new_n1906, new_n1907,
    new_n1908, new_n1910, new_n1911, new_n1912, new_n1913, new_n1915,
    new_n1916, new_n1917, new_n1918, new_n1920, new_n1921, new_n1922,
    new_n1923, new_n1924, new_n1925, new_n1927, new_n1928, new_n1929,
    new_n1930, new_n1931, new_n1932, new_n1933, new_n1934, new_n1935,
    new_n1936, new_n1937, new_n1938, new_n1939, new_n1940, new_n1941,
    new_n1942, new_n1943, new_n1944, new_n1945, new_n1946, new_n1947,
    new_n1948, new_n1949, new_n1950, new_n1951, new_n1952, new_n1954,
    new_n1955, new_n1956, new_n1957, new_n1958, new_n1959, new_n1960,
    new_n1961, new_n1962, new_n1963, new_n1964, new_n1965, new_n1966,
    new_n1967, new_n1968, new_n1969, new_n1970, new_n1971, new_n1972,
    new_n1973, new_n1974, new_n1975, new_n1976, new_n1977, new_n1978,
    new_n1979, new_n1981, new_n1982, new_n1983, new_n1984, new_n1985,
    new_n1986, new_n1987, new_n1988, new_n1989, new_n1990, new_n1991,
    new_n1992, new_n1993, new_n1994, new_n1995, new_n1996, new_n1997,
    new_n1998, new_n1999, new_n2000, new_n2001, new_n2002, new_n2003,
    new_n2004, new_n2005, new_n2006, new_n2007, new_n2008, new_n2009,
    new_n2010, new_n2011, new_n2012, new_n2013, new_n2014, new_n2015,
    new_n2016, new_n2017, new_n2018, new_n2019, new_n2020, new_n2021,
    new_n2022, new_n2023, new_n2024, new_n2025, new_n2026, new_n2027,
    new_n2028, new_n2029, new_n2030, new_n2031, new_n2032, new_n2033,
    new_n2034, new_n2035, new_n2036, new_n2037, new_n2038, new_n2039,
    new_n2040, new_n2041, new_n2042, new_n2043, new_n2044, new_n2045,
    new_n2046, new_n2047, new_n2048, new_n2049, new_n2050, new_n2051,
    new_n2052, new_n2053, new_n2054, new_n2055, new_n2056, new_n2057,
    new_n2058, new_n2059, new_n2060, new_n2061, new_n2062, new_n2063,
    new_n2064, new_n2065, new_n2066, new_n2067, new_n2068, new_n2069,
    new_n2070, new_n2071, new_n2072, new_n2073, new_n2074, new_n2075,
    new_n2076, new_n2077, new_n2078, new_n2079, new_n2080, new_n2081,
    new_n2082, new_n2083, new_n2084, new_n2085, new_n2086, new_n2087,
    new_n2088, new_n2089, new_n2090, new_n2091, new_n2092, new_n2093,
    new_n2094, new_n2095, new_n2096, new_n2097, new_n2098, new_n2099,
    new_n2100, new_n2101, new_n2102, new_n2103, new_n2104, new_n2105,
    new_n2106, new_n2107, new_n2108, new_n2109, new_n2110, new_n2111,
    new_n2112, new_n2113, new_n2114, new_n2115, new_n2116, new_n2117,
    new_n2118, new_n2119, new_n2120, new_n2121, new_n2122, new_n2123,
    new_n2125, new_n2126, new_n2127, new_n2128, new_n2130, new_n2131,
    new_n2132, new_n2133, new_n2135, new_n2136, new_n2137, new_n2138,
    new_n2139, new_n2140, new_n2141, new_n2142, new_n2144, new_n2145,
    new_n2146, new_n2147, new_n2148, new_n2149, new_n2150, new_n2151,
    new_n2152, new_n2153, new_n2154, new_n2155, new_n2156, new_n2157,
    new_n2158, new_n2159, new_n2160, new_n2161, new_n2162, new_n2163,
    new_n2164, new_n2165, new_n2166, new_n2167, new_n2168, new_n2169,
    new_n2170, new_n2172, new_n2173, new_n2174, new_n2175, new_n2176,
    new_n2177, new_n2178, new_n2179, new_n2180, new_n2181, new_n2182,
    new_n2183, new_n2184, new_n2185, new_n2186, new_n2187, new_n2188,
    new_n2189, new_n2190, new_n2191, new_n2192, new_n2193, new_n2194,
    new_n2195, new_n2196, new_n2197, new_n2198, new_n2199, new_n2200,
    new_n2202, new_n2203, new_n2204, new_n2205, new_n2206, new_n2207,
    new_n2208, new_n2209, new_n2210, new_n2211, new_n2212, new_n2213,
    new_n2214, new_n2215, new_n2216, new_n2217, new_n2218, new_n2219,
    new_n2220, new_n2221, new_n2222, new_n2223, new_n2224, new_n2225,
    new_n2226, new_n2227, new_n2228, new_n2229, new_n2231, new_n2232,
    new_n2233, new_n2234, new_n2235, new_n2236, new_n2237, new_n2238,
    new_n2239, new_n2240, new_n2241, new_n2242, new_n2243, new_n2244,
    new_n2245, new_n2246, new_n2247, new_n2248, new_n2249, new_n2250,
    new_n2251, new_n2252, new_n2253, new_n2254, new_n2255, new_n2256,
    new_n2257, new_n2258, new_n2260, new_n2262, new_n2263, new_n2265,
    new_n2266, new_n2267, new_n2268, new_n2270, new_n2271, new_n2272,
    new_n2273, new_n2274, new_n2275, new_n2276, new_n2277, new_n2278,
    new_n2279, new_n2280, new_n2281, new_n2282, new_n2283, new_n2284,
    new_n2285, new_n2286, new_n2287, new_n2288, new_n2289, new_n2290,
    new_n2291, new_n2292, new_n2293, new_n2294, new_n2295, new_n2296,
    new_n2297, new_n2298, new_n2299, new_n2300, new_n2301, new_n2302,
    new_n2303, new_n2304, new_n2305, new_n2306, new_n2307, new_n2308,
    new_n2309, new_n2310, new_n2311, new_n2312, new_n2313, new_n2314,
    new_n2315, new_n2316, new_n2317, new_n2318, new_n2319, new_n2320,
    new_n2321, new_n2322, new_n2323, new_n2324, new_n2325, new_n2326,
    new_n2327, new_n2328, new_n2329, new_n2331, new_n2332, new_n2333,
    new_n2334, new_n2336, new_n2337, new_n2338, new_n2339, new_n2341,
    new_n2342, new_n2343, new_n2344, new_n2346, new_n2347, new_n2348,
    new_n2349, new_n2351, new_n2352, new_n2353, new_n2354, new_n2355,
    new_n2356, new_n2357, new_n2358, new_n2360, new_n2361, new_n2362,
    new_n2363, new_n2364, new_n2365, new_n2366, new_n2367, new_n2369,
    new_n2370, new_n2371, new_n2372, new_n2373, new_n2374, new_n2376,
    new_n2377, new_n2378, new_n2379, new_n2380, new_n2381, new_n2382,
    new_n2383, new_n2384, new_n2385, new_n2386, new_n2387, new_n2388,
    new_n2389, new_n2390, new_n2391, new_n2392, new_n2393, new_n2394,
    new_n2395, new_n2396, new_n2397, new_n2398, new_n2399, new_n2400,
    new_n2401, new_n2402, new_n2403, new_n2404, new_n2405, new_n2406,
    new_n2407, new_n2408, new_n2409, new_n2410, new_n2411, new_n2412,
    new_n2413, new_n2414, new_n2415, new_n2416, new_n2417, new_n2418,
    new_n2419, new_n2420, new_n2421, new_n2422, new_n2423, new_n2424,
    new_n2425, new_n2426, new_n2427, new_n2428, new_n2429, new_n2430,
    new_n2431, new_n2432, new_n2433, new_n2435, new_n2436, new_n2437,
    new_n2438, new_n2439, new_n2440, new_n2441, new_n2442, new_n2443,
    new_n2444, new_n2445, new_n2446, new_n2447, new_n2448, new_n2449,
    new_n2450, new_n2451, new_n2452, new_n2453, new_n2454, new_n2455,
    new_n2456, new_n2457, new_n2458, new_n2459, new_n2460, new_n2461,
    new_n2462, new_n2464, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2492, new_n2493,
    new_n2494, new_n2495, new_n2496, new_n2497, new_n2498, new_n2499,
    new_n2500, new_n2501, new_n2502, new_n2503, new_n2504, new_n2505,
    new_n2506, new_n2507, new_n2508, new_n2509, new_n2510, new_n2511,
    new_n2512, new_n2513, new_n2514, new_n2515, new_n2516, new_n2517,
    new_n2518, new_n2519, new_n2521, new_n2522, new_n2523, new_n2524,
    new_n2525, new_n2526, new_n2527, new_n2528, new_n2529, new_n2530,
    new_n2531, new_n2532, new_n2533, new_n2534, new_n2535, new_n2536,
    new_n2537, new_n2538, new_n2539, new_n2540, new_n2541, new_n2542,
    new_n2543, new_n2544, new_n2545, new_n2546, new_n2547, new_n2549,
    new_n2550, new_n2552, new_n2553, new_n2554, new_n2555, new_n2556,
    new_n2557, new_n2558, new_n2559, new_n2560, new_n2561, new_n2562,
    new_n2563, new_n2564, new_n2565, new_n2566, new_n2567, new_n2568,
    new_n2569, new_n2570, new_n2571, new_n2572, new_n2573, new_n2574,
    new_n2575, new_n2576, new_n2577, new_n2578, new_n2579, new_n2580,
    new_n2581, new_n2582, new_n2583, new_n2584, new_n2585, new_n2586,
    new_n2587, new_n2588, new_n2589, new_n2590, new_n2591, new_n2592,
    new_n2593, new_n2594, new_n2596, new_n2597, new_n2598, new_n2599,
    new_n2600, new_n2601, new_n2602, new_n2603, new_n2604, new_n2605,
    new_n2606, new_n2607, new_n2608, new_n2609, new_n2610, new_n2611,
    new_n2612, new_n2613, new_n2614, new_n2615, new_n2616, new_n2617,
    new_n2618, new_n2619, new_n2620, new_n2621, new_n2622, new_n2623,
    new_n2624, new_n2625, new_n2626, new_n2627, new_n2628, new_n2629,
    new_n2630, new_n2631, new_n2632, new_n2633, new_n2634, new_n2635,
    new_n2636, new_n2637, new_n2638, new_n2639, new_n2640, new_n2641,
    new_n2642, new_n2643, new_n2644, new_n2645, new_n2646, new_n2647,
    new_n2648, new_n2649, new_n2650, new_n2651, new_n2652, new_n2653,
    new_n2654, new_n2655, new_n2656, new_n2657, new_n2658, new_n2659,
    new_n2660, new_n2661, new_n2662, new_n2663, new_n2664, new_n2665,
    new_n2666, new_n2667, new_n2668, new_n2669, new_n2670, new_n2671,
    new_n2672, new_n2673, new_n2674, new_n2675, new_n2676, new_n2677,
    new_n2678, new_n2679, new_n2680, new_n2681, new_n2682, new_n2683,
    new_n2684, new_n2685, new_n2686, new_n2687, new_n2688, new_n2689,
    new_n2690, new_n2691, new_n2692, new_n2693, new_n2694, new_n2695,
    new_n2696, new_n2697, new_n2698, new_n2699, new_n2700, new_n2701,
    new_n2702, new_n2703, new_n2704, new_n2705, new_n2706, new_n2707,
    new_n2708, new_n2709, new_n2710, new_n2711, new_n2712, new_n2713,
    new_n2714, new_n2715, new_n2716, new_n2717, new_n2718, new_n2719,
    new_n2720, new_n2721, new_n2722, new_n2723, new_n2724, new_n2725,
    new_n2726, new_n2727, new_n2728, new_n2729, new_n2730, new_n2731,
    new_n2732, new_n2734, new_n2735, new_n2736, new_n2737, new_n2739,
    new_n2740, new_n2741, new_n2742, new_n2744, new_n2745, new_n2746,
    new_n2747, new_n2749, new_n2750, new_n2751, new_n2752, new_n2754,
    new_n2755, new_n2756, new_n2757, new_n2758, new_n2759, new_n2761,
    new_n2762, new_n2763, new_n2764, new_n2765, new_n2766, new_n2768,
    new_n2769, new_n2770, new_n2771, new_n2772, new_n2773, new_n2774,
    new_n2775, new_n2776, new_n2777, new_n2778, new_n2779, new_n2780,
    new_n2781, new_n2782, new_n2783, new_n2784, new_n2785, new_n2786,
    new_n2787, new_n2788, new_n2789, new_n2790, new_n2791, new_n2792,
    new_n2793, new_n2794, new_n2795, new_n2796, new_n2797, new_n2798,
    new_n2799, new_n2800, new_n2801, new_n2802, new_n2803, new_n2804,
    new_n2805, new_n2806, new_n2807, new_n2808, new_n2809, new_n2810,
    new_n2811, new_n2812, new_n2813, new_n2814, new_n2815, new_n2816,
    new_n2817, new_n2818, new_n2819, new_n2820, new_n2821, new_n2822,
    new_n2823, new_n2824, new_n2825, new_n2826, new_n2827, new_n2828,
    new_n2829, new_n2830, new_n2831, new_n2832, new_n2833, new_n2835,
    new_n2836, new_n2837, new_n2839, new_n2840, new_n2841, new_n2842,
    new_n2843, new_n2844, new_n2845, new_n2846, new_n2847, new_n2848,
    new_n2849, new_n2850, new_n2851, new_n2852, new_n2853, new_n2854,
    new_n2855, new_n2856, new_n2857, new_n2858, new_n2859, new_n2860,
    new_n2861, new_n2862, new_n2863, new_n2864, new_n2865, new_n2867,
    new_n2868, new_n2869, new_n2870, new_n2871, new_n2872, new_n2873,
    new_n2874, new_n2875, new_n2876, new_n2877, new_n2878, new_n2879,
    new_n2880, new_n2881, new_n2882, new_n2883, new_n2884, new_n2885,
    new_n2886, new_n2887, new_n2888, new_n2889, new_n2890, new_n2891,
    new_n2892, new_n2894, new_n2895, new_n2896, new_n2897, new_n2898,
    new_n2899, new_n2900, new_n2901, new_n2902, new_n2903, new_n2904,
    new_n2905, new_n2906, new_n2907, new_n2908, new_n2909, new_n2910,
    new_n2911, new_n2912, new_n2913, new_n2914, new_n2915, new_n2916,
    new_n2917, new_n2918, new_n2919, new_n2920, new_n2921, new_n2923,
    new_n2924, new_n2925, new_n2926, new_n2927, new_n2928, new_n2929,
    new_n2930, new_n2931, new_n2932, new_n2933, new_n2934, new_n2935,
    new_n2936, new_n2937, new_n2938, new_n2939, new_n2940, new_n2941,
    new_n2942, new_n2943, new_n2944, new_n2945, new_n2946, new_n2947,
    new_n2948, new_n2950, new_n2951, new_n2952, new_n2953, new_n2954,
    new_n2955, new_n2956, new_n2957, new_n2958, new_n2959, new_n2961,
    new_n2962, new_n2964, new_n2965, new_n2966, new_n2967, new_n2968,
    new_n2969, new_n2970, new_n2971, new_n2972, new_n2973, new_n2974,
    new_n2975, new_n2976, new_n2977, new_n2978, new_n2979, new_n2980,
    new_n2981, new_n2982, new_n2983, new_n2984, new_n2985, new_n2986,
    new_n2987, new_n2988, new_n2989, new_n2990, new_n2991, new_n2992,
    new_n2993, new_n2994, new_n2995, new_n2996, new_n2997, new_n2998,
    new_n2999, new_n3000, new_n3001, new_n3002, new_n3003, new_n3004,
    new_n3005, new_n3006, new_n3007, new_n3008, new_n3009, new_n3010,
    new_n3011, new_n3012, new_n3013, new_n3014, new_n3015, new_n3016,
    new_n3017, new_n3019, new_n3020, new_n3021, new_n3022, new_n3023,
    new_n3024, new_n3025, new_n3026, new_n3027, new_n3028, new_n3029,
    new_n3030, new_n3031, new_n3032, new_n3033, new_n3034, new_n3035,
    new_n3036, new_n3037, new_n3038, new_n3039, new_n3040, new_n3041,
    new_n3042, new_n3043, new_n3044, new_n3045, new_n3046, new_n3047,
    new_n3048, new_n3049, new_n3050, new_n3051, new_n3052, new_n3053,
    new_n3054, new_n3055, new_n3056, new_n3057, new_n3058, new_n3059,
    new_n3060, new_n3061, new_n3063, new_n3064, new_n3065, new_n3066,
    new_n3068, new_n3069, new_n3070, new_n3071, new_n3073, new_n3074,
    new_n3075, new_n3076, new_n3078, new_n3079, new_n3080, new_n3081,
    new_n3083, new_n3084, new_n3085, new_n3086, new_n3088, new_n3089,
    new_n3090, new_n3091, new_n3092, new_n3093, new_n3094, new_n3095,
    new_n3096, new_n3097, new_n3098, new_n3099, new_n3100, new_n3101,
    new_n3102, new_n3103, new_n3104, new_n3105, new_n3106, new_n3107,
    new_n3108, new_n3109, new_n3110, new_n3111, new_n3112, new_n3113,
    new_n3114, new_n3115, new_n3116, new_n3117, new_n3118, new_n3119,
    new_n3120, new_n3121, new_n3122, new_n3123, new_n3124, new_n3125,
    new_n3126, new_n3127, new_n3128, new_n3129, new_n3130, new_n3131,
    new_n3132, new_n3133, new_n3134, new_n3135, new_n3136, new_n3137,
    new_n3138, new_n3139, new_n3140, new_n3141, new_n3142, new_n3143,
    new_n3144, new_n3145, new_n3146, new_n3147, new_n3148, new_n3149,
    new_n3150, new_n3151, new_n3152, new_n3153, new_n3154, new_n3155,
    new_n3156, new_n3157, new_n3158, new_n3159, new_n3160, new_n3161,
    new_n3162, new_n3163, new_n3164, new_n3165, new_n3166, new_n3167,
    new_n3168, new_n3169, new_n3170, new_n3171, new_n3172, new_n3173,
    new_n3174, new_n3175, new_n3176, new_n3177, new_n3178, new_n3179,
    new_n3180, new_n3181, new_n3182, new_n3183, new_n3184, new_n3185,
    new_n3186, new_n3187, new_n3188, new_n3189, new_n3190, new_n3191,
    new_n3192, new_n3193, new_n3194, new_n3195, new_n3196, new_n3197,
    new_n3198, new_n3199, new_n3200, new_n3201, new_n3202, new_n3203,
    new_n3204, new_n3205, new_n3206, new_n3207, new_n3208, new_n3209,
    new_n3210, new_n3211, new_n3212, new_n3213, new_n3214, new_n3215,
    new_n3216, new_n3217, new_n3218, new_n3219, new_n3220, new_n3221,
    new_n3222, new_n3223, new_n3224, new_n3225, new_n3226, new_n3227,
    new_n3228, new_n3229, new_n3230, new_n3231, new_n3232, new_n3233,
    new_n3235, new_n3236, new_n3237, new_n3238, new_n3239, new_n3240,
    new_n3242, new_n3243, new_n3244, new_n3245, new_n3246, new_n3247,
    new_n3248, new_n3249, new_n3250, new_n3251, new_n3252, new_n3253,
    new_n3254, new_n3255, new_n3256, new_n3257, new_n3258, new_n3259,
    new_n3260, new_n3261, new_n3262, new_n3263, new_n3264, new_n3265,
    new_n3266, new_n3267, new_n3268, new_n3269, new_n3270, new_n3271,
    new_n3272, new_n3273, new_n3274, new_n3275, new_n3276, new_n3277,
    new_n3278, new_n3279, new_n3280, new_n3281, new_n3282, new_n3283,
    new_n3284, new_n3285, new_n3286, new_n3287, new_n3288, new_n3289,
    new_n3290, new_n3291, new_n3292, new_n3293, new_n3294, new_n3295,
    new_n3296, new_n3297, new_n3298, new_n3299, new_n3300, new_n3301,
    new_n3302, new_n3304, new_n3305, new_n3306, new_n3307, new_n3308,
    new_n3309, new_n3311, new_n3312, new_n3313, new_n3314, new_n3315,
    new_n3317, new_n3318, new_n3319, new_n3320, new_n3321, new_n3322,
    new_n3323, new_n3324, new_n3325, new_n3326, new_n3327, new_n3328,
    new_n3329, new_n3330, new_n3331, new_n3332, new_n3333, new_n3334,
    new_n3335, new_n3336, new_n3337, new_n3338, new_n3339, new_n3340,
    new_n3341, new_n3342, new_n3343, new_n3344, new_n3346, new_n3347,
    new_n3348, new_n3349, new_n3350, new_n3351, new_n3352, new_n3353,
    new_n3354, new_n3355, new_n3356, new_n3357, new_n3358, new_n3359,
    new_n3360, new_n3361, new_n3362, new_n3363, new_n3364, new_n3365,
    new_n3366, new_n3367, new_n3368, new_n3369, new_n3370, new_n3371,
    new_n3373, new_n3374, new_n3375, new_n3376, new_n3377, new_n3378,
    new_n3379, new_n3380, new_n3381, new_n3382, new_n3383, new_n3384,
    new_n3385, new_n3386, new_n3387, new_n3388, new_n3389, new_n3390,
    new_n3391, new_n3392, new_n3393, new_n3394, new_n3395, new_n3396,
    new_n3397, new_n3398, new_n3399, new_n3401, new_n3402, new_n3403,
    new_n3404, new_n3405, new_n3406, new_n3407, new_n3408, new_n3409,
    new_n3410, new_n3411, new_n3412, new_n3413, new_n3414, new_n3415,
    new_n3416, new_n3417, new_n3418, new_n3419, new_n3420, new_n3421,
    new_n3422, new_n3423, new_n3424, new_n3425, new_n3426, new_n3427,
    new_n3429, new_n3430, new_n3431, new_n3432, new_n3433, new_n3435,
    new_n3436, new_n3438, new_n3439, new_n3440, new_n3441, new_n3443,
    new_n3444, new_n3445, new_n3446, new_n3447, new_n3448, new_n3449,
    new_n3450, new_n3451, new_n3452, new_n3453, new_n3454, new_n3455,
    new_n3456, new_n3457, new_n3458, new_n3459, new_n3460, new_n3461,
    new_n3462, new_n3463, new_n3464, new_n3465, new_n3466, new_n3467,
    new_n3468, new_n3469, new_n3470, new_n3471, new_n3472, new_n3473,
    new_n3474, new_n3475, new_n3476, new_n3477, new_n3478, new_n3479,
    new_n3480, new_n3481, new_n3482, new_n3483, new_n3485, new_n3486,
    new_n3487, new_n3488, new_n3490, new_n3491, new_n3492, new_n3493,
    new_n3495, new_n3496, new_n3497, new_n3498, new_n3500, new_n3501,
    new_n3502, new_n3503, new_n3505, new_n3506, new_n3507, new_n3508,
    new_n3509, new_n3510, new_n3512, new_n3513, new_n3514, new_n3515,
    new_n3516, new_n3517, new_n3519, new_n3520, new_n3521, new_n3522,
    new_n3523, new_n3524, new_n3525, new_n3526, new_n3527, new_n3528,
    new_n3529, new_n3530, new_n3531, new_n3532, new_n3533, new_n3534,
    new_n3535, new_n3536, new_n3537, new_n3538, new_n3539, new_n3540,
    new_n3541, new_n3542, new_n3543, new_n3544, new_n3545, new_n3546,
    new_n3547, new_n3548, new_n3549, new_n3550, new_n3551, new_n3552,
    new_n3553, new_n3554, new_n3555, new_n3556, new_n3557, new_n3558,
    new_n3559, new_n3560, new_n3561, new_n3562, new_n3563, new_n3564,
    new_n3565, new_n3566, new_n3567, new_n3569, new_n3570, new_n3571,
    new_n3572, new_n3573, new_n3574, new_n3575, new_n3576, new_n3577,
    new_n3578, new_n3579, new_n3580, new_n3581, new_n3582, new_n3583,
    new_n3584, new_n3585, new_n3586, new_n3587, new_n3588, new_n3589,
    new_n3590, new_n3591, new_n3592, new_n3593, new_n3595, new_n3596,
    new_n3597, new_n3598, new_n3599, new_n3600, new_n3601, new_n3602,
    new_n3603, new_n3604, new_n3605, new_n3606, new_n3607, new_n3608,
    new_n3609, new_n3610, new_n3611, new_n3612, new_n3613, new_n3614,
    new_n3615, new_n3616, new_n3617, new_n3618, new_n3620, new_n3621,
    new_n3622, new_n3623, new_n3624, new_n3625, new_n3626, new_n3627,
    new_n3628, new_n3629, new_n3630, new_n3631, new_n3632, new_n3633,
    new_n3634, new_n3635, new_n3636, new_n3637, new_n3638, new_n3639,
    new_n3640, new_n3641, new_n3642, new_n3643, new_n3644, new_n3645,
    new_n3647, new_n3648, new_n3649, new_n3650, new_n3651, new_n3652,
    new_n3653, new_n3654, new_n3655, new_n3656, new_n3657, new_n3658,
    new_n3659, new_n3660, new_n3661, new_n3662, new_n3663, new_n3664,
    new_n3665, new_n3666, new_n3667, new_n3668, new_n3669, new_n3670,
    new_n3671, new_n3672, new_n3674, new_n3675, new_n3677, new_n3678,
    new_n3679, new_n3680, new_n3681, new_n3682, new_n3683, new_n3684,
    new_n3685, new_n3686, new_n3687, new_n3688, new_n3689, new_n3690,
    new_n3691, new_n3692, new_n3693, new_n3694, new_n3695, new_n3696,
    new_n3697, new_n3698, new_n3699, new_n3700, new_n3701, new_n3702,
    new_n3703, new_n3704, new_n3705, new_n3706, new_n3707, new_n3708,
    new_n3709, new_n3710, new_n3711, new_n3712, new_n3713, new_n3714,
    new_n3715, new_n3716, new_n3717, new_n3718, new_n3719, new_n3720,
    new_n3722, new_n3723, new_n3724, new_n3725, new_n3727, new_n3728,
    new_n3729, new_n3730, new_n3732, new_n3733, new_n3734, new_n3735,
    new_n3737, new_n3738, new_n3739, new_n3740, new_n3741, new_n3742,
    new_n3743, new_n3744, new_n3746, new_n3747, new_n3748, new_n3749,
    new_n3750, new_n3751, new_n3752, new_n3753, new_n3754, new_n3755,
    new_n3756, new_n3757, new_n3758, new_n3759, new_n3760, new_n3761,
    new_n3762, new_n3763, new_n3764, new_n3765, new_n3766, new_n3767,
    new_n3768, new_n3769, new_n3770, new_n3771, new_n3772, new_n3773,
    new_n3774, new_n3775, new_n3776, new_n3777, new_n3778, new_n3779,
    new_n3780, new_n3781, new_n3782, new_n3783, new_n3784, new_n3785,
    new_n3786, new_n3787, new_n3789, new_n3790, new_n3791, new_n3792,
    new_n3793, new_n3794, new_n3795, new_n3796, new_n3798, new_n3799,
    new_n3800, new_n3801, new_n3802, new_n3803, new_n3805, new_n3806,
    new_n3807, new_n3808, new_n3809, new_n3810, new_n3811, new_n3812,
    new_n3813, new_n3814, new_n3815, new_n3816, new_n3817, new_n3818,
    new_n3819, new_n3820, new_n3821, new_n3822, new_n3823, new_n3824,
    new_n3825, new_n3826, new_n3827, new_n3828, new_n3829, new_n3830,
    new_n3832, new_n3833, new_n3834, new_n3835, new_n3836, new_n3837,
    new_n3838, new_n3839, new_n3840, new_n3841, new_n3842, new_n3843,
    new_n3844, new_n3845, new_n3846, new_n3847, new_n3848, new_n3849,
    new_n3850, new_n3851, new_n3852, new_n3853, new_n3854, new_n3855,
    new_n3856, new_n3858, new_n3859, new_n3860, new_n3861, new_n3862,
    new_n3863, new_n3864, new_n3865, new_n3866, new_n3867, new_n3868,
    new_n3869, new_n3870, new_n3871, new_n3872, new_n3873, new_n3874,
    new_n3875, new_n3876, new_n3877, new_n3878, new_n3879, new_n3880,
    new_n3881, new_n3882, new_n3884, new_n3885, new_n3886, new_n3887,
    new_n3888, new_n3889, new_n3890, new_n3891, new_n3892, new_n3893,
    new_n3894, new_n3895, new_n3896, new_n3897, new_n3899, new_n3900,
    new_n3902, new_n3903, new_n3904, new_n3905, new_n3907, new_n3908,
    new_n3909, new_n3910, new_n3912, new_n3913, new_n3914, new_n3915,
    new_n3917, new_n3918, new_n3919, new_n3920, new_n3921, new_n3922,
    new_n3924, new_n3925, new_n3926, new_n3927, new_n3928, new_n3929,
    new_n3931, new_n3932, new_n3933, new_n3934, new_n3935, new_n3936,
    new_n3937, new_n3938, new_n3939, new_n3940, new_n3941, new_n3942,
    new_n3943, new_n3944, new_n3945, new_n3946, new_n3947, new_n3948,
    new_n3949, new_n3950, new_n3951, new_n3952, new_n3953, new_n3954,
    new_n3955, new_n3956, new_n3957, new_n3958, new_n3959, new_n3960,
    new_n3961, new_n3962, new_n3963, new_n3964, new_n3965, new_n3966,
    new_n3967, new_n3968, new_n3969, new_n3970, new_n3971, new_n3972,
    new_n3973, new_n3974, new_n3975, new_n3976, new_n3977, new_n3978,
    new_n3980, new_n3981, new_n3982, new_n3983, new_n3984, new_n3985,
    new_n3986, new_n3987, new_n3988, new_n3989, new_n3990, new_n3991,
    new_n3992, new_n3993, new_n3994, new_n3995, new_n3996, new_n3997,
    new_n3998, new_n3999, new_n4000, new_n4001, new_n4002, new_n4003,
    new_n4005, new_n4006, new_n4007, new_n4008, new_n4009, new_n4010,
    new_n4011, new_n4012, new_n4013, new_n4014, new_n4015, new_n4016,
    new_n4017, new_n4018, new_n4019, new_n4020, new_n4021, new_n4022,
    new_n4023, new_n4024, new_n4025, new_n4026, new_n4027, new_n4028,
    new_n4029, new_n4031, new_n4032, new_n4033, new_n4034, new_n4035,
    new_n4036, new_n4037, new_n4038, new_n4039, new_n4040, new_n4041,
    new_n4042, new_n4043, new_n4044, new_n4045, new_n4046, new_n4047,
    new_n4048, new_n4049, new_n4050, new_n4051, new_n4052, new_n4053,
    new_n4054, new_n4056, new_n4057, new_n4059, new_n4060, new_n4061,
    new_n4062, new_n4064, new_n4065, new_n4066, new_n4067, new_n4069,
    new_n4070, new_n4071, new_n4072, new_n4074, new_n4075, new_n4076,
    new_n4077, new_n4078, new_n4079, new_n4080, new_n4081, new_n4083,
    new_n4084, new_n4085, new_n4086, new_n4087, new_n4088, new_n4089,
    new_n4090, new_n4091, new_n4092, new_n4093, new_n4094, new_n4095,
    new_n4096, new_n4097, new_n4098, new_n4099, new_n4100, new_n4101,
    new_n4102, new_n4103, new_n4104, new_n4105, new_n4106, new_n4107,
    new_n4108, new_n4109, new_n4110, new_n4111, new_n4112, new_n4113,
    new_n4114, new_n4115, new_n4116, new_n4117, new_n4118, new_n4119,
    new_n4120, new_n4121, new_n4122, new_n4123, new_n4124, new_n4125,
    new_n4126, new_n4127, new_n4128, new_n4129, new_n4130, new_n4131,
    new_n4132, new_n4133, new_n4134, new_n4135, new_n4136, new_n4137,
    new_n4138, new_n4139, new_n4140, new_n4141, new_n4143, new_n4144,
    new_n4145, new_n4146, new_n4147, new_n4148, new_n4150, new_n4151,
    new_n4152, new_n4153, new_n4154, new_n4155, new_n4156, new_n4157,
    new_n4158, new_n4159, new_n4160, new_n4161, new_n4162, new_n4163,
    new_n4164, new_n4165, new_n4166, new_n4167, new_n4168, new_n4169,
    new_n4170, new_n4171, new_n4172, new_n4173, new_n4174, new_n4176,
    new_n4177, new_n4178, new_n4179, new_n4180, new_n4181, new_n4182,
    new_n4183, new_n4184, new_n4185, new_n4186, new_n4187, new_n4188,
    new_n4189, new_n4190, new_n4191, new_n4192, new_n4193, new_n4194,
    new_n4195, new_n4196, new_n4197, new_n4198, new_n4199, new_n4201,
    new_n4202, new_n4203, new_n4204, new_n4205, new_n4206, new_n4207,
    new_n4208, new_n4209, new_n4210, new_n4211, new_n4212, new_n4213,
    new_n4214, new_n4215, new_n4216, new_n4217, new_n4218, new_n4219,
    new_n4220, new_n4221, new_n4222, new_n4223, new_n4224, new_n4226,
    new_n4227, new_n4228, new_n4229, new_n4230, new_n4231, new_n4232,
    new_n4233, new_n4234, new_n4235, new_n4236, new_n4237, new_n4238,
    new_n4239, new_n4240, new_n4241, new_n4242, new_n4243, new_n4244,
    new_n4245, new_n4246, new_n4247, new_n4248, new_n4249, new_n4251,
    new_n4252, new_n4254, new_n4255, new_n4256, new_n4257, new_n4258,
    new_n4259, new_n4260, new_n4261, new_n4262, new_n4263, new_n4264,
    new_n4265, new_n4266, new_n4267, new_n4268, new_n4269, new_n4270,
    new_n4271, new_n4272, new_n4273, new_n4274, new_n4275, new_n4276,
    new_n4277, new_n4278, new_n4279, new_n4280, new_n4281, new_n4282,
    new_n4283, new_n4284, new_n4285, new_n4286, new_n4287, new_n4288,
    new_n4289, new_n4290, new_n4291, new_n4292, new_n4294, new_n4295,
    new_n4296, new_n4297, new_n4299, new_n4300, new_n4301, new_n4302,
    new_n4304, new_n4305, new_n4306, new_n4307, new_n4309, new_n4310,
    new_n4311, new_n4312, new_n4313, new_n4314, new_n4316, new_n4317,
    new_n4318, new_n4319, new_n4320, new_n4321, new_n4322, new_n4323,
    new_n4325, new_n4326, new_n4327, new_n4328, new_n4329, new_n4330,
    new_n4332, new_n4333, new_n4334, new_n4335, new_n4336, new_n4337,
    new_n4338, new_n4339, new_n4341, new_n4342, new_n4343, new_n4345,
    new_n4346, new_n4347, new_n4348, new_n4350, new_n4351, new_n4352,
    new_n4353, new_n4355, new_n4356, new_n4357, new_n4358, new_n4359,
    new_n4360, new_n4362, new_n4363, new_n4364, new_n4365, new_n4366,
    new_n4367, new_n4368, new_n4369, new_n4370, new_n4371, new_n4372,
    new_n4373, new_n4374, new_n4375, new_n4376, new_n4377, new_n4378,
    new_n4379, new_n4380, new_n4381, new_n4382, new_n4383, new_n4384,
    new_n4385, new_n4386, new_n4387, new_n4388, new_n4389, new_n4390,
    new_n4391, new_n4392, new_n4393, new_n4394, new_n4395, new_n4396,
    new_n4397, new_n4398, new_n4399, new_n4400, new_n4401, new_n4402,
    new_n4403, new_n4404, new_n4405, new_n4406, new_n4407, new_n4408,
    new_n4409, new_n4410, new_n4412, new_n4413, new_n4414, new_n4416,
    new_n4417, new_n4418, new_n4419, new_n4420, new_n4421, new_n4423,
    new_n4424, new_n4425, new_n4426, new_n4427, new_n4428, new_n4429,
    new_n4430, new_n4432, new_n4433, new_n4434, new_n4435, new_n4436,
    new_n4437, new_n4438, new_n4439, new_n4440, new_n4441, new_n4442,
    new_n4443, new_n4444, new_n4445, new_n4446, new_n4447, new_n4448,
    new_n4449, new_n4450, new_n4451, new_n4452, new_n4453, new_n4454,
    new_n4455, new_n4456, new_n4457, new_n4458, new_n4459, new_n4460,
    new_n4461, new_n4462, new_n4463, new_n4464, new_n4465, new_n4466,
    new_n4467, new_n4469, new_n4470, new_n4471, new_n4472, new_n4473,
    new_n4474, new_n4475, new_n4476, new_n4477, new_n4478, new_n4479,
    new_n4481, new_n4482, new_n4483, new_n4484, new_n4485, new_n4486,
    new_n4487, new_n4488, new_n4489, new_n4490, new_n4491, new_n4492,
    new_n4493, new_n4494, new_n4495, new_n4496, new_n4497, new_n4498,
    new_n4499, new_n4500, new_n4501, new_n4502, new_n4503, new_n4504,
    new_n4505, new_n4506, new_n4507, new_n4508, new_n4509, new_n4510,
    new_n4511, new_n4512, new_n4513, new_n4514, new_n4515, new_n4516,
    new_n4517, new_n4518, new_n4519, new_n4520, new_n4521, new_n4522,
    new_n4523, new_n4525, new_n4526, new_n4527, new_n4529, new_n4530,
    new_n4531, new_n4532, new_n4533, new_n4534, new_n4535, new_n4536,
    new_n4537, new_n4538, new_n4539, new_n4540, new_n4541, new_n4542,
    new_n4543, new_n4544, new_n4545, new_n4546, new_n4547, new_n4548,
    new_n4549, new_n4550, new_n4551, new_n4552, new_n4553, new_n4554,
    new_n4555, new_n4556, new_n4557, new_n4558, new_n4559, new_n4560,
    new_n4561, new_n4562, new_n4563, new_n4564, new_n4565, new_n4566,
    new_n4567, new_n4568, new_n4569, new_n4570, new_n4571, new_n4572,
    new_n4573, new_n4574, new_n4576, new_n4577, new_n4578, new_n4579,
    new_n4581, new_n4582, new_n4583, new_n4584, new_n4585, new_n4586,
    new_n4588, new_n4589, new_n4590, new_n4591, new_n4592, new_n4593,
    new_n4595, new_n4596, new_n4597, new_n4598, new_n4599, new_n4600,
    new_n4601, new_n4602, new_n4603, new_n4604, new_n4605, new_n4606,
    new_n4607, new_n4608, new_n4609, new_n4610, new_n4611, new_n4612,
    new_n4613, new_n4614, new_n4615, new_n4616, new_n4617, new_n4618,
    new_n4619, new_n4620, new_n4621, new_n4622, new_n4623, new_n4624,
    new_n4625, new_n4626, new_n4627, new_n4628, new_n4629, new_n4630,
    new_n4631, new_n4632, new_n4633, new_n4635, new_n4636, new_n4637,
    new_n4638, new_n4640, new_n4641, new_n4642, new_n4643, new_n4644,
    new_n4645, new_n4646, new_n4647, new_n4648, new_n4649, new_n4650,
    new_n4651, new_n4652, new_n4653, new_n4654, new_n4655, new_n4656,
    new_n4657, new_n4658, new_n4659, new_n4660, new_n4661, new_n4662,
    new_n4663, new_n4664, new_n4665, new_n4666, new_n4667, new_n4668,
    new_n4669, new_n4670, new_n4671, new_n4672, new_n4673, new_n4674,
    new_n4675, new_n4676, new_n4677, new_n4678, new_n4680, new_n4681,
    new_n4682, new_n4683, new_n4685, new_n4686, new_n4687, new_n4688,
    new_n4690, new_n4691, new_n4692, new_n4693, new_n4694, new_n4695,
    new_n4696, new_n4697, new_n4698, new_n4699, new_n4700, new_n4701,
    new_n4702, new_n4703, new_n4704, new_n4705, new_n4706, new_n4707,
    new_n4708, new_n4709, new_n4710, new_n4711, new_n4712, new_n4713,
    new_n4714, new_n4715, new_n4716, new_n4717, new_n4718, new_n4719,
    new_n4720, new_n4721, new_n4722, new_n4723, new_n4724, new_n4725,
    new_n4726, new_n4727, new_n4728, new_n4729, new_n4731, new_n4732,
    new_n4733, new_n4734, new_n4735, new_n4736, new_n4738, new_n4739,
    new_n4740, new_n4741, new_n4742, new_n4743, new_n4744, new_n4745,
    new_n4746, new_n4747, new_n4748, new_n4749, new_n4750, new_n4751,
    new_n4752, new_n4753, new_n4754, new_n4755, new_n4756, new_n4757,
    new_n4758, new_n4759, new_n4760, new_n4761, new_n4763, new_n4764,
    new_n4766, new_n4767, new_n4768, new_n4769, new_n4771, new_n4772,
    new_n4773, new_n4774, new_n4776, new_n4777, new_n4778, new_n4779,
    new_n4780, new_n4781, new_n4782, new_n4783, new_n4784, new_n4785,
    new_n4786, new_n4787, new_n4788, new_n4789, new_n4790, new_n4791,
    new_n4792, new_n4793, new_n4794, new_n4795, new_n4796, new_n4797,
    new_n4798, new_n4799, new_n4800, new_n4801, new_n4802, new_n4803,
    new_n4804, new_n4805, new_n4806, new_n4807, new_n4808, new_n4809,
    new_n4810, new_n4811, new_n4812, new_n4814, new_n4815, new_n4816,
    new_n4817, new_n4819, new_n4820, new_n4821, new_n4822, new_n4824,
    new_n4825, new_n4826, new_n4827, new_n4828, new_n4829, new_n4831,
    new_n4832, new_n4833, new_n4834, new_n4835, new_n4836, new_n4837,
    new_n4838, new_n4840, new_n4841, new_n4842, new_n4843, new_n4844,
    new_n4845, new_n4847, new_n4848, new_n4849, new_n4850, new_n4851,
    new_n4853, new_n4854, new_n4855, new_n4856, new_n4857, new_n4858,
    new_n4859, new_n4860, new_n4861, new_n4862, new_n4863, new_n4864,
    new_n4865, new_n4866, new_n4867, new_n4868, new_n4869, new_n4870,
    new_n4871, new_n4872, new_n4873, new_n4874, new_n4875, new_n4876,
    new_n4878, new_n4879, new_n4880, new_n4881, new_n4882, new_n4883,
    new_n4884, new_n4885, new_n4886, new_n4887, new_n4888, new_n4889,
    new_n4890, new_n4891, new_n4892, new_n4893, new_n4894, new_n4895,
    new_n4896, new_n4897, new_n4898, new_n4899, new_n4900, new_n4901,
    new_n4902, new_n4904, new_n4905, new_n4906, new_n4907, new_n4909,
    new_n4910, new_n4911, new_n4912, new_n4914, new_n4915, new_n4916,
    new_n4917, new_n4919, new_n4920, new_n4921, new_n4922, new_n4924,
    new_n4925, new_n4926, new_n4927, new_n4928, new_n4929, new_n4930,
    new_n4931, new_n4933, new_n4934, new_n4935, new_n4936, new_n4937,
    new_n4938, new_n4940, new_n4941, new_n4942, new_n4943, new_n4944,
    new_n4945, new_n4946, new_n4947, new_n4948, new_n4949, new_n4950,
    new_n4951, new_n4952, new_n4953, new_n4954, new_n4955, new_n4956,
    new_n4957, new_n4958, new_n4959, new_n4960, new_n4961, new_n4962,
    new_n4963, new_n4964, new_n4966, new_n4967, new_n4968, new_n4969,
    new_n4971, new_n4972, new_n4973, new_n4974, new_n4976, new_n4977,
    new_n4978, new_n4979, new_n4981, new_n4982, new_n4983, new_n4984,
    new_n4986, new_n4987, new_n4988, new_n4989, new_n4990, new_n4991,
    new_n4993, new_n4994, new_n4995, new_n4996, new_n4997, new_n4998,
    new_n4999, new_n5000, new_n5002, new_n5003, new_n5004, new_n5005,
    new_n5007, new_n5008, new_n5009, new_n5010, new_n5012, new_n5013,
    new_n5014, new_n5015, new_n5016, new_n5017, new_n5019, new_n5020,
    new_n5022, new_n5023, new_n5025, new_n5026, new_n5027, new_n5028,
    new_n5030, new_n5031, new_n5032, new_n5033, new_n5034, new_n5035,
    new_n5036, new_n5037, new_n5039, new_n5040, new_n5041, new_n5042,
    new_n5044, new_n5045, new_n5046, new_n5047, new_n5048, new_n5049,
    new_n5051, new_n5052, new_n5054, new_n5055, new_n5056, new_n5057,
    new_n5059, new_n5060, new_n5061, new_n5062, new_n5063, new_n5064,
    new_n5065, new_n5066, new_n5068, new_n5069, new_n5070, new_n5071,
    new_n5072, new_n5073, new_n5074, new_n5075, new_n5076, new_n5077,
    new_n5078, new_n5079, new_n5080, new_n5081, new_n5082, new_n5083,
    new_n5084, new_n5085, new_n5086, new_n5087, new_n5088, new_n5089,
    new_n5090, new_n5091, new_n5092, new_n5094, new_n5095, new_n5097,
    new_n5098, new_n5100, new_n5101, new_n5103, new_n5104, new_n5106,
    new_n5107, new_n5108, new_n5109, new_n5111, new_n5112, new_n5113,
    new_n5114, new_n5115, new_n5116, new_n5117, new_n5118, new_n5119,
    new_n5120, new_n5121, new_n5122, new_n5123, new_n5124, new_n5125,
    new_n5126, new_n5127, new_n5128, new_n5129, new_n5130, new_n5131,
    new_n5132, new_n5133, new_n5134, new_n5136, new_n5137, new_n5138,
    new_n5139, new_n5140, new_n5141, new_n5142, new_n5143, new_n5144,
    new_n5145, new_n5146, new_n5147, new_n5148, new_n5149, new_n5150,
    new_n5151, new_n5152, new_n5153, new_n5154, new_n5155, new_n5156,
    new_n5157, new_n5158, new_n5159, new_n5161, new_n5162, new_n5164,
    new_n5165, new_n5167, new_n5168, new_n5170, new_n5171, new_n5172,
    new_n5173, new_n5174, new_n5175, new_n5177, new_n5178, new_n5179,
    new_n5180, new_n5181, new_n5182, new_n5183, new_n5184, new_n5185,
    new_n5186, new_n5187, new_n5188, new_n5189, new_n5190, new_n5191,
    new_n5192, new_n5193, new_n5194, new_n5195, new_n5196, new_n5197,
    new_n5198, new_n5199, new_n5200, new_n5202, new_n5203, new_n5204,
    new_n5205, new_n5206, new_n5207, new_n5208, new_n5209, new_n5210,
    new_n5211, new_n5212, new_n5213, new_n5214, new_n5215, new_n5216,
    new_n5217, new_n5218, new_n5219, new_n5220, new_n5221, new_n5222,
    new_n5223, new_n5224, new_n5225, new_n5227, new_n5228, new_n5230,
    new_n5231;
  assign new_n502 = pcount_3_ & pencrypt_0_;
  assign new_n503 = pcount_1_ & new_n502;
  assign new_n504 = pcount_2_ & new_n503;
  assign new_n505 = pcount_0_ & new_n504;
  assign new_n506 = ~pencrypt_mode_0_ & new_n505;
  assign new_n507 = pcount_3_ & ~pencrypt_0_;
  assign new_n508 = pcount_1_ & new_n507;
  assign new_n509 = pcount_2_ & new_n508;
  assign new_n510 = pcount_0_ & new_n509;
  assign new_n511 = pencrypt_mode_0_ & new_n510;
  assign new_n512 = ~new_n506 & ~new_n511;
  assign new_n513 = ~pcount_3_ & ~pcount_1_;
  assign new_n514 = ~pcount_2_ & new_n513;
  assign new_n515 = ~pcount_0_ & new_n514;
  assign new_n516 = pcount_3_ & pcount_1_;
  assign new_n517 = pcount_2_ & new_n516;
  assign new_n518 = ~pcount_0_ & new_n517;
  assign new_n519 = ~pcount_3_ & pcount_1_;
  assign new_n520 = pcount_2_ & new_n519;
  assign new_n521 = pcount_0_ & new_n520;
  assign new_n522 = pcount_0_ & new_n517;
  assign new_n523 = ~new_n515 & ~new_n518;
  assign new_n524 = ~new_n521 & ~new_n522;
  assign new_n525 = new_n523 & new_n524;
  assign new_n526 = pcount_3_ & pload_key_0_;
  assign new_n527 = pcount_1_ & new_n526;
  assign new_n528 = pcount_2_ & new_n527;
  assign new_n529 = pcount_0_ & new_n528;
  assign new_n530 = new_n512 & ~new_n525;
  assign new_n531 = pc_5_ & new_n530;
  assign new_n532 = ~pencrypt_mode_0_ & new_n531;
  assign new_n533 = ~new_n529 & new_n532;
  assign new_n534 = ~preset_0_ & new_n533;
  assign new_n535 = new_n512 & new_n525;
  assign new_n536 = pc_8_ & new_n535;
  assign new_n537 = pencrypt_mode_0_ & new_n536;
  assign new_n538 = ~new_n529 & new_n537;
  assign new_n539 = ~preset_0_ & new_n538;
  assign new_n540 = ~preset_0_ & pc_6_;
  assign new_n541 = ~new_n512 & new_n540;
  assign new_n542 = ~new_n529 & new_n541;
  assign new_n543 = pc_7_ & new_n530;
  assign new_n544 = pencrypt_mode_0_ & new_n543;
  assign new_n545 = ~new_n529 & new_n544;
  assign new_n546 = ~preset_0_ & new_n545;
  assign new_n547 = ~preset_0_ & pdata_in_0_;
  assign new_n548 = pencrypt_0_ & new_n547;
  assign new_n549 = new_n529 & new_n548;
  assign new_n550 = pc_4_ & new_n535;
  assign new_n551 = ~pencrypt_mode_0_ & new_n550;
  assign new_n552 = ~new_n529 & new_n551;
  assign new_n553 = ~preset_0_ & new_n552;
  assign new_n554 = ~preset_0_ & ~pencrypt_0_;
  assign new_n555 = pinreg_0_ & new_n554;
  assign new_n556 = new_n529 & new_n555;
  assign new_n557 = ~new_n549 & ~new_n553;
  assign new_n558 = ~new_n556 & new_n557;
  assign new_n559 = ~new_n534 & ~new_n539;
  assign new_n560 = ~new_n542 & ~new_n546;
  assign new_n561 = new_n559 & new_n560;
  assign pc_new_6_ = ~new_n558 | ~new_n561;
  assign new_n563 = pc_21_ & new_n535;
  assign new_n564 = pencrypt_mode_0_ & new_n563;
  assign new_n565 = ~new_n529 & new_n564;
  assign new_n566 = ~preset_0_ & new_n565;
  assign new_n567 = pc_17_ & new_n535;
  assign new_n568 = ~pencrypt_mode_0_ & new_n567;
  assign new_n569 = ~new_n529 & new_n568;
  assign new_n570 = ~preset_0_ & new_n569;
  assign new_n571 = pc_20_ & new_n530;
  assign new_n572 = pencrypt_mode_0_ & new_n571;
  assign new_n573 = ~new_n529 & new_n572;
  assign new_n574 = ~preset_0_ & new_n573;
  assign new_n575 = pc_18_ & new_n530;
  assign new_n576 = ~pencrypt_mode_0_ & new_n575;
  assign new_n577 = ~new_n529 & new_n576;
  assign new_n578 = ~preset_0_ & new_n577;
  assign new_n579 = ~preset_0_ & pc_19_;
  assign new_n580 = ~new_n512 & new_n579;
  assign new_n581 = ~new_n529 & new_n580;
  assign new_n582 = ~preset_0_ & pencrypt_0_;
  assign new_n583 = pinreg_18_ & new_n582;
  assign new_n584 = new_n529 & new_n583;
  assign new_n585 = pinreg_26_ & new_n554;
  assign new_n586 = new_n529 & new_n585;
  assign new_n587 = ~new_n581 & ~new_n584;
  assign new_n588 = ~new_n586 & new_n587;
  assign new_n589 = ~new_n566 & ~new_n570;
  assign new_n590 = ~new_n574 & ~new_n578;
  assign new_n591 = new_n589 & new_n590;
  assign pc_new_19_ = ~new_n588 | ~new_n591;
  assign new_n593 = pd_7_ & new_n535;
  assign new_n594 = pencrypt_mode_0_ & new_n593;
  assign new_n595 = ~new_n529 & new_n594;
  assign new_n596 = ~preset_0_ & new_n595;
  assign new_n597 = pd_3_ & new_n535;
  assign new_n598 = ~pencrypt_mode_0_ & new_n597;
  assign new_n599 = ~new_n529 & new_n598;
  assign new_n600 = ~preset_0_ & new_n599;
  assign new_n601 = pd_6_ & new_n530;
  assign new_n602 = pencrypt_mode_0_ & new_n601;
  assign new_n603 = ~new_n529 & new_n602;
  assign new_n604 = ~preset_0_ & new_n603;
  assign new_n605 = pd_4_ & new_n530;
  assign new_n606 = ~pencrypt_mode_0_ & new_n605;
  assign new_n607 = ~new_n529 & new_n606;
  assign new_n608 = ~preset_0_ & new_n607;
  assign new_n609 = ~preset_0_ & pd_5_;
  assign new_n610 = ~new_n512 & new_n609;
  assign new_n611 = ~new_n529 & new_n610;
  assign new_n612 = pinreg_14_ & new_n554;
  assign new_n613 = new_n529 & new_n612;
  assign new_n614 = pinreg_6_ & new_n582;
  assign new_n615 = new_n529 & new_n614;
  assign new_n616 = ~new_n611 & ~new_n613;
  assign new_n617 = ~new_n615 & new_n616;
  assign new_n618 = ~new_n596 & ~new_n600;
  assign new_n619 = ~new_n604 & ~new_n608;
  assign new_n620 = new_n618 & new_n619;
  assign pd_new_5_ = ~new_n617 | ~new_n620;
  assign new_n622 = pinreg_3_ & new_n522;
  assign new_n623 = pdata_46_ & ~new_n522;
  assign pdata_new_14_ = new_n622 | new_n623;
  assign new_n625 = pinreg_31_ & new_n522;
  assign new_n626 = pdata_59_ & ~new_n522;
  assign pdata_new_27_ = new_n625 | new_n626;
  assign new_n628 = ~pcount_0_ & pinreg_6_;
  assign new_n629 = ~new_n522 & new_n628;
  assign new_n630 = pcount_0_ & pdata_in_6_;
  assign new_n631 = ~new_n522 & new_n630;
  assign pinreg_new_6_ = new_n629 | new_n631;
  assign new_n633 = ~pcount_0_ & pinreg_19_;
  assign new_n634 = ~new_n522 & new_n633;
  assign new_n635 = pcount_0_ & pinreg_11_;
  assign new_n636 = ~new_n522 & new_n635;
  assign pinreg_new_19_ = new_n634 | new_n636;
  assign new_n638 = pd_27_ & ~pdata_58_;
  assign new_n639 = ~pd_27_ & pdata_58_;
  assign new_n640 = ~new_n638 & ~new_n639;
  assign new_n641 = ~pdata_59_ & pd_5_;
  assign new_n642 = pdata_59_ & ~pd_5_;
  assign new_n643 = ~new_n641 & ~new_n642;
  assign new_n644 = pd_20_ & ~pdata_56_;
  assign new_n645 = ~pd_20_ & pdata_56_;
  assign new_n646 = ~new_n644 & ~new_n645;
  assign new_n647 = pd_10_ & ~pdata_57_;
  assign new_n648 = ~pd_10_ & pdata_57_;
  assign new_n649 = ~new_n647 & ~new_n648;
  assign new_n650 = pd_15_ & ~pdata_55_;
  assign new_n651 = ~pd_15_ & pdata_55_;
  assign new_n652 = ~new_n650 & ~new_n651;
  assign new_n653 = ~pdata_60_ & pd_24_;
  assign new_n654 = pdata_60_ & ~pd_24_;
  assign new_n655 = ~new_n653 & ~new_n654;
  assign new_n656 = new_n640 & new_n643;
  assign new_n657 = ~new_n646 & new_n656;
  assign new_n658 = new_n649 & new_n657;
  assign new_n659 = new_n652 & new_n658;
  assign new_n660 = new_n655 & new_n659;
  assign new_n661 = ~new_n640 & new_n643;
  assign new_n662 = ~new_n646 & new_n661;
  assign new_n663 = new_n649 & new_n662;
  assign new_n664 = new_n652 & new_n663;
  assign new_n665 = new_n655 & new_n664;
  assign new_n666 = new_n646 & new_n656;
  assign new_n667 = ~new_n649 & new_n666;
  assign new_n668 = new_n652 & new_n667;
  assign new_n669 = new_n655 & new_n668;
  assign new_n670 = ~new_n640 & ~new_n643;
  assign new_n671 = new_n646 & new_n670;
  assign new_n672 = ~new_n649 & new_n671;
  assign new_n673 = new_n652 & new_n672;
  assign new_n674 = new_n655 & new_n673;
  assign new_n675 = new_n640 & ~new_n643;
  assign new_n676 = new_n646 & new_n675;
  assign new_n677 = new_n649 & new_n676;
  assign new_n678 = new_n652 & new_n677;
  assign new_n679 = new_n655 & new_n678;
  assign new_n680 = ~new_n649 & new_n662;
  assign new_n681 = ~new_n652 & new_n680;
  assign new_n682 = ~new_n655 & new_n681;
  assign new_n683 = ~new_n649 & new_n676;
  assign new_n684 = ~new_n652 & new_n683;
  assign new_n685 = new_n655 & new_n684;
  assign new_n686 = ~new_n646 & new_n670;
  assign new_n687 = new_n649 & new_n686;
  assign new_n688 = ~new_n652 & new_n687;
  assign new_n689 = ~new_n655 & new_n688;
  assign new_n690 = new_n646 & new_n661;
  assign new_n691 = ~new_n649 & new_n690;
  assign new_n692 = ~new_n652 & new_n691;
  assign new_n693 = new_n655 & new_n692;
  assign new_n694 = ~new_n652 & new_n667;
  assign new_n695 = ~new_n655 & new_n694;
  assign new_n696 = ~new_n646 & new_n675;
  assign new_n697 = new_n649 & new_n696;
  assign new_n698 = ~new_n652 & new_n697;
  assign new_n699 = new_n655 & new_n698;
  assign new_n700 = new_n652 & new_n691;
  assign new_n701 = ~new_n655 & new_n700;
  assign new_n702 = ~new_n649 & new_n696;
  assign new_n703 = ~new_n652 & new_n702;
  assign new_n704 = new_n655 & new_n703;
  assign new_n705 = ~new_n652 & new_n672;
  assign new_n706 = ~new_n655 & new_n705;
  assign new_n707 = ~new_n655 & new_n664;
  assign new_n708 = new_n649 & new_n690;
  assign new_n709 = ~new_n652 & new_n708;
  assign new_n710 = ~new_n655 & new_n709;
  assign new_n711 = new_n652 & new_n702;
  assign new_n712 = ~new_n655 & new_n711;
  assign new_n713 = ~new_n655 & new_n698;
  assign new_n714 = new_n655 & new_n709;
  assign new_n715 = ~new_n652 & new_n658;
  assign new_n716 = ~new_n655 & new_n715;
  assign new_n717 = new_n649 & new_n671;
  assign new_n718 = ~new_n652 & new_n717;
  assign new_n719 = new_n655 & new_n718;
  assign new_n720 = ~new_n649 & new_n686;
  assign new_n721 = new_n652 & new_n720;
  assign new_n722 = new_n655 & new_n721;
  assign new_n723 = new_n649 & new_n666;
  assign new_n724 = ~new_n652 & new_n723;
  assign new_n725 = new_n655 & new_n724;
  assign new_n726 = ~new_n652 & new_n677;
  assign new_n727 = ~new_n655 & new_n726;
  assign new_n728 = new_n652 & new_n683;
  assign new_n729 = ~new_n655 & new_n728;
  assign new_n730 = new_n655 & new_n681;
  assign new_n731 = new_n652 & new_n697;
  assign new_n732 = ~new_n655 & new_n731;
  assign new_n733 = new_n652 & new_n717;
  assign new_n734 = ~new_n655 & new_n733;
  assign new_n735 = new_n652 & new_n723;
  assign new_n736 = ~new_n655 & new_n735;
  assign new_n737 = new_n652 & new_n708;
  assign new_n738 = ~new_n655 & new_n737;
  assign new_n739 = new_n652 & new_n687;
  assign new_n740 = new_n655 & new_n739;
  assign new_n741 = ~new_n649 & new_n657;
  assign new_n742 = new_n652 & new_n741;
  assign new_n743 = new_n655 & new_n742;
  assign new_n744 = ~new_n740 & ~new_n743;
  assign new_n745 = ~new_n736 & ~new_n738;
  assign new_n746 = new_n744 & new_n745;
  assign new_n747 = ~new_n732 & ~new_n734;
  assign new_n748 = ~new_n729 & ~new_n730;
  assign new_n749 = new_n747 & new_n748;
  assign new_n750 = new_n746 & new_n749;
  assign new_n751 = ~new_n725 & ~new_n727;
  assign new_n752 = ~new_n719 & ~new_n722;
  assign new_n753 = new_n751 & new_n752;
  assign new_n754 = ~new_n714 & ~new_n716;
  assign new_n755 = ~new_n712 & ~new_n713;
  assign new_n756 = new_n754 & new_n755;
  assign new_n757 = new_n753 & new_n756;
  assign new_n758 = new_n750 & new_n757;
  assign new_n759 = ~new_n707 & ~new_n710;
  assign new_n760 = ~new_n704 & ~new_n706;
  assign new_n761 = new_n759 & new_n760;
  assign new_n762 = ~new_n699 & ~new_n701;
  assign new_n763 = ~new_n693 & ~new_n695;
  assign new_n764 = new_n762 & new_n763;
  assign new_n765 = new_n761 & new_n764;
  assign new_n766 = ~new_n660 & ~new_n665;
  assign new_n767 = ~new_n669 & ~new_n674;
  assign new_n768 = new_n766 & new_n767;
  assign new_n769 = ~new_n679 & ~new_n682;
  assign new_n770 = ~new_n685 & ~new_n689;
  assign new_n771 = new_n769 & new_n770;
  assign new_n772 = new_n768 & new_n771;
  assign new_n773 = new_n765 & new_n772;
  assign new_n774 = new_n758 & new_n773;
  assign new_n775 = pdata_6_ & new_n774;
  assign new_n776 = new_n522 & new_n775;
  assign new_n777 = ~pcount_0_ & poutreg_9_;
  assign new_n778 = ~new_n522 & new_n777;
  assign new_n779 = ~pdata_6_ & ~new_n774;
  assign new_n780 = new_n522 & new_n779;
  assign new_n781 = pcount_0_ & poutreg_17_;
  assign new_n782 = ~new_n522 & new_n781;
  assign new_n783 = ~new_n776 & ~new_n778;
  assign new_n784 = ~new_n780 & ~new_n782;
  assign poutreg_new_9_ = ~new_n783 | ~new_n784;
  assign new_n786 = pc_6_ & new_n530;
  assign new_n787 = ~pencrypt_mode_0_ & new_n786;
  assign new_n788 = ~new_n529 & new_n787;
  assign new_n789 = ~preset_0_ & new_n788;
  assign new_n790 = pc_9_ & new_n535;
  assign new_n791 = pencrypt_mode_0_ & new_n790;
  assign new_n792 = ~new_n529 & new_n791;
  assign new_n793 = ~preset_0_ & new_n792;
  assign new_n794 = ~preset_0_ & pc_7_;
  assign new_n795 = ~new_n512 & new_n794;
  assign new_n796 = ~new_n529 & new_n795;
  assign new_n797 = pc_8_ & new_n530;
  assign new_n798 = pencrypt_mode_0_ & new_n797;
  assign new_n799 = ~new_n529 & new_n798;
  assign new_n800 = ~preset_0_ & new_n799;
  assign new_n801 = ~pencrypt_0_ & new_n547;
  assign new_n802 = new_n529 & new_n801;
  assign new_n803 = pc_5_ & new_n535;
  assign new_n804 = ~pencrypt_mode_0_ & new_n803;
  assign new_n805 = ~new_n529 & new_n804;
  assign new_n806 = ~preset_0_ & new_n805;
  assign new_n807 = pinreg_49_ & new_n582;
  assign new_n808 = new_n529 & new_n807;
  assign new_n809 = ~new_n802 & ~new_n806;
  assign new_n810 = ~new_n808 & new_n809;
  assign new_n811 = ~new_n789 & ~new_n793;
  assign new_n812 = ~new_n796 & ~new_n800;
  assign new_n813 = new_n811 & new_n812;
  assign pc_new_7_ = ~new_n810 | ~new_n813;
  assign new_n815 = pd_5_ & new_n530;
  assign new_n816 = ~pencrypt_mode_0_ & new_n815;
  assign new_n817 = ~new_n529 & new_n816;
  assign new_n818 = ~preset_0_ & new_n817;
  assign new_n819 = pd_8_ & new_n535;
  assign new_n820 = pencrypt_mode_0_ & new_n819;
  assign new_n821 = ~new_n529 & new_n820;
  assign new_n822 = ~preset_0_ & new_n821;
  assign new_n823 = ~preset_0_ & pd_6_;
  assign new_n824 = ~new_n512 & new_n823;
  assign new_n825 = ~new_n529 & new_n824;
  assign new_n826 = pd_7_ & new_n530;
  assign new_n827 = pencrypt_mode_0_ & new_n826;
  assign new_n828 = ~new_n529 & new_n827;
  assign new_n829 = ~preset_0_ & new_n828;
  assign new_n830 = ~preset_0_ & pdata_in_6_;
  assign new_n831 = pencrypt_0_ & new_n830;
  assign new_n832 = new_n529 & new_n831;
  assign new_n833 = pd_4_ & new_n535;
  assign new_n834 = ~pencrypt_mode_0_ & new_n833;
  assign new_n835 = ~new_n529 & new_n834;
  assign new_n836 = ~preset_0_ & new_n835;
  assign new_n837 = pinreg_6_ & new_n554;
  assign new_n838 = new_n529 & new_n837;
  assign new_n839 = ~new_n832 & ~new_n836;
  assign new_n840 = ~new_n838 & new_n839;
  assign new_n841 = ~new_n818 & ~new_n822;
  assign new_n842 = ~new_n825 & ~new_n829;
  assign new_n843 = new_n841 & new_n842;
  assign pd_new_6_ = ~new_n840 | ~new_n843;
  assign new_n845 = pd_21_ & new_n535;
  assign new_n846 = pencrypt_mode_0_ & new_n845;
  assign new_n847 = ~new_n529 & new_n846;
  assign new_n848 = ~preset_0_ & new_n847;
  assign new_n849 = pd_17_ & new_n535;
  assign new_n850 = ~pencrypt_mode_0_ & new_n849;
  assign new_n851 = ~new_n529 & new_n850;
  assign new_n852 = ~preset_0_ & new_n851;
  assign new_n853 = pd_20_ & new_n530;
  assign new_n854 = pencrypt_mode_0_ & new_n853;
  assign new_n855 = ~new_n529 & new_n854;
  assign new_n856 = ~preset_0_ & new_n855;
  assign new_n857 = pd_18_ & new_n530;
  assign new_n858 = ~pencrypt_mode_0_ & new_n857;
  assign new_n859 = ~new_n529 & new_n858;
  assign new_n860 = ~preset_0_ & new_n859;
  assign new_n861 = ~preset_0_ & pd_19_;
  assign new_n862 = ~new_n512 & new_n861;
  assign new_n863 = ~new_n529 & new_n862;
  assign new_n864 = pinreg_20_ & new_n582;
  assign new_n865 = new_n529 & new_n864;
  assign new_n866 = pinreg_28_ & new_n554;
  assign new_n867 = new_n529 & new_n866;
  assign new_n868 = ~new_n863 & ~new_n865;
  assign new_n869 = ~new_n867 & new_n868;
  assign new_n870 = ~new_n848 & ~new_n852;
  assign new_n871 = ~new_n856 & ~new_n860;
  assign new_n872 = new_n870 & new_n871;
  assign pd_new_19_ = ~new_n869 | ~new_n872;
  assign new_n874 = pinreg_11_ & new_n522;
  assign new_n875 = pdata_45_ & ~new_n522;
  assign pdata_new_13_ = new_n874 | new_n875;
  assign new_n877 = pinreg_23_ & new_n522;
  assign new_n878 = pdata_60_ & ~new_n522;
  assign pdata_new_28_ = new_n877 | new_n878;
  assign new_n880 = pd_8_ & ~pdata_50_;
  assign new_n881 = ~pd_8_ & pdata_50_;
  assign new_n882 = ~new_n880 & ~new_n881;
  assign new_n883 = pd_18_ & ~pdata_51_;
  assign new_n884 = ~pd_18_ & pdata_51_;
  assign new_n885 = ~new_n883 & ~new_n884;
  assign new_n886 = ~pdata_48_ & pd_23_;
  assign new_n887 = pdata_48_ & ~pd_23_;
  assign new_n888 = ~new_n886 & ~new_n887;
  assign new_n889 = pd_2_ & ~pdata_49_;
  assign new_n890 = ~pd_2_ & pdata_49_;
  assign new_n891 = ~new_n889 & ~new_n890;
  assign new_n892 = ~pdata_47_ & pd_12_;
  assign new_n893 = pdata_47_ & ~pd_12_;
  assign new_n894 = ~new_n892 & ~new_n893;
  assign new_n895 = pd_26_ & ~pdata_52_;
  assign new_n896 = ~pd_26_ & pdata_52_;
  assign new_n897 = ~new_n895 & ~new_n896;
  assign new_n898 = ~new_n882 & ~new_n885;
  assign new_n899 = ~new_n888 & new_n898;
  assign new_n900 = new_n891 & new_n899;
  assign new_n901 = new_n894 & new_n900;
  assign new_n902 = new_n897 & new_n901;
  assign new_n903 = new_n882 & new_n885;
  assign new_n904 = ~new_n888 & new_n903;
  assign new_n905 = ~new_n891 & new_n904;
  assign new_n906 = new_n894 & new_n905;
  assign new_n907 = new_n897 & new_n906;
  assign new_n908 = new_n882 & ~new_n885;
  assign new_n909 = new_n888 & new_n908;
  assign new_n910 = ~new_n891 & new_n909;
  assign new_n911 = new_n894 & new_n910;
  assign new_n912 = new_n897 & new_n911;
  assign new_n913 = ~new_n882 & new_n885;
  assign new_n914 = new_n888 & new_n913;
  assign new_n915 = ~new_n891 & new_n914;
  assign new_n916 = new_n894 & new_n915;
  assign new_n917 = new_n897 & new_n916;
  assign new_n918 = new_n891 & new_n909;
  assign new_n919 = new_n894 & new_n918;
  assign new_n920 = new_n897 & new_n919;
  assign new_n921 = ~new_n894 & new_n905;
  assign new_n922 = ~new_n897 & new_n921;
  assign new_n923 = ~new_n894 & new_n910;
  assign new_n924 = new_n897 & new_n923;
  assign new_n925 = ~new_n894 & new_n900;
  assign new_n926 = ~new_n897 & new_n925;
  assign new_n927 = new_n891 & new_n904;
  assign new_n928 = ~new_n894 & new_n927;
  assign new_n929 = new_n897 & new_n928;
  assign new_n930 = ~new_n888 & new_n913;
  assign new_n931 = ~new_n891 & new_n930;
  assign new_n932 = new_n894 & new_n931;
  assign new_n933 = ~new_n897 & new_n932;
  assign new_n934 = ~new_n888 & new_n908;
  assign new_n935 = new_n891 & new_n934;
  assign new_n936 = ~new_n894 & new_n935;
  assign new_n937 = new_n897 & new_n936;
  assign new_n938 = ~new_n894 & new_n918;
  assign new_n939 = ~new_n897 & new_n938;
  assign new_n940 = new_n891 & new_n930;
  assign new_n941 = ~new_n894 & new_n940;
  assign new_n942 = new_n897 & new_n941;
  assign new_n943 = ~new_n897 & new_n923;
  assign new_n944 = ~new_n897 & new_n901;
  assign new_n945 = new_n891 & new_n914;
  assign new_n946 = ~new_n894 & new_n945;
  assign new_n947 = ~new_n897 & new_n946;
  assign new_n948 = ~new_n891 & new_n934;
  assign new_n949 = new_n894 & new_n948;
  assign new_n950 = ~new_n897 & new_n949;
  assign new_n951 = ~new_n897 & new_n936;
  assign new_n952 = new_n888 & new_n898;
  assign new_n953 = new_n891 & new_n952;
  assign new_n954 = ~new_n894 & new_n953;
  assign new_n955 = new_n897 & new_n954;
  assign new_n956 = ~new_n891 & new_n952;
  assign new_n957 = ~new_n894 & new_n956;
  assign new_n958 = ~new_n897 & new_n957;
  assign new_n959 = new_n888 & new_n903;
  assign new_n960 = ~new_n891 & new_n959;
  assign new_n961 = ~new_n894 & new_n960;
  assign new_n962 = new_n897 & new_n961;
  assign new_n963 = new_n897 & new_n957;
  assign new_n964 = new_n894 & new_n927;
  assign new_n965 = new_n897 & new_n964;
  assign new_n966 = new_n891 & new_n959;
  assign new_n967 = ~new_n894 & new_n966;
  assign new_n968 = ~new_n897 & new_n967;
  assign new_n969 = ~new_n897 & new_n916;
  assign new_n970 = ~new_n891 & new_n899;
  assign new_n971 = ~new_n894 & new_n970;
  assign new_n972 = new_n897 & new_n971;
  assign new_n973 = new_n894 & new_n940;
  assign new_n974 = ~new_n897 & new_n973;
  assign new_n975 = new_n894 & new_n953;
  assign new_n976 = ~new_n897 & new_n975;
  assign new_n977 = new_n894 & new_n966;
  assign new_n978 = ~new_n897 & new_n977;
  assign new_n979 = ~new_n897 & new_n919;
  assign new_n980 = new_n897 & new_n932;
  assign new_n981 = new_n894 & new_n970;
  assign new_n982 = new_n897 & new_n981;
  assign new_n983 = ~new_n980 & ~new_n982;
  assign new_n984 = ~new_n978 & ~new_n979;
  assign new_n985 = new_n983 & new_n984;
  assign new_n986 = ~new_n974 & ~new_n976;
  assign new_n987 = ~new_n969 & ~new_n972;
  assign new_n988 = new_n986 & new_n987;
  assign new_n989 = new_n985 & new_n988;
  assign new_n990 = ~new_n965 & ~new_n968;
  assign new_n991 = ~new_n962 & ~new_n963;
  assign new_n992 = new_n990 & new_n991;
  assign new_n993 = ~new_n955 & ~new_n958;
  assign new_n994 = ~new_n950 & ~new_n951;
  assign new_n995 = new_n993 & new_n994;
  assign new_n996 = new_n992 & new_n995;
  assign new_n997 = new_n989 & new_n996;
  assign new_n998 = ~new_n944 & ~new_n947;
  assign new_n999 = ~new_n942 & ~new_n943;
  assign new_n1000 = new_n998 & new_n999;
  assign new_n1001 = ~new_n937 & ~new_n939;
  assign new_n1002 = ~new_n929 & ~new_n933;
  assign new_n1003 = new_n1001 & new_n1002;
  assign new_n1004 = new_n1000 & new_n1003;
  assign new_n1005 = ~new_n902 & ~new_n907;
  assign new_n1006 = ~new_n912 & ~new_n917;
  assign new_n1007 = new_n1005 & new_n1006;
  assign new_n1008 = ~new_n920 & ~new_n922;
  assign new_n1009 = ~new_n924 & ~new_n926;
  assign new_n1010 = new_n1008 & new_n1009;
  assign new_n1011 = new_n1007 & new_n1010;
  assign new_n1012 = new_n1004 & new_n1011;
  assign new_n1013 = new_n997 & new_n1012;
  assign new_n1014 = ~pdata_7_ & ~new_n1013;
  assign new_n1015 = ~new_n522 & new_n1014;
  assign new_n1016 = pdata_7_ & new_n1013;
  assign new_n1017 = ~new_n522 & new_n1016;
  assign new_n1018 = pdata_in_0_ & new_n522;
  assign new_n1019 = ~new_n1015 & ~new_n1017;
  assign pdata_new_39_ = new_n1018 | ~new_n1019;
  assign new_n1021 = ~pcount_0_ & pinreg_5_;
  assign new_n1022 = ~new_n522 & new_n1021;
  assign new_n1023 = pcount_0_ & pdata_in_5_;
  assign new_n1024 = ~new_n522 & new_n1023;
  assign pinreg_new_5_ = new_n1022 | new_n1024;
  assign new_n1026 = ~pcount_0_ & pinreg_18_;
  assign new_n1027 = ~new_n522 & new_n1026;
  assign new_n1028 = pcount_0_ & pinreg_10_;
  assign new_n1029 = ~new_n522 & new_n1028;
  assign pinreg_new_18_ = new_n1027 | new_n1029;
  assign new_n1031 = new_n894 & new_n935;
  assign new_n1032 = new_n897 & new_n1031;
  assign new_n1033 = new_n894 & new_n960;
  assign new_n1034 = new_n897 & new_n1033;
  assign new_n1035 = new_n894 & new_n956;
  assign new_n1036 = new_n897 & new_n1035;
  assign new_n1037 = ~new_n894 & new_n931;
  assign new_n1038 = ~new_n897 & new_n1037;
  assign new_n1039 = ~new_n897 & new_n1033;
  assign new_n1040 = new_n897 & new_n925;
  assign new_n1041 = ~new_n894 & new_n948;
  assign new_n1042 = ~new_n897 & new_n1041;
  assign new_n1043 = new_n897 & new_n921;
  assign new_n1044 = ~new_n897 & new_n954;
  assign new_n1045 = ~new_n897 & new_n981;
  assign new_n1046 = ~new_n897 & new_n928;
  assign new_n1047 = ~new_n894 & new_n915;
  assign new_n1048 = new_n897 & new_n1047;
  assign new_n1049 = new_n894 & new_n945;
  assign new_n1050 = new_n897 & new_n1049;
  assign new_n1051 = new_n897 & new_n967;
  assign new_n1052 = ~new_n897 & new_n964;
  assign new_n1053 = ~new_n897 & new_n911;
  assign new_n1054 = ~new_n907 & ~new_n980;
  assign new_n1055 = ~new_n976 & ~new_n978;
  assign new_n1056 = new_n1054 & new_n1055;
  assign new_n1057 = ~new_n1052 & ~new_n1053;
  assign new_n1058 = new_n987 & new_n1057;
  assign new_n1059 = new_n1056 & new_n1058;
  assign new_n1060 = ~new_n947 & ~new_n1051;
  assign new_n1061 = ~new_n1048 & ~new_n1050;
  assign new_n1062 = new_n1060 & new_n1061;
  assign new_n1063 = ~new_n924 & ~new_n958;
  assign new_n1064 = ~new_n1045 & ~new_n1046;
  assign new_n1065 = new_n1063 & new_n1064;
  assign new_n1066 = new_n1062 & new_n1065;
  assign new_n1067 = new_n1059 & new_n1066;
  assign new_n1068 = ~new_n974 & ~new_n1044;
  assign new_n1069 = ~new_n943 & ~new_n1043;
  assign new_n1070 = new_n1068 & new_n1069;
  assign new_n1071 = ~new_n1040 & ~new_n1042;
  assign new_n1072 = ~new_n942 & ~new_n1039;
  assign new_n1073 = new_n1071 & new_n1072;
  assign new_n1074 = new_n1070 & new_n1073;
  assign new_n1075 = ~new_n902 & ~new_n1032;
  assign new_n1076 = ~new_n1034 & ~new_n1036;
  assign new_n1077 = new_n1075 & new_n1076;
  assign new_n1078 = ~new_n920 & ~new_n1038;
  assign new_n1079 = ~new_n929 & ~new_n951;
  assign new_n1080 = new_n1078 & new_n1079;
  assign new_n1081 = new_n1077 & new_n1080;
  assign new_n1082 = new_n1074 & new_n1081;
  assign new_n1083 = new_n1067 & new_n1082;
  assign new_n1084 = pdata_13_ & new_n1083;
  assign new_n1085 = new_n522 & new_n1084;
  assign new_n1086 = pcount_0_ & poutreg_27_;
  assign new_n1087 = ~new_n522 & new_n1086;
  assign new_n1088 = ~pdata_13_ & ~new_n1083;
  assign new_n1089 = new_n522 & new_n1088;
  assign new_n1090 = ~pcount_0_ & poutreg_19_;
  assign new_n1091 = ~new_n522 & new_n1090;
  assign new_n1092 = ~new_n1085 & ~new_n1087;
  assign new_n1093 = ~new_n1089 & ~new_n1091;
  assign poutreg_new_19_ = ~new_n1092 | ~new_n1093;
  assign new_n1095 = pc_6_ & new_n535;
  assign new_n1096 = pencrypt_mode_0_ & new_n1095;
  assign new_n1097 = ~new_n529 & new_n1096;
  assign new_n1098 = ~preset_0_ & new_n1097;
  assign new_n1099 = pc_2_ & new_n535;
  assign new_n1100 = ~pencrypt_mode_0_ & new_n1099;
  assign new_n1101 = ~new_n529 & new_n1100;
  assign new_n1102 = ~preset_0_ & new_n1101;
  assign new_n1103 = pencrypt_mode_0_ & new_n531;
  assign new_n1104 = ~new_n529 & new_n1103;
  assign new_n1105 = ~preset_0_ & new_n1104;
  assign new_n1106 = pc_3_ & new_n530;
  assign new_n1107 = ~pencrypt_mode_0_ & new_n1106;
  assign new_n1108 = ~new_n529 & new_n1107;
  assign new_n1109 = ~preset_0_ & new_n1108;
  assign new_n1110 = ~preset_0_ & pc_4_;
  assign new_n1111 = ~new_n512 & new_n1110;
  assign new_n1112 = ~new_n529 & new_n1111;
  assign new_n1113 = pinreg_16_ & new_n554;
  assign new_n1114 = new_n529 & new_n1113;
  assign new_n1115 = pinreg_8_ & new_n582;
  assign new_n1116 = new_n529 & new_n1115;
  assign new_n1117 = ~new_n1112 & ~new_n1114;
  assign new_n1118 = ~new_n1116 & new_n1117;
  assign new_n1119 = ~new_n1098 & ~new_n1102;
  assign new_n1120 = ~new_n1105 & ~new_n1109;
  assign new_n1121 = new_n1119 & new_n1120;
  assign pc_new_4_ = ~new_n1118 | ~new_n1121;
  assign new_n1123 = pd_5_ & new_n535;
  assign new_n1124 = pencrypt_mode_0_ & new_n1123;
  assign new_n1125 = ~new_n529 & new_n1124;
  assign new_n1126 = ~preset_0_ & new_n1125;
  assign new_n1127 = pd_1_ & new_n535;
  assign new_n1128 = ~pencrypt_mode_0_ & new_n1127;
  assign new_n1129 = ~new_n529 & new_n1128;
  assign new_n1130 = ~preset_0_ & new_n1129;
  assign new_n1131 = pencrypt_mode_0_ & new_n605;
  assign new_n1132 = ~new_n529 & new_n1131;
  assign new_n1133 = ~preset_0_ & new_n1132;
  assign new_n1134 = pd_2_ & new_n530;
  assign new_n1135 = ~pencrypt_mode_0_ & new_n1134;
  assign new_n1136 = ~new_n529 & new_n1135;
  assign new_n1137 = ~preset_0_ & new_n1136;
  assign new_n1138 = ~preset_0_ & pd_3_;
  assign new_n1139 = ~new_n512 & new_n1138;
  assign new_n1140 = ~new_n529 & new_n1139;
  assign new_n1141 = pinreg_22_ & new_n582;
  assign new_n1142 = new_n529 & new_n1141;
  assign new_n1143 = pinreg_30_ & new_n554;
  assign new_n1144 = new_n529 & new_n1143;
  assign new_n1145 = ~new_n1140 & ~new_n1142;
  assign new_n1146 = ~new_n1144 & new_n1145;
  assign new_n1147 = ~new_n1126 & ~new_n1130;
  assign new_n1148 = ~new_n1133 & ~new_n1137;
  assign new_n1149 = new_n1147 & new_n1148;
  assign pd_new_3_ = ~new_n1146 | ~new_n1149;
  assign new_n1151 = pinreg_43_ & new_n522;
  assign new_n1152 = pdata_41_ & ~new_n522;
  assign pdata_new_9_ = new_n1151 | new_n1152;
  assign new_n1154 = pinreg_19_ & new_n522;
  assign new_n1155 = pdata_44_ & ~new_n522;
  assign pdata_new_12_ = new_n1154 | new_n1155;
  assign new_n1157 = pinreg_47_ & new_n522;
  assign new_n1158 = pdata_57_ & ~new_n522;
  assign pdata_new_25_ = new_n1157 | new_n1158;
  assign new_n1160 = ~pcount_0_ & pinreg_8_;
  assign new_n1161 = ~new_n522 & new_n1160;
  assign new_n1162 = pinreg_0_ & pcount_0_;
  assign new_n1163 = ~new_n522 & new_n1162;
  assign pinreg_new_8_ = new_n1161 | new_n1163;
  assign new_n1165 = pcount_0_ & pinreg_9_;
  assign new_n1166 = ~new_n522 & new_n1165;
  assign new_n1167 = ~pcount_0_ & pinreg_17_;
  assign new_n1168 = ~new_n522 & new_n1167;
  assign pinreg_new_17_ = new_n1166 | new_n1168;
  assign new_n1170 = new_n655 & new_n731;
  assign new_n1171 = new_n655 & new_n733;
  assign new_n1172 = ~new_n652 & new_n720;
  assign new_n1173 = ~new_n655 & new_n1172;
  assign new_n1174 = new_n655 & new_n694;
  assign new_n1175 = ~new_n652 & new_n741;
  assign new_n1176 = ~new_n655 & new_n1175;
  assign new_n1177 = new_n655 & new_n705;
  assign new_n1178 = new_n652 & new_n680;
  assign new_n1179 = ~new_n655 & new_n1178;
  assign new_n1180 = new_n655 & new_n715;
  assign new_n1181 = ~new_n655 & new_n718;
  assign new_n1182 = ~new_n655 & new_n692;
  assign new_n1183 = ~new_n655 & new_n739;
  assign new_n1184 = new_n655 & new_n688;
  assign new_n1185 = new_n655 & new_n700;
  assign new_n1186 = ~new_n655 & new_n673;
  assign new_n1187 = ~new_n655 & new_n659;
  assign new_n1188 = new_n655 & new_n711;
  assign new_n1189 = ~new_n665 & ~new_n1188;
  assign new_n1190 = new_n745 & new_n1189;
  assign new_n1191 = ~new_n729 & ~new_n1187;
  assign new_n1192 = ~new_n730 & ~new_n1186;
  assign new_n1193 = new_n1191 & new_n1192;
  assign new_n1194 = new_n1190 & new_n1193;
  assign new_n1195 = ~new_n727 & ~new_n1185;
  assign new_n1196 = ~new_n719 & ~new_n1184;
  assign new_n1197 = new_n1195 & new_n1196;
  assign new_n1198 = ~new_n689 & ~new_n712;
  assign new_n1199 = new_n754 & new_n1198;
  assign new_n1200 = new_n1197 & new_n1199;
  assign new_n1201 = new_n1194 & new_n1200;
  assign new_n1202 = ~new_n710 & ~new_n1183;
  assign new_n1203 = ~new_n699 & ~new_n1182;
  assign new_n1204 = new_n1202 & new_n1203;
  assign new_n1205 = ~new_n1180 & ~new_n1181;
  assign new_n1206 = ~new_n1177 & ~new_n1179;
  assign new_n1207 = new_n1205 & new_n1206;
  assign new_n1208 = new_n1204 & new_n1207;
  assign new_n1209 = ~new_n674 & ~new_n1170;
  assign new_n1210 = ~new_n669 & ~new_n1171;
  assign new_n1211 = new_n1209 & new_n1210;
  assign new_n1212 = ~new_n679 & ~new_n1173;
  assign new_n1213 = ~new_n1174 & ~new_n1176;
  assign new_n1214 = new_n1212 & new_n1213;
  assign new_n1215 = new_n1211 & new_n1214;
  assign new_n1216 = new_n1208 & new_n1215;
  assign new_n1217 = new_n1201 & new_n1216;
  assign new_n1218 = pdata_31_ & new_n1217;
  assign new_n1219 = new_n522 & new_n1218;
  assign new_n1220 = ~pcount_0_ & poutreg_7_;
  assign new_n1221 = ~new_n522 & new_n1220;
  assign new_n1222 = ~pdata_31_ & ~new_n1217;
  assign new_n1223 = new_n522 & new_n1222;
  assign new_n1224 = pcount_0_ & poutreg_15_;
  assign new_n1225 = ~new_n522 & new_n1224;
  assign new_n1226 = ~new_n1219 & ~new_n1221;
  assign new_n1227 = ~new_n1223 & ~new_n1225;
  assign poutreg_new_7_ = ~new_n1226 | ~new_n1227;
  assign new_n1229 = pc_7_ & new_n535;
  assign new_n1230 = pencrypt_mode_0_ & new_n1229;
  assign new_n1231 = ~new_n529 & new_n1230;
  assign new_n1232 = ~preset_0_ & new_n1231;
  assign new_n1233 = pc_3_ & new_n535;
  assign new_n1234 = ~pencrypt_mode_0_ & new_n1233;
  assign new_n1235 = ~new_n529 & new_n1234;
  assign new_n1236 = ~preset_0_ & new_n1235;
  assign new_n1237 = pencrypt_mode_0_ & new_n786;
  assign new_n1238 = ~new_n529 & new_n1237;
  assign new_n1239 = ~preset_0_ & new_n1238;
  assign new_n1240 = pc_4_ & new_n530;
  assign new_n1241 = ~pencrypt_mode_0_ & new_n1240;
  assign new_n1242 = ~new_n529 & new_n1241;
  assign new_n1243 = ~preset_0_ & new_n1242;
  assign new_n1244 = ~preset_0_ & pc_5_;
  assign new_n1245 = ~new_n512 & new_n1244;
  assign new_n1246 = ~new_n529 & new_n1245;
  assign new_n1247 = pinreg_0_ & new_n582;
  assign new_n1248 = new_n529 & new_n1247;
  assign new_n1249 = pinreg_8_ & new_n554;
  assign new_n1250 = new_n529 & new_n1249;
  assign new_n1251 = ~new_n1246 & ~new_n1248;
  assign new_n1252 = ~new_n1250 & new_n1251;
  assign new_n1253 = ~new_n1232 & ~new_n1236;
  assign new_n1254 = ~new_n1239 & ~new_n1243;
  assign new_n1255 = new_n1253 & new_n1254;
  assign pc_new_5_ = ~new_n1252 | ~new_n1255;
  assign new_n1257 = pd_6_ & new_n535;
  assign new_n1258 = pencrypt_mode_0_ & new_n1257;
  assign new_n1259 = ~new_n529 & new_n1258;
  assign new_n1260 = ~preset_0_ & new_n1259;
  assign new_n1261 = pd_2_ & new_n535;
  assign new_n1262 = ~pencrypt_mode_0_ & new_n1261;
  assign new_n1263 = ~new_n529 & new_n1262;
  assign new_n1264 = ~preset_0_ & new_n1263;
  assign new_n1265 = pencrypt_mode_0_ & new_n815;
  assign new_n1266 = ~new_n529 & new_n1265;
  assign new_n1267 = ~preset_0_ & new_n1266;
  assign new_n1268 = pd_3_ & new_n530;
  assign new_n1269 = ~pencrypt_mode_0_ & new_n1268;
  assign new_n1270 = ~new_n529 & new_n1269;
  assign new_n1271 = ~preset_0_ & new_n1270;
  assign new_n1272 = ~preset_0_ & pd_4_;
  assign new_n1273 = ~new_n512 & new_n1272;
  assign new_n1274 = ~new_n529 & new_n1273;
  assign new_n1275 = pinreg_14_ & new_n582;
  assign new_n1276 = new_n529 & new_n1275;
  assign new_n1277 = pinreg_22_ & new_n554;
  assign new_n1278 = new_n529 & new_n1277;
  assign new_n1279 = ~new_n1274 & ~new_n1276;
  assign new_n1280 = ~new_n1278 & new_n1279;
  assign new_n1281 = ~new_n1260 & ~new_n1264;
  assign new_n1282 = ~new_n1267 & ~new_n1271;
  assign new_n1283 = new_n1281 & new_n1282;
  assign pd_new_4_ = ~new_n1280 | ~new_n1283;
  assign new_n1285 = pinreg_27_ & new_n522;
  assign new_n1286 = pdata_43_ & ~new_n522;
  assign pdata_new_11_ = new_n1285 | new_n1286;
  assign new_n1288 = pinreg_39_ & new_n522;
  assign new_n1289 = pdata_58_ & ~new_n522;
  assign pdata_new_26_ = new_n1288 | new_n1289;
  assign new_n1291 = ~pcount_0_ & pinreg_7_;
  assign new_n1292 = ~new_n522 & new_n1291;
  assign new_n1293 = pcount_0_ & pdata_in_7_;
  assign new_n1294 = ~new_n522 & new_n1293;
  assign pinreg_new_7_ = new_n1292 | new_n1294;
  assign new_n1296 = pcount_0_ & pinreg_8_;
  assign new_n1297 = ~new_n522 & new_n1296;
  assign new_n1298 = ~pcount_0_ & pinreg_16_;
  assign new_n1299 = ~new_n522 & new_n1298;
  assign pinreg_new_16_ = new_n1297 | new_n1299;
  assign new_n1301 = pcount_0_ & poutreg_16_;
  assign new_n1302 = ~new_n522 & new_n1301;
  assign new_n1303 = ~pcount_0_ & poutreg_8_;
  assign new_n1304 = ~new_n522 & new_n1303;
  assign new_n1305 = pdata_38_ & new_n522;
  assign new_n1306 = ~new_n1302 & ~new_n1304;
  assign poutreg_new_8_ = new_n1305 | ~new_n1306;
  assign new_n1308 = pencrypt_mode_0_ & new_n550;
  assign new_n1309 = ~new_n529 & new_n1308;
  assign new_n1310 = ~preset_0_ & new_n1309;
  assign new_n1311 = pc_0_ & new_n535;
  assign new_n1312 = ~pencrypt_mode_0_ & new_n1311;
  assign new_n1313 = ~new_n529 & new_n1312;
  assign new_n1314 = ~preset_0_ & new_n1313;
  assign new_n1315 = pencrypt_mode_0_ & new_n1106;
  assign new_n1316 = ~new_n529 & new_n1315;
  assign new_n1317 = ~preset_0_ & new_n1316;
  assign new_n1318 = pc_1_ & new_n530;
  assign new_n1319 = ~pencrypt_mode_0_ & new_n1318;
  assign new_n1320 = ~new_n529 & new_n1319;
  assign new_n1321 = ~preset_0_ & new_n1320;
  assign new_n1322 = ~preset_0_ & pc_2_;
  assign new_n1323 = ~new_n512 & new_n1322;
  assign new_n1324 = ~new_n529 & new_n1323;
  assign new_n1325 = pinreg_24_ & new_n582;
  assign new_n1326 = new_n529 & new_n1325;
  assign new_n1327 = pinreg_32_ & new_n554;
  assign new_n1328 = new_n529 & new_n1327;
  assign new_n1329 = ~new_n1324 & ~new_n1326;
  assign new_n1330 = ~new_n1328 & new_n1329;
  assign new_n1331 = ~new_n1310 & ~new_n1314;
  assign new_n1332 = ~new_n1317 & ~new_n1321;
  assign new_n1333 = new_n1331 & new_n1332;
  assign pc_new_2_ = ~new_n1330 | ~new_n1333;
  assign new_n1335 = pencrypt_mode_0_ & new_n597;
  assign new_n1336 = ~new_n529 & new_n1335;
  assign new_n1337 = ~preset_0_ & new_n1336;
  assign new_n1338 = pd_27_ & new_n535;
  assign new_n1339 = ~pencrypt_mode_0_ & new_n1338;
  assign new_n1340 = ~new_n529 & new_n1339;
  assign new_n1341 = ~preset_0_ & new_n1340;
  assign new_n1342 = pencrypt_mode_0_ & new_n1134;
  assign new_n1343 = ~new_n529 & new_n1342;
  assign new_n1344 = ~preset_0_ & new_n1343;
  assign new_n1345 = pd_0_ & new_n530;
  assign new_n1346 = ~pencrypt_mode_0_ & new_n1345;
  assign new_n1347 = ~new_n529 & new_n1346;
  assign new_n1348 = ~preset_0_ & new_n1347;
  assign new_n1349 = ~preset_0_ & pd_1_;
  assign new_n1350 = ~new_n512 & new_n1349;
  assign new_n1351 = ~new_n529 & new_n1350;
  assign new_n1352 = pinreg_38_ & new_n582;
  assign new_n1353 = new_n529 & new_n1352;
  assign new_n1354 = pinreg_46_ & new_n554;
  assign new_n1355 = new_n529 & new_n1354;
  assign new_n1356 = ~new_n1351 & ~new_n1353;
  assign new_n1357 = ~new_n1355 & new_n1356;
  assign new_n1358 = ~new_n1337 & ~new_n1341;
  assign new_n1359 = ~new_n1344 & ~new_n1348;
  assign new_n1360 = new_n1358 & new_n1359;
  assign pd_new_1_ = ~new_n1357 | ~new_n1360;
  assign new_n1362 = pinreg_35_ & new_n522;
  assign new_n1363 = pdata_42_ & ~new_n522;
  assign pdata_new_10_ = new_n1362 | new_n1363;
  assign new_n1365 = pd_7_ & ~pdata_62_;
  assign new_n1366 = ~pd_7_ & pdata_62_;
  assign new_n1367 = ~new_n1365 & ~new_n1366;
  assign new_n1368 = pd_0_ & ~pdata_63_;
  assign new_n1369 = ~pd_0_ & pdata_63_;
  assign new_n1370 = ~new_n1368 & ~new_n1369;
  assign new_n1371 = ~pdata_60_ & pd_13_;
  assign new_n1372 = pdata_60_ & ~pd_13_;
  assign new_n1373 = ~new_n1371 & ~new_n1372;
  assign new_n1374 = pd_21_ & ~pdata_61_;
  assign new_n1375 = ~pd_21_ & pdata_61_;
  assign new_n1376 = ~new_n1374 & ~new_n1375;
  assign new_n1377 = ~pdata_59_ & pd_17_;
  assign new_n1378 = pdata_59_ & ~pd_17_;
  assign new_n1379 = ~new_n1377 & ~new_n1378;
  assign new_n1380 = ~pdata_32_ & pd_3_;
  assign new_n1381 = pdata_32_ & ~pd_3_;
  assign new_n1382 = ~new_n1380 & ~new_n1381;
  assign new_n1383 = new_n1367 & new_n1370;
  assign new_n1384 = ~new_n1373 & new_n1383;
  assign new_n1385 = new_n1376 & new_n1384;
  assign new_n1386 = new_n1379 & new_n1385;
  assign new_n1387 = new_n1382 & new_n1386;
  assign new_n1388 = new_n1367 & ~new_n1370;
  assign new_n1389 = ~new_n1373 & new_n1388;
  assign new_n1390 = new_n1376 & new_n1389;
  assign new_n1391 = new_n1379 & new_n1390;
  assign new_n1392 = new_n1382 & new_n1391;
  assign new_n1393 = new_n1373 & new_n1388;
  assign new_n1394 = ~new_n1376 & new_n1393;
  assign new_n1395 = new_n1379 & new_n1394;
  assign new_n1396 = new_n1382 & new_n1395;
  assign new_n1397 = ~new_n1367 & new_n1370;
  assign new_n1398 = new_n1373 & new_n1397;
  assign new_n1399 = ~new_n1376 & new_n1398;
  assign new_n1400 = new_n1379 & new_n1399;
  assign new_n1401 = new_n1382 & new_n1400;
  assign new_n1402 = new_n1373 & new_n1383;
  assign new_n1403 = new_n1376 & new_n1402;
  assign new_n1404 = new_n1379 & new_n1403;
  assign new_n1405 = new_n1382 & new_n1404;
  assign new_n1406 = ~new_n1367 & ~new_n1370;
  assign new_n1407 = ~new_n1373 & new_n1406;
  assign new_n1408 = ~new_n1376 & new_n1407;
  assign new_n1409 = ~new_n1379 & new_n1408;
  assign new_n1410 = ~new_n1382 & new_n1409;
  assign new_n1411 = ~new_n1379 & new_n1394;
  assign new_n1412 = new_n1382 & new_n1411;
  assign new_n1413 = ~new_n1373 & new_n1397;
  assign new_n1414 = new_n1376 & new_n1413;
  assign new_n1415 = ~new_n1379 & new_n1414;
  assign new_n1416 = ~new_n1382 & new_n1415;
  assign new_n1417 = ~new_n1379 & new_n1399;
  assign new_n1418 = new_n1382 & new_n1417;
  assign new_n1419 = ~new_n1382 & new_n1417;
  assign new_n1420 = new_n1382 & new_n1415;
  assign new_n1421 = new_n1373 & new_n1406;
  assign new_n1422 = new_n1376 & new_n1421;
  assign new_n1423 = new_n1379 & new_n1422;
  assign new_n1424 = ~new_n1382 & new_n1423;
  assign new_n1425 = new_n1376 & new_n1407;
  assign new_n1426 = ~new_n1379 & new_n1425;
  assign new_n1427 = new_n1382 & new_n1426;
  assign new_n1428 = ~new_n1376 & new_n1421;
  assign new_n1429 = ~new_n1379 & new_n1428;
  assign new_n1430 = ~new_n1382 & new_n1429;
  assign new_n1431 = ~new_n1376 & new_n1389;
  assign new_n1432 = new_n1379 & new_n1431;
  assign new_n1433 = ~new_n1382 & new_n1432;
  assign new_n1434 = ~new_n1382 & new_n1411;
  assign new_n1435 = ~new_n1376 & new_n1413;
  assign new_n1436 = new_n1379 & new_n1435;
  assign new_n1437 = ~new_n1382 & new_n1436;
  assign new_n1438 = ~new_n1379 & new_n1390;
  assign new_n1439 = ~new_n1382 & new_n1438;
  assign new_n1440 = new_n1376 & new_n1393;
  assign new_n1441 = ~new_n1379 & new_n1440;
  assign new_n1442 = new_n1382 & new_n1441;
  assign new_n1443 = ~new_n1379 & new_n1385;
  assign new_n1444 = ~new_n1382 & new_n1443;
  assign new_n1445 = ~new_n1376 & new_n1402;
  assign new_n1446 = ~new_n1379 & new_n1445;
  assign new_n1447 = new_n1382 & new_n1446;
  assign new_n1448 = new_n1382 & new_n1409;
  assign new_n1449 = new_n1376 & new_n1398;
  assign new_n1450 = new_n1379 & new_n1449;
  assign new_n1451 = new_n1382 & new_n1450;
  assign new_n1452 = ~new_n1379 & new_n1449;
  assign new_n1453 = ~new_n1382 & new_n1452;
  assign new_n1454 = ~new_n1382 & new_n1386;
  assign new_n1455 = ~new_n1376 & new_n1384;
  assign new_n1456 = ~new_n1379 & new_n1455;
  assign new_n1457 = new_n1382 & new_n1456;
  assign new_n1458 = new_n1379 & new_n1425;
  assign new_n1459 = ~new_n1382 & new_n1458;
  assign new_n1460 = new_n1379 & new_n1445;
  assign new_n1461 = ~new_n1382 & new_n1460;
  assign new_n1462 = new_n1379 & new_n1440;
  assign new_n1463 = ~new_n1382 & new_n1462;
  assign new_n1464 = ~new_n1382 & new_n1450;
  assign new_n1465 = new_n1382 & new_n1458;
  assign new_n1466 = new_n1382 & new_n1436;
  assign new_n1467 = ~new_n1465 & ~new_n1466;
  assign new_n1468 = ~new_n1463 & ~new_n1464;
  assign new_n1469 = new_n1467 & new_n1468;
  assign new_n1470 = ~new_n1459 & ~new_n1461;
  assign new_n1471 = ~new_n1454 & ~new_n1457;
  assign new_n1472 = new_n1470 & new_n1471;
  assign new_n1473 = new_n1469 & new_n1472;
  assign new_n1474 = ~new_n1451 & ~new_n1453;
  assign new_n1475 = ~new_n1447 & ~new_n1448;
  assign new_n1476 = new_n1474 & new_n1475;
  assign new_n1477 = ~new_n1442 & ~new_n1444;
  assign new_n1478 = ~new_n1437 & ~new_n1439;
  assign new_n1479 = new_n1477 & new_n1478;
  assign new_n1480 = new_n1476 & new_n1479;
  assign new_n1481 = new_n1473 & new_n1480;
  assign new_n1482 = ~new_n1433 & ~new_n1434;
  assign new_n1483 = ~new_n1427 & ~new_n1430;
  assign new_n1484 = new_n1482 & new_n1483;
  assign new_n1485 = ~new_n1420 & ~new_n1424;
  assign new_n1486 = ~new_n1418 & ~new_n1419;
  assign new_n1487 = new_n1485 & new_n1486;
  assign new_n1488 = new_n1484 & new_n1487;
  assign new_n1489 = ~new_n1387 & ~new_n1392;
  assign new_n1490 = ~new_n1396 & ~new_n1401;
  assign new_n1491 = new_n1489 & new_n1490;
  assign new_n1492 = ~new_n1405 & ~new_n1410;
  assign new_n1493 = ~new_n1412 & ~new_n1416;
  assign new_n1494 = new_n1492 & new_n1493;
  assign new_n1495 = new_n1491 & new_n1494;
  assign new_n1496 = new_n1488 & new_n1495;
  assign new_n1497 = new_n1481 & new_n1496;
  assign new_n1498 = ~pdata_4_ & ~new_n1497;
  assign new_n1499 = ~new_n522 & new_n1498;
  assign new_n1500 = pdata_4_ & new_n1497;
  assign new_n1501 = ~new_n522 & new_n1500;
  assign new_n1502 = pinreg_16_ & new_n522;
  assign new_n1503 = ~new_n1499 & ~new_n1501;
  assign pdata_new_36_ = new_n1502 | ~new_n1503;
  assign new_n1505 = ~pcount_0_ & pinreg_2_;
  assign new_n1506 = ~new_n522 & new_n1505;
  assign new_n1507 = pcount_0_ & pdata_in_2_;
  assign new_n1508 = ~new_n522 & new_n1507;
  assign pinreg_new_2_ = new_n1506 | new_n1508;
  assign new_n1510 = pcount_0_ & pinreg_7_;
  assign new_n1511 = ~new_n522 & new_n1510;
  assign new_n1512 = ~pcount_0_ & pinreg_15_;
  assign new_n1513 = ~new_n522 & new_n1512;
  assign pinreg_new_15_ = new_n1511 | new_n1513;
  assign new_n1515 = ~pcount_0_ & poutreg_16_;
  assign new_n1516 = ~new_n522 & new_n1515;
  assign new_n1517 = pcount_0_ & poutreg_24_;
  assign new_n1518 = ~new_n522 & new_n1517;
  assign new_n1519 = pdata_37_ & new_n522;
  assign new_n1520 = ~new_n1516 & ~new_n1518;
  assign poutreg_new_16_ = new_n1519 | ~new_n1520;
  assign new_n1522 = pencrypt_mode_0_ & new_n803;
  assign new_n1523 = ~new_n529 & new_n1522;
  assign new_n1524 = ~preset_0_ & new_n1523;
  assign new_n1525 = pc_1_ & new_n535;
  assign new_n1526 = ~pencrypt_mode_0_ & new_n1525;
  assign new_n1527 = ~new_n529 & new_n1526;
  assign new_n1528 = ~preset_0_ & new_n1527;
  assign new_n1529 = pencrypt_mode_0_ & new_n1240;
  assign new_n1530 = ~new_n529 & new_n1529;
  assign new_n1531 = ~preset_0_ & new_n1530;
  assign new_n1532 = pc_2_ & new_n530;
  assign new_n1533 = ~pencrypt_mode_0_ & new_n1532;
  assign new_n1534 = ~new_n529 & new_n1533;
  assign new_n1535 = ~preset_0_ & new_n1534;
  assign new_n1536 = ~preset_0_ & pc_3_;
  assign new_n1537 = ~new_n512 & new_n1536;
  assign new_n1538 = ~new_n529 & new_n1537;
  assign new_n1539 = pinreg_16_ & new_n582;
  assign new_n1540 = new_n529 & new_n1539;
  assign new_n1541 = pinreg_24_ & new_n554;
  assign new_n1542 = new_n529 & new_n1541;
  assign new_n1543 = ~new_n1538 & ~new_n1540;
  assign new_n1544 = ~new_n1542 & new_n1543;
  assign new_n1545 = ~new_n1524 & ~new_n1528;
  assign new_n1546 = ~new_n1531 & ~new_n1535;
  assign new_n1547 = new_n1545 & new_n1546;
  assign pc_new_3_ = ~new_n1544 | ~new_n1547;
  assign new_n1549 = pencrypt_mode_0_ & new_n833;
  assign new_n1550 = ~new_n529 & new_n1549;
  assign new_n1551 = ~preset_0_ & new_n1550;
  assign new_n1552 = pd_0_ & new_n535;
  assign new_n1553 = ~pencrypt_mode_0_ & new_n1552;
  assign new_n1554 = ~new_n529 & new_n1553;
  assign new_n1555 = ~preset_0_ & new_n1554;
  assign new_n1556 = pencrypt_mode_0_ & new_n1268;
  assign new_n1557 = ~new_n529 & new_n1556;
  assign new_n1558 = ~preset_0_ & new_n1557;
  assign new_n1559 = pd_1_ & new_n530;
  assign new_n1560 = ~pencrypt_mode_0_ & new_n1559;
  assign new_n1561 = ~new_n529 & new_n1560;
  assign new_n1562 = ~preset_0_ & new_n1561;
  assign new_n1563 = ~preset_0_ & pd_2_;
  assign new_n1564 = ~new_n512 & new_n1563;
  assign new_n1565 = ~new_n529 & new_n1564;
  assign new_n1566 = pinreg_30_ & new_n582;
  assign new_n1567 = new_n529 & new_n1566;
  assign new_n1568 = pinreg_38_ & new_n554;
  assign new_n1569 = new_n529 & new_n1568;
  assign new_n1570 = ~new_n1565 & ~new_n1567;
  assign new_n1571 = ~new_n1569 & new_n1570;
  assign new_n1572 = ~new_n1551 & ~new_n1555;
  assign new_n1573 = ~new_n1558 & ~new_n1562;
  assign new_n1574 = new_n1572 & new_n1573;
  assign pd_new_2_ = ~new_n1571 | ~new_n1574;
  assign new_n1576 = pd_16_ & ~pdata_54_;
  assign new_n1577 = ~pd_16_ & pdata_54_;
  assign new_n1578 = ~new_n1576 & ~new_n1577;
  assign new_n1579 = pd_4_ & ~pdata_55_;
  assign new_n1580 = ~pd_4_ & pdata_55_;
  assign new_n1581 = ~new_n1579 & ~new_n1580;
  assign new_n1582 = pd_11_ & ~pdata_52_;
  assign new_n1583 = ~pd_11_ & pdata_52_;
  assign new_n1584 = ~new_n1582 & ~new_n1583;
  assign new_n1585 = pd_22_ & ~pdata_53_;
  assign new_n1586 = ~pd_22_ & pdata_53_;
  assign new_n1587 = ~new_n1585 & ~new_n1586;
  assign new_n1588 = pd_1_ & ~pdata_51_;
  assign new_n1589 = ~pd_1_ & pdata_51_;
  assign new_n1590 = ~new_n1588 & ~new_n1589;
  assign new_n1591 = pd_19_ & ~pdata_56_;
  assign new_n1592 = ~pd_19_ & pdata_56_;
  assign new_n1593 = ~new_n1591 & ~new_n1592;
  assign new_n1594 = new_n1578 & new_n1581;
  assign new_n1595 = new_n1584 & new_n1594;
  assign new_n1596 = ~new_n1587 & new_n1595;
  assign new_n1597 = new_n1590 & new_n1596;
  assign new_n1598 = new_n1593 & new_n1597;
  assign new_n1599 = new_n1578 & ~new_n1581;
  assign new_n1600 = ~new_n1584 & new_n1599;
  assign new_n1601 = new_n1587 & new_n1600;
  assign new_n1602 = new_n1590 & new_n1601;
  assign new_n1603 = new_n1593 & new_n1602;
  assign new_n1604 = ~new_n1578 & new_n1581;
  assign new_n1605 = new_n1584 & new_n1604;
  assign new_n1606 = new_n1587 & new_n1605;
  assign new_n1607 = new_n1590 & new_n1606;
  assign new_n1608 = new_n1593 & new_n1607;
  assign new_n1609 = ~new_n1578 & ~new_n1581;
  assign new_n1610 = new_n1584 & new_n1609;
  assign new_n1611 = new_n1587 & new_n1610;
  assign new_n1612 = new_n1590 & new_n1611;
  assign new_n1613 = new_n1593 & new_n1612;
  assign new_n1614 = new_n1587 & new_n1595;
  assign new_n1615 = new_n1590 & new_n1614;
  assign new_n1616 = new_n1593 & new_n1615;
  assign new_n1617 = ~new_n1584 & new_n1609;
  assign new_n1618 = ~new_n1587 & new_n1617;
  assign new_n1619 = ~new_n1590 & new_n1618;
  assign new_n1620 = ~new_n1593 & new_n1619;
  assign new_n1621 = ~new_n1590 & new_n1606;
  assign new_n1622 = new_n1593 & new_n1621;
  assign new_n1623 = ~new_n1590 & new_n1601;
  assign new_n1624 = ~new_n1593 & new_n1623;
  assign new_n1625 = ~new_n1587 & new_n1605;
  assign new_n1626 = ~new_n1590 & new_n1625;
  assign new_n1627 = new_n1593 & new_n1626;
  assign new_n1628 = ~new_n1584 & new_n1604;
  assign new_n1629 = ~new_n1587 & new_n1628;
  assign new_n1630 = ~new_n1590 & new_n1629;
  assign new_n1631 = ~new_n1593 & new_n1630;
  assign new_n1632 = new_n1587 & new_n1617;
  assign new_n1633 = ~new_n1590 & new_n1632;
  assign new_n1634 = new_n1593 & new_n1633;
  assign new_n1635 = new_n1590 & new_n1618;
  assign new_n1636 = ~new_n1593 & new_n1635;
  assign new_n1637 = ~new_n1587 & new_n1600;
  assign new_n1638 = ~new_n1590 & new_n1637;
  assign new_n1639 = new_n1593 & new_n1638;
  assign new_n1640 = ~new_n1593 & new_n1626;
  assign new_n1641 = new_n1590 & new_n1632;
  assign new_n1642 = ~new_n1593 & new_n1641;
  assign new_n1643 = ~new_n1590 & new_n1596;
  assign new_n1644 = ~new_n1593 & new_n1643;
  assign new_n1645 = new_n1590 & new_n1637;
  assign new_n1646 = ~new_n1593 & new_n1645;
  assign new_n1647 = ~new_n1584 & new_n1594;
  assign new_n1648 = new_n1587 & new_n1647;
  assign new_n1649 = ~new_n1590 & new_n1648;
  assign new_n1650 = ~new_n1593 & new_n1649;
  assign new_n1651 = ~new_n1590 & new_n1614;
  assign new_n1652 = new_n1593 & new_n1651;
  assign new_n1653 = ~new_n1587 & new_n1610;
  assign new_n1654 = ~new_n1590 & new_n1653;
  assign new_n1655 = ~new_n1593 & new_n1654;
  assign new_n1656 = new_n1584 & new_n1599;
  assign new_n1657 = new_n1587 & new_n1656;
  assign new_n1658 = ~new_n1590 & new_n1657;
  assign new_n1659 = new_n1593 & new_n1658;
  assign new_n1660 = new_n1590 & new_n1653;
  assign new_n1661 = new_n1593 & new_n1660;
  assign new_n1662 = ~new_n1587 & new_n1656;
  assign new_n1663 = ~new_n1590 & new_n1662;
  assign new_n1664 = new_n1593 & new_n1663;
  assign new_n1665 = ~new_n1590 & new_n1611;
  assign new_n1666 = ~new_n1593 & new_n1665;
  assign new_n1667 = new_n1590 & new_n1625;
  assign new_n1668 = ~new_n1593 & new_n1667;
  assign new_n1669 = new_n1593 & new_n1630;
  assign new_n1670 = new_n1587 & new_n1628;
  assign new_n1671 = new_n1590 & new_n1670;
  assign new_n1672 = ~new_n1593 & new_n1671;
  assign new_n1673 = new_n1590 & new_n1662;
  assign new_n1674 = ~new_n1593 & new_n1673;
  assign new_n1675 = ~new_n1593 & new_n1615;
  assign new_n1676 = new_n1590 & new_n1657;
  assign new_n1677 = ~new_n1593 & new_n1676;
  assign new_n1678 = ~new_n1587 & new_n1647;
  assign new_n1679 = new_n1590 & new_n1678;
  assign new_n1680 = new_n1593 & new_n1679;
  assign new_n1681 = new_n1593 & new_n1635;
  assign new_n1682 = ~new_n1680 & ~new_n1681;
  assign new_n1683 = ~new_n1675 & ~new_n1677;
  assign new_n1684 = new_n1682 & new_n1683;
  assign new_n1685 = ~new_n1672 & ~new_n1674;
  assign new_n1686 = ~new_n1668 & ~new_n1669;
  assign new_n1687 = new_n1685 & new_n1686;
  assign new_n1688 = new_n1684 & new_n1687;
  assign new_n1689 = ~new_n1664 & ~new_n1666;
  assign new_n1690 = ~new_n1659 & ~new_n1661;
  assign new_n1691 = new_n1689 & new_n1690;
  assign new_n1692 = ~new_n1652 & ~new_n1655;
  assign new_n1693 = ~new_n1646 & ~new_n1650;
  assign new_n1694 = new_n1692 & new_n1693;
  assign new_n1695 = new_n1691 & new_n1694;
  assign new_n1696 = new_n1688 & new_n1695;
  assign new_n1697 = ~new_n1642 & ~new_n1644;
  assign new_n1698 = ~new_n1639 & ~new_n1640;
  assign new_n1699 = new_n1697 & new_n1698;
  assign new_n1700 = ~new_n1634 & ~new_n1636;
  assign new_n1701 = ~new_n1627 & ~new_n1631;
  assign new_n1702 = new_n1700 & new_n1701;
  assign new_n1703 = new_n1699 & new_n1702;
  assign new_n1704 = ~new_n1598 & ~new_n1603;
  assign new_n1705 = ~new_n1608 & ~new_n1613;
  assign new_n1706 = new_n1704 & new_n1705;
  assign new_n1707 = ~new_n1616 & ~new_n1620;
  assign new_n1708 = ~new_n1622 & ~new_n1624;
  assign new_n1709 = new_n1707 & new_n1708;
  assign new_n1710 = new_n1706 & new_n1709;
  assign new_n1711 = new_n1703 & new_n1710;
  assign new_n1712 = new_n1696 & new_n1711;
  assign new_n1713 = ~pdata_3_ & ~new_n1712;
  assign new_n1714 = ~new_n522 & new_n1713;
  assign new_n1715 = pdata_3_ & new_n1712;
  assign new_n1716 = ~new_n522 & new_n1715;
  assign new_n1717 = pinreg_24_ & new_n522;
  assign new_n1718 = ~new_n1714 & ~new_n1716;
  assign pdata_new_35_ = new_n1717 | ~new_n1718;
  assign new_n1720 = pinreg_1_ & ~pcount_0_;
  assign new_n1721 = ~new_n522 & new_n1720;
  assign new_n1722 = pcount_0_ & pdata_in_1_;
  assign new_n1723 = ~new_n522 & new_n1722;
  assign pinreg_new_1_ = new_n1721 | new_n1723;
  assign new_n1725 = pcount_0_ & pinreg_6_;
  assign new_n1726 = ~new_n522 & new_n1725;
  assign new_n1727 = ~pcount_0_ & pinreg_14_;
  assign new_n1728 = ~new_n522 & new_n1727;
  assign pinreg_new_14_ = new_n1726 | new_n1728;
  assign new_n1730 = ~pdata_34_ & pc_23_;
  assign new_n1731 = pdata_34_ & ~pc_23_;
  assign new_n1732 = ~new_n1730 & ~new_n1731;
  assign new_n1733 = ~pdata_35_ & pc_0_;
  assign new_n1734 = pdata_35_ & ~pc_0_;
  assign new_n1735 = ~new_n1733 & ~new_n1734;
  assign new_n1736 = ~pdata_32_ & pc_16_;
  assign new_n1737 = pdata_32_ & ~pc_16_;
  assign new_n1738 = ~new_n1736 & ~new_n1737;
  assign new_n1739 = ~pdata_33_ & pc_10_;
  assign new_n1740 = pdata_33_ & ~pc_10_;
  assign new_n1741 = ~new_n1739 & ~new_n1740;
  assign new_n1742 = pc_13_ & ~pdata_63_;
  assign new_n1743 = ~pc_13_ & pdata_63_;
  assign new_n1744 = ~new_n1742 & ~new_n1743;
  assign new_n1745 = ~pdata_36_ & pc_4_;
  assign new_n1746 = pdata_36_ & ~pc_4_;
  assign new_n1747 = ~new_n1745 & ~new_n1746;
  assign new_n1748 = new_n1732 & ~new_n1735;
  assign new_n1749 = new_n1738 & new_n1748;
  assign new_n1750 = new_n1741 & new_n1749;
  assign new_n1751 = new_n1744 & new_n1750;
  assign new_n1752 = ~new_n1747 & new_n1751;
  assign new_n1753 = ~new_n1732 & new_n1735;
  assign new_n1754 = new_n1738 & new_n1753;
  assign new_n1755 = new_n1741 & new_n1754;
  assign new_n1756 = new_n1744 & new_n1755;
  assign new_n1757 = ~new_n1747 & new_n1756;
  assign new_n1758 = ~new_n1738 & new_n1748;
  assign new_n1759 = ~new_n1741 & new_n1758;
  assign new_n1760 = new_n1744 & new_n1759;
  assign new_n1761 = new_n1747 & new_n1760;
  assign new_n1762 = ~new_n1732 & ~new_n1735;
  assign new_n1763 = ~new_n1738 & new_n1762;
  assign new_n1764 = ~new_n1741 & new_n1763;
  assign new_n1765 = new_n1744 & new_n1764;
  assign new_n1766 = new_n1747 & new_n1765;
  assign new_n1767 = new_n1732 & new_n1735;
  assign new_n1768 = ~new_n1738 & new_n1767;
  assign new_n1769 = ~new_n1741 & new_n1768;
  assign new_n1770 = new_n1744 & new_n1769;
  assign new_n1771 = new_n1747 & new_n1770;
  assign new_n1772 = new_n1741 & new_n1768;
  assign new_n1773 = new_n1744 & new_n1772;
  assign new_n1774 = new_n1747 & new_n1773;
  assign new_n1775 = ~new_n1744 & new_n1769;
  assign new_n1776 = new_n1747 & new_n1775;
  assign new_n1777 = ~new_n1741 & new_n1754;
  assign new_n1778 = new_n1744 & new_n1777;
  assign new_n1779 = new_n1747 & new_n1778;
  assign new_n1780 = ~new_n1738 & new_n1753;
  assign new_n1781 = ~new_n1741 & new_n1780;
  assign new_n1782 = ~new_n1744 & new_n1781;
  assign new_n1783 = new_n1747 & new_n1782;
  assign new_n1784 = ~new_n1744 & new_n1777;
  assign new_n1785 = ~new_n1747 & new_n1784;
  assign new_n1786 = new_n1738 & new_n1767;
  assign new_n1787 = new_n1741 & new_n1786;
  assign new_n1788 = ~new_n1744 & new_n1787;
  assign new_n1789 = ~new_n1747 & new_n1788;
  assign new_n1790 = new_n1738 & new_n1762;
  assign new_n1791 = ~new_n1741 & new_n1790;
  assign new_n1792 = new_n1744 & new_n1791;
  assign new_n1793 = ~new_n1747 & new_n1792;
  assign new_n1794 = ~new_n1741 & new_n1749;
  assign new_n1795 = ~new_n1744 & new_n1794;
  assign new_n1796 = ~new_n1747 & new_n1795;
  assign new_n1797 = new_n1741 & new_n1780;
  assign new_n1798 = ~new_n1744 & new_n1797;
  assign new_n1799 = ~new_n1747 & new_n1798;
  assign new_n1800 = ~new_n1744 & new_n1791;
  assign new_n1801 = new_n1747 & new_n1800;
  assign new_n1802 = new_n1741 & new_n1758;
  assign new_n1803 = ~new_n1744 & new_n1802;
  assign new_n1804 = ~new_n1747 & new_n1803;
  assign new_n1805 = ~new_n1744 & new_n1772;
  assign new_n1806 = new_n1747 & new_n1805;
  assign new_n1807 = ~new_n1744 & new_n1764;
  assign new_n1808 = ~new_n1747 & new_n1807;
  assign new_n1809 = new_n1747 & new_n1798;
  assign new_n1810 = new_n1744 & new_n1794;
  assign new_n1811 = new_n1747 & new_n1810;
  assign new_n1812 = new_n1741 & new_n1763;
  assign new_n1813 = ~new_n1744 & new_n1812;
  assign new_n1814 = new_n1747 & new_n1813;
  assign new_n1815 = new_n1741 & new_n1790;
  assign new_n1816 = new_n1744 & new_n1815;
  assign new_n1817 = new_n1747 & new_n1816;
  assign new_n1818 = ~new_n1744 & new_n1750;
  assign new_n1819 = new_n1747 & new_n1818;
  assign new_n1820 = ~new_n1747 & new_n1805;
  assign new_n1821 = new_n1744 & new_n1781;
  assign new_n1822 = ~new_n1747 & new_n1821;
  assign new_n1823 = ~new_n1747 & new_n1800;
  assign new_n1824 = ~new_n1741 & new_n1786;
  assign new_n1825 = ~new_n1744 & new_n1824;
  assign new_n1826 = new_n1747 & new_n1825;
  assign new_n1827 = new_n1747 & new_n1756;
  assign new_n1828 = ~new_n1747 & new_n1770;
  assign new_n1829 = ~new_n1747 & new_n1760;
  assign new_n1830 = ~new_n1747 & new_n1778;
  assign new_n1831 = new_n1744 & new_n1812;
  assign new_n1832 = ~new_n1747 & new_n1831;
  assign new_n1833 = ~new_n1830 & ~new_n1832;
  assign new_n1834 = ~new_n1828 & ~new_n1829;
  assign new_n1835 = new_n1833 & new_n1834;
  assign new_n1836 = ~new_n1826 & ~new_n1827;
  assign new_n1837 = ~new_n1822 & ~new_n1823;
  assign new_n1838 = new_n1836 & new_n1837;
  assign new_n1839 = new_n1835 & new_n1838;
  assign new_n1840 = ~new_n1819 & ~new_n1820;
  assign new_n1841 = ~new_n1814 & ~new_n1817;
  assign new_n1842 = new_n1840 & new_n1841;
  assign new_n1843 = ~new_n1809 & ~new_n1811;
  assign new_n1844 = ~new_n1806 & ~new_n1808;
  assign new_n1845 = new_n1843 & new_n1844;
  assign new_n1846 = new_n1842 & new_n1845;
  assign new_n1847 = new_n1839 & new_n1846;
  assign new_n1848 = ~new_n1801 & ~new_n1804;
  assign new_n1849 = ~new_n1796 & ~new_n1799;
  assign new_n1850 = new_n1848 & new_n1849;
  assign new_n1851 = ~new_n1789 & ~new_n1793;
  assign new_n1852 = ~new_n1783 & ~new_n1785;
  assign new_n1853 = new_n1851 & new_n1852;
  assign new_n1854 = new_n1850 & new_n1853;
  assign new_n1855 = ~new_n1752 & ~new_n1757;
  assign new_n1856 = ~new_n1761 & ~new_n1766;
  assign new_n1857 = new_n1855 & new_n1856;
  assign new_n1858 = ~new_n1771 & ~new_n1774;
  assign new_n1859 = ~new_n1776 & ~new_n1779;
  assign new_n1860 = new_n1858 & new_n1859;
  assign new_n1861 = new_n1857 & new_n1860;
  assign new_n1862 = new_n1854 & new_n1861;
  assign new_n1863 = new_n1847 & new_n1862;
  assign new_n1864 = pdata_30_ & new_n1863;
  assign new_n1865 = new_n522 & new_n1864;
  assign new_n1866 = pcount_0_ & poutreg_23_;
  assign new_n1867 = ~new_n522 & new_n1866;
  assign new_n1868 = ~pdata_30_ & ~new_n1863;
  assign new_n1869 = new_n522 & new_n1868;
  assign new_n1870 = ~pcount_0_ & poutreg_15_;
  assign new_n1871 = ~new_n522 & new_n1870;
  assign new_n1872 = ~new_n1865 & ~new_n1867;
  assign new_n1873 = ~new_n1869 & ~new_n1871;
  assign poutreg_new_15_ = ~new_n1872 | ~new_n1873;
  assign new_n1875 = pencrypt_mode_0_ & new_n1099;
  assign new_n1876 = ~new_n529 & new_n1875;
  assign new_n1877 = ~preset_0_ & new_n1876;
  assign new_n1878 = pc_26_ & new_n535;
  assign new_n1879 = ~pencrypt_mode_0_ & new_n1878;
  assign new_n1880 = ~new_n529 & new_n1879;
  assign new_n1881 = ~preset_0_ & new_n1880;
  assign new_n1882 = pencrypt_mode_0_ & new_n1318;
  assign new_n1883 = ~new_n529 & new_n1882;
  assign new_n1884 = ~preset_0_ & new_n1883;
  assign new_n1885 = pc_27_ & new_n530;
  assign new_n1886 = ~pencrypt_mode_0_ & new_n1885;
  assign new_n1887 = ~new_n529 & new_n1886;
  assign new_n1888 = ~preset_0_ & new_n1887;
  assign new_n1889 = ~preset_0_ & pc_0_;
  assign new_n1890 = ~new_n512 & new_n1889;
  assign new_n1891 = ~new_n529 & new_n1890;
  assign new_n1892 = pinreg_40_ & new_n582;
  assign new_n1893 = new_n529 & new_n1892;
  assign new_n1894 = pinreg_48_ & new_n554;
  assign new_n1895 = new_n529 & new_n1894;
  assign new_n1896 = ~new_n1891 & ~new_n1893;
  assign new_n1897 = ~new_n1895 & new_n1896;
  assign new_n1898 = ~new_n1877 & ~new_n1881;
  assign new_n1899 = ~new_n1884 & ~new_n1888;
  assign new_n1900 = new_n1898 & new_n1899;
  assign pc_new_0_ = ~new_n1897 | ~new_n1900;
  assign new_n1902 = pinreg_15_ & new_n522;
  assign new_n1903 = pdata_61_ & ~new_n522;
  assign pdata_new_29_ = new_n1902 | new_n1903;
  assign new_n1905 = ~new_n522 & new_n779;
  assign new_n1906 = ~new_n522 & new_n775;
  assign new_n1907 = pinreg_0_ & new_n522;
  assign new_n1908 = ~new_n1905 & ~new_n1906;
  assign pdata_new_38_ = new_n1907 | ~new_n1908;
  assign new_n1910 = ~pcount_0_ & pinreg_4_;
  assign new_n1911 = ~new_n522 & new_n1910;
  assign new_n1912 = pcount_0_ & pdata_in_4_;
  assign new_n1913 = ~new_n522 & new_n1912;
  assign pinreg_new_4_ = new_n1911 | new_n1913;
  assign new_n1915 = pcount_0_ & pinreg_5_;
  assign new_n1916 = ~new_n522 & new_n1915;
  assign new_n1917 = ~pcount_0_ & pinreg_13_;
  assign new_n1918 = ~new_n522 & new_n1917;
  assign pinreg_new_13_ = new_n1916 | new_n1918;
  assign new_n1920 = ~pcount_0_ & poutreg_18_;
  assign new_n1921 = ~new_n522 & new_n1920;
  assign new_n1922 = pcount_0_ & poutreg_26_;
  assign new_n1923 = ~new_n522 & new_n1922;
  assign new_n1924 = pdata_45_ & new_n522;
  assign new_n1925 = ~new_n1921 & ~new_n1923;
  assign poutreg_new_18_ = new_n1924 | ~new_n1925;
  assign new_n1927 = pencrypt_mode_0_ & new_n1233;
  assign new_n1928 = ~new_n529 & new_n1927;
  assign new_n1929 = ~preset_0_ & new_n1928;
  assign new_n1930 = pc_27_ & new_n535;
  assign new_n1931 = ~pencrypt_mode_0_ & new_n1930;
  assign new_n1932 = ~new_n529 & new_n1931;
  assign new_n1933 = ~preset_0_ & new_n1932;
  assign new_n1934 = pencrypt_mode_0_ & new_n1532;
  assign new_n1935 = ~new_n529 & new_n1934;
  assign new_n1936 = ~preset_0_ & new_n1935;
  assign new_n1937 = pc_0_ & new_n530;
  assign new_n1938 = ~pencrypt_mode_0_ & new_n1937;
  assign new_n1939 = ~new_n529 & new_n1938;
  assign new_n1940 = ~preset_0_ & new_n1939;
  assign new_n1941 = ~preset_0_ & pc_1_;
  assign new_n1942 = ~new_n512 & new_n1941;
  assign new_n1943 = ~new_n529 & new_n1942;
  assign new_n1944 = pinreg_32_ & new_n582;
  assign new_n1945 = new_n529 & new_n1944;
  assign new_n1946 = pinreg_40_ & new_n554;
  assign new_n1947 = new_n529 & new_n1946;
  assign new_n1948 = ~new_n1943 & ~new_n1945;
  assign new_n1949 = ~new_n1947 & new_n1948;
  assign new_n1950 = ~new_n1929 & ~new_n1933;
  assign new_n1951 = ~new_n1936 & ~new_n1940;
  assign new_n1952 = new_n1950 & new_n1951;
  assign pc_new_1_ = ~new_n1949 | ~new_n1952;
  assign new_n1954 = pencrypt_mode_0_ & new_n1261;
  assign new_n1955 = ~new_n529 & new_n1954;
  assign new_n1956 = ~preset_0_ & new_n1955;
  assign new_n1957 = pd_26_ & new_n535;
  assign new_n1958 = ~pencrypt_mode_0_ & new_n1957;
  assign new_n1959 = ~new_n529 & new_n1958;
  assign new_n1960 = ~preset_0_ & new_n1959;
  assign new_n1961 = pencrypt_mode_0_ & new_n1559;
  assign new_n1962 = ~new_n529 & new_n1961;
  assign new_n1963 = ~preset_0_ & new_n1962;
  assign new_n1964 = pd_27_ & new_n530;
  assign new_n1965 = ~pencrypt_mode_0_ & new_n1964;
  assign new_n1966 = ~new_n529 & new_n1965;
  assign new_n1967 = ~preset_0_ & new_n1966;
  assign new_n1968 = ~preset_0_ & pd_0_;
  assign new_n1969 = ~new_n512 & new_n1968;
  assign new_n1970 = ~new_n529 & new_n1969;
  assign new_n1971 = pinreg_46_ & new_n582;
  assign new_n1972 = new_n529 & new_n1971;
  assign new_n1973 = pinreg_54_ & new_n554;
  assign new_n1974 = new_n529 & new_n1973;
  assign new_n1975 = ~new_n1970 & ~new_n1972;
  assign new_n1976 = ~new_n1974 & new_n1975;
  assign new_n1977 = ~new_n1956 & ~new_n1960;
  assign new_n1978 = ~new_n1963 & ~new_n1967;
  assign new_n1979 = new_n1977 & new_n1978;
  assign pd_new_0_ = ~new_n1976 | ~new_n1979;
  assign new_n1981 = ~pdata_42_ & pc_3_;
  assign new_n1982 = pdata_42_ & ~pc_3_;
  assign new_n1983 = ~new_n1981 & ~new_n1982;
  assign new_n1984 = ~pdata_43_ & pc_25_;
  assign new_n1985 = pdata_43_ & ~pc_25_;
  assign new_n1986 = ~new_n1984 & ~new_n1985;
  assign new_n1987 = ~pdata_40_ & pc_18_;
  assign new_n1988 = pdata_40_ & ~pc_18_;
  assign new_n1989 = ~new_n1987 & ~new_n1988;
  assign new_n1990 = ~pdata_41_ & pc_11_;
  assign new_n1991 = pdata_41_ & ~pc_11_;
  assign new_n1992 = ~new_n1990 & ~new_n1991;
  assign new_n1993 = pc_22_ & ~pdata_39_;
  assign new_n1994 = ~pc_22_ & pdata_39_;
  assign new_n1995 = ~new_n1993 & ~new_n1994;
  assign new_n1996 = ~pdata_44_ & pc_7_;
  assign new_n1997 = pdata_44_ & ~pc_7_;
  assign new_n1998 = ~new_n1996 & ~new_n1997;
  assign new_n1999 = ~new_n1983 & ~new_n1986;
  assign new_n2000 = new_n1989 & new_n1999;
  assign new_n2001 = ~new_n1992 & new_n2000;
  assign new_n2002 = new_n1995 & new_n2001;
  assign new_n2003 = new_n1998 & new_n2002;
  assign new_n2004 = new_n1983 & ~new_n1986;
  assign new_n2005 = ~new_n1989 & new_n2004;
  assign new_n2006 = new_n1992 & new_n2005;
  assign new_n2007 = new_n1995 & new_n2006;
  assign new_n2008 = new_n1998 & new_n2007;
  assign new_n2009 = new_n1989 & new_n2004;
  assign new_n2010 = ~new_n1992 & new_n2009;
  assign new_n2011 = new_n1995 & new_n2010;
  assign new_n2012 = new_n1998 & new_n2011;
  assign new_n2013 = ~new_n1983 & new_n1986;
  assign new_n2014 = new_n1989 & new_n2013;
  assign new_n2015 = ~new_n1992 & new_n2014;
  assign new_n2016 = new_n1995 & new_n2015;
  assign new_n2017 = new_n1998 & new_n2016;
  assign new_n2018 = new_n1992 & new_n2014;
  assign new_n2019 = new_n1995 & new_n2018;
  assign new_n2020 = new_n1998 & new_n2019;
  assign new_n2021 = ~new_n1992 & new_n2005;
  assign new_n2022 = ~new_n1995 & new_n2021;
  assign new_n2023 = ~new_n1998 & new_n2022;
  assign new_n2024 = ~new_n1995 & new_n2010;
  assign new_n2025 = new_n1998 & new_n2024;
  assign new_n2026 = new_n1983 & new_n1986;
  assign new_n2027 = ~new_n1989 & new_n2026;
  assign new_n2028 = ~new_n1992 & new_n2027;
  assign new_n2029 = ~new_n1995 & new_n2028;
  assign new_n2030 = ~new_n1998 & new_n2029;
  assign new_n2031 = ~new_n1995 & new_n2015;
  assign new_n2032 = new_n1998 & new_n2031;
  assign new_n2033 = new_n1989 & new_n2026;
  assign new_n2034 = new_n1992 & new_n2033;
  assign new_n2035 = ~new_n1995 & new_n2034;
  assign new_n2036 = ~new_n1998 & new_n2035;
  assign new_n2037 = new_n1992 & new_n2027;
  assign new_n2038 = ~new_n1995 & new_n2037;
  assign new_n2039 = new_n1998 & new_n2038;
  assign new_n2040 = ~new_n1989 & new_n1999;
  assign new_n2041 = ~new_n1992 & new_n2040;
  assign new_n2042 = new_n1995 & new_n2041;
  assign new_n2043 = ~new_n1998 & new_n2042;
  assign new_n2044 = new_n1998 & new_n2029;
  assign new_n2045 = ~new_n1995 & new_n2001;
  assign new_n2046 = ~new_n1998 & new_n2045;
  assign new_n2047 = new_n1995 & new_n2021;
  assign new_n2048 = ~new_n1998 & new_n2047;
  assign new_n2049 = ~new_n1998 & new_n2024;
  assign new_n2050 = ~new_n1989 & new_n2013;
  assign new_n2051 = ~new_n1992 & new_n2050;
  assign new_n2052 = new_n1995 & new_n2051;
  assign new_n2053 = ~new_n1998 & new_n2052;
  assign new_n2054 = new_n1992 & new_n2040;
  assign new_n2055 = ~new_n1995 & new_n2054;
  assign new_n2056 = ~new_n1998 & new_n2055;
  assign new_n2057 = new_n1998 & new_n2035;
  assign new_n2058 = ~new_n1995 & new_n2006;
  assign new_n2059 = ~new_n1998 & new_n2058;
  assign new_n2060 = new_n1992 & new_n2000;
  assign new_n2061 = ~new_n1995 & new_n2060;
  assign new_n2062 = new_n1998 & new_n2061;
  assign new_n2063 = new_n1998 & new_n2058;
  assign new_n2064 = new_n1995 & new_n2037;
  assign new_n2065 = new_n1998 & new_n2064;
  assign new_n2066 = ~new_n1995 & new_n2018;
  assign new_n2067 = ~new_n1998 & new_n2066;
  assign new_n2068 = ~new_n1992 & new_n2033;
  assign new_n2069 = new_n1995 & new_n2068;
  assign new_n2070 = ~new_n1998 & new_n2069;
  assign new_n2071 = ~new_n1995 & new_n2041;
  assign new_n2072 = new_n1998 & new_n2071;
  assign new_n2073 = new_n1992 & new_n2050;
  assign new_n2074 = new_n1995 & new_n2073;
  assign new_n2075 = ~new_n1998 & new_n2074;
  assign new_n2076 = new_n1995 & new_n2060;
  assign new_n2077 = ~new_n1998 & new_n2076;
  assign new_n2078 = new_n1995 & new_n2034;
  assign new_n2079 = ~new_n1998 & new_n2078;
  assign new_n2080 = new_n1992 & new_n2009;
  assign new_n2081 = new_n1995 & new_n2080;
  assign new_n2082 = ~new_n1998 & new_n2081;
  assign new_n2083 = new_n1995 & new_n2054;
  assign new_n2084 = new_n1998 & new_n2083;
  assign new_n2085 = new_n1995 & new_n2028;
  assign new_n2086 = new_n1998 & new_n2085;
  assign new_n2087 = ~new_n2084 & ~new_n2086;
  assign new_n2088 = ~new_n2079 & ~new_n2082;
  assign new_n2089 = new_n2087 & new_n2088;
  assign new_n2090 = ~new_n2075 & ~new_n2077;
  assign new_n2091 = ~new_n2070 & ~new_n2072;
  assign new_n2092 = new_n2090 & new_n2091;
  assign new_n2093 = new_n2089 & new_n2092;
  assign new_n2094 = ~new_n2065 & ~new_n2067;
  assign new_n2095 = ~new_n2062 & ~new_n2063;
  assign new_n2096 = new_n2094 & new_n2095;
  assign new_n2097 = ~new_n2057 & ~new_n2059;
  assign new_n2098 = ~new_n2053 & ~new_n2056;
  assign new_n2099 = new_n2097 & new_n2098;
  assign new_n2100 = new_n2096 & new_n2099;
  assign new_n2101 = new_n2093 & new_n2100;
  assign new_n2102 = ~new_n2048 & ~new_n2049;
  assign new_n2103 = ~new_n2044 & ~new_n2046;
  assign new_n2104 = new_n2102 & new_n2103;
  assign new_n2105 = ~new_n2039 & ~new_n2043;
  assign new_n2106 = ~new_n2032 & ~new_n2036;
  assign new_n2107 = new_n2105 & new_n2106;
  assign new_n2108 = new_n2104 & new_n2107;
  assign new_n2109 = ~new_n2003 & ~new_n2008;
  assign new_n2110 = ~new_n2012 & ~new_n2017;
  assign new_n2111 = new_n2109 & new_n2110;
  assign new_n2112 = ~new_n2020 & ~new_n2023;
  assign new_n2113 = ~new_n2025 & ~new_n2030;
  assign new_n2114 = new_n2112 & new_n2113;
  assign new_n2115 = new_n2111 & new_n2114;
  assign new_n2116 = new_n2108 & new_n2115;
  assign new_n2117 = new_n2101 & new_n2116;
  assign new_n2118 = ~pdata_5_ & ~new_n2117;
  assign new_n2119 = ~new_n522 & new_n2118;
  assign new_n2120 = pdata_5_ & new_n2117;
  assign new_n2121 = ~new_n522 & new_n2120;
  assign new_n2122 = pinreg_8_ & new_n522;
  assign new_n2123 = ~new_n2119 & ~new_n2121;
  assign pdata_new_37_ = new_n2122 | ~new_n2123;
  assign new_n2125 = ~pcount_0_ & pinreg_3_;
  assign new_n2126 = ~new_n522 & new_n2125;
  assign new_n2127 = pcount_0_ & pdata_in_3_;
  assign new_n2128 = ~new_n522 & new_n2127;
  assign pinreg_new_3_ = new_n2126 | new_n2128;
  assign new_n2130 = pcount_0_ & pinreg_4_;
  assign new_n2131 = ~new_n522 & new_n2130;
  assign new_n2132 = ~pcount_0_ & pinreg_12_;
  assign new_n2133 = ~new_n522 & new_n2132;
  assign pinreg_new_12_ = new_n2131 | new_n2133;
  assign new_n2135 = new_n522 & new_n2120;
  assign new_n2136 = pcount_0_ & poutreg_25_;
  assign new_n2137 = ~new_n522 & new_n2136;
  assign new_n2138 = new_n522 & new_n2118;
  assign new_n2139 = ~pcount_0_ & poutreg_17_;
  assign new_n2140 = ~new_n522 & new_n2139;
  assign new_n2141 = ~new_n2135 & ~new_n2137;
  assign new_n2142 = ~new_n2138 & ~new_n2140;
  assign poutreg_new_17_ = ~new_n2141 | ~new_n2142;
  assign new_n2144 = pc_13_ & new_n535;
  assign new_n2145 = pencrypt_mode_0_ & new_n2144;
  assign new_n2146 = ~new_n529 & new_n2145;
  assign new_n2147 = ~preset_0_ & new_n2146;
  assign new_n2148 = ~pencrypt_mode_0_ & new_n790;
  assign new_n2149 = ~new_n529 & new_n2148;
  assign new_n2150 = ~preset_0_ & new_n2149;
  assign new_n2151 = pc_12_ & new_n530;
  assign new_n2152 = pencrypt_mode_0_ & new_n2151;
  assign new_n2153 = ~new_n529 & new_n2152;
  assign new_n2154 = ~preset_0_ & new_n2153;
  assign new_n2155 = pc_10_ & new_n530;
  assign new_n2156 = ~pencrypt_mode_0_ & new_n2155;
  assign new_n2157 = ~new_n529 & new_n2156;
  assign new_n2158 = ~preset_0_ & new_n2157;
  assign new_n2159 = ~preset_0_ & pc_11_;
  assign new_n2160 = ~new_n512 & new_n2159;
  assign new_n2161 = ~new_n529 & new_n2160;
  assign new_n2162 = pinreg_17_ & new_n582;
  assign new_n2163 = new_n529 & new_n2162;
  assign new_n2164 = pinreg_25_ & new_n554;
  assign new_n2165 = new_n529 & new_n2164;
  assign new_n2166 = ~new_n2161 & ~new_n2163;
  assign new_n2167 = ~new_n2165 & new_n2166;
  assign new_n2168 = ~new_n2147 & ~new_n2150;
  assign new_n2169 = ~new_n2154 & ~new_n2158;
  assign new_n2170 = new_n2168 & new_n2169;
  assign pc_new_11_ = ~new_n2167 | ~new_n2170;
  assign new_n2172 = pc_21_ & new_n530;
  assign new_n2173 = ~pencrypt_mode_0_ & new_n2172;
  assign new_n2174 = ~new_n529 & new_n2173;
  assign new_n2175 = ~preset_0_ & new_n2174;
  assign new_n2176 = pc_24_ & new_n535;
  assign new_n2177 = pencrypt_mode_0_ & new_n2176;
  assign new_n2178 = ~new_n529 & new_n2177;
  assign new_n2179 = ~preset_0_ & new_n2178;
  assign new_n2180 = ~preset_0_ & pc_22_;
  assign new_n2181 = ~new_n512 & new_n2180;
  assign new_n2182 = ~new_n529 & new_n2181;
  assign new_n2183 = pc_23_ & new_n530;
  assign new_n2184 = pencrypt_mode_0_ & new_n2183;
  assign new_n2185 = ~new_n529 & new_n2184;
  assign new_n2186 = ~preset_0_ & new_n2185;
  assign new_n2187 = ~preset_0_ & pdata_in_2_;
  assign new_n2188 = pencrypt_0_ & new_n2187;
  assign new_n2189 = new_n529 & new_n2188;
  assign new_n2190 = pc_20_ & new_n535;
  assign new_n2191 = ~pencrypt_mode_0_ & new_n2190;
  assign new_n2192 = ~new_n529 & new_n2191;
  assign new_n2193 = ~preset_0_ & new_n2192;
  assign new_n2194 = pinreg_2_ & new_n554;
  assign new_n2195 = new_n529 & new_n2194;
  assign new_n2196 = ~new_n2189 & ~new_n2193;
  assign new_n2197 = ~new_n2195 & new_n2196;
  assign new_n2198 = ~new_n2175 & ~new_n2179;
  assign new_n2199 = ~new_n2182 & ~new_n2186;
  assign new_n2200 = new_n2198 & new_n2199;
  assign pc_new_22_ = ~new_n2197 | ~new_n2200;
  assign new_n2202 = pd_14_ & new_n535;
  assign new_n2203 = pencrypt_mode_0_ & new_n2202;
  assign new_n2204 = ~new_n529 & new_n2203;
  assign new_n2205 = ~preset_0_ & new_n2204;
  assign new_n2206 = pd_10_ & new_n535;
  assign new_n2207 = ~pencrypt_mode_0_ & new_n2206;
  assign new_n2208 = ~new_n529 & new_n2207;
  assign new_n2209 = ~preset_0_ & new_n2208;
  assign new_n2210 = pd_13_ & new_n530;
  assign new_n2211 = pencrypt_mode_0_ & new_n2210;
  assign new_n2212 = ~new_n529 & new_n2211;
  assign new_n2213 = ~preset_0_ & new_n2212;
  assign new_n2214 = pd_11_ & new_n530;
  assign new_n2215 = ~pencrypt_mode_0_ & new_n2214;
  assign new_n2216 = ~new_n529 & new_n2215;
  assign new_n2217 = ~preset_0_ & new_n2216;
  assign new_n2218 = ~preset_0_ & pd_12_;
  assign new_n2219 = ~new_n512 & new_n2218;
  assign new_n2220 = ~new_n529 & new_n2219;
  assign new_n2221 = pinreg_13_ & new_n582;
  assign new_n2222 = new_n529 & new_n2221;
  assign new_n2223 = pinreg_21_ & new_n554;
  assign new_n2224 = new_n529 & new_n2223;
  assign new_n2225 = ~new_n2220 & ~new_n2222;
  assign new_n2226 = ~new_n2224 & new_n2225;
  assign new_n2227 = ~new_n2205 & ~new_n2209;
  assign new_n2228 = ~new_n2213 & ~new_n2217;
  assign new_n2229 = new_n2227 & new_n2228;
  assign pd_new_12_ = ~new_n2226 | ~new_n2229;
  assign new_n2231 = pd_22_ & new_n530;
  assign new_n2232 = ~pencrypt_mode_0_ & new_n2231;
  assign new_n2233 = ~new_n529 & new_n2232;
  assign new_n2234 = ~preset_0_ & new_n2233;
  assign new_n2235 = pd_25_ & new_n535;
  assign new_n2236 = pencrypt_mode_0_ & new_n2235;
  assign new_n2237 = ~new_n529 & new_n2236;
  assign new_n2238 = ~preset_0_ & new_n2237;
  assign new_n2239 = ~preset_0_ & pd_23_;
  assign new_n2240 = ~new_n512 & new_n2239;
  assign new_n2241 = ~new_n529 & new_n2240;
  assign new_n2242 = pd_24_ & new_n530;
  assign new_n2243 = pencrypt_mode_0_ & new_n2242;
  assign new_n2244 = ~new_n529 & new_n2243;
  assign new_n2245 = ~preset_0_ & new_n2244;
  assign new_n2246 = ~preset_0_ & pdata_in_4_;
  assign new_n2247 = ~pencrypt_0_ & new_n2246;
  assign new_n2248 = new_n529 & new_n2247;
  assign new_n2249 = ~pencrypt_mode_0_ & new_n845;
  assign new_n2250 = ~new_n529 & new_n2249;
  assign new_n2251 = ~preset_0_ & new_n2250;
  assign new_n2252 = pinreg_19_ & new_n582;
  assign new_n2253 = new_n529 & new_n2252;
  assign new_n2254 = ~new_n2248 & ~new_n2251;
  assign new_n2255 = ~new_n2253 & new_n2254;
  assign new_n2256 = ~new_n2234 & ~new_n2238;
  assign new_n2257 = ~new_n2241 & ~new_n2245;
  assign new_n2258 = new_n2256 & new_n2257;
  assign pd_new_23_ = ~new_n2255 | ~new_n2258;
  assign new_n2260 = ~pcount_0_ & ~preset_0_;
  assign pcount_new_0_ = ~new_n529 & new_n2260;
  assign new_n2262 = pinreg_25_ & new_n522;
  assign new_n2263 = pdata_35_ & ~new_n522;
  assign pdata_new_3_ = new_n2262 | new_n2263;
  assign new_n2265 = ~new_n522 & new_n1088;
  assign new_n2266 = ~new_n522 & new_n1084;
  assign new_n2267 = pinreg_10_ & new_n522;
  assign new_n2268 = ~new_n2265 & ~new_n2266;
  assign pdata_new_45_ = new_n2267 | ~new_n2268;
  assign new_n2270 = new_n1379 & new_n1455;
  assign new_n2271 = new_n1382 & new_n2270;
  assign new_n2272 = new_n1382 & new_n1460;
  assign new_n2273 = ~new_n1379 & new_n1435;
  assign new_n2274 = ~new_n1382 & new_n2273;
  assign new_n2275 = ~new_n1379 & new_n1431;
  assign new_n2276 = ~new_n1382 & new_n2275;
  assign new_n2277 = new_n1382 & new_n1438;
  assign new_n2278 = ~new_n1382 & new_n1446;
  assign new_n2279 = new_n1379 & new_n1428;
  assign new_n2280 = ~new_n1382 & new_n2279;
  assign new_n2281 = new_n1379 & new_n1414;
  assign new_n2282 = ~new_n1382 & new_n2281;
  assign new_n2283 = ~new_n1379 & new_n1422;
  assign new_n2284 = ~new_n1382 & new_n2283;
  assign new_n2285 = ~new_n1379 & new_n1403;
  assign new_n2286 = new_n1382 & new_n2285;
  assign new_n2287 = new_n1382 & new_n1423;
  assign new_n2288 = new_n1382 & new_n1452;
  assign new_n2289 = new_n1382 & new_n2273;
  assign new_n2290 = ~new_n1382 & new_n1391;
  assign new_n2291 = ~new_n1382 & new_n1400;
  assign new_n2292 = new_n1379 & new_n1408;
  assign new_n2293 = new_n1382 & new_n2292;
  assign new_n2294 = ~new_n1466 & ~new_n2293;
  assign new_n2295 = new_n1468 & new_n2294;
  assign new_n2296 = ~new_n2290 & ~new_n2291;
  assign new_n2297 = ~new_n1454 & ~new_n2289;
  assign new_n2298 = new_n2296 & new_n2297;
  assign new_n2299 = new_n2295 & new_n2298;
  assign new_n2300 = ~new_n1453 & ~new_n2288;
  assign new_n2301 = ~new_n1412 & ~new_n2287;
  assign new_n2302 = new_n2300 & new_n2301;
  assign new_n2303 = ~new_n1444 & ~new_n2286;
  assign new_n2304 = ~new_n1433 & ~new_n1439;
  assign new_n2305 = new_n2303 & new_n2304;
  assign new_n2306 = new_n2302 & new_n2305;
  assign new_n2307 = new_n2299 & new_n2306;
  assign new_n2308 = ~new_n2282 & ~new_n2284;
  assign new_n2309 = ~new_n1430 & ~new_n1457;
  assign new_n2310 = new_n2308 & new_n2309;
  assign new_n2311 = ~new_n1427 & ~new_n2280;
  assign new_n2312 = ~new_n2277 & ~new_n2278;
  assign new_n2313 = new_n2311 & new_n2312;
  assign new_n2314 = new_n2310 & new_n2313;
  assign new_n2315 = ~new_n1465 & ~new_n2271;
  assign new_n2316 = ~new_n1396 & ~new_n2272;
  assign new_n2317 = new_n2315 & new_n2316;
  assign new_n2318 = ~new_n1405 & ~new_n2274;
  assign new_n2319 = ~new_n1418 & ~new_n2276;
  assign new_n2320 = new_n2318 & new_n2319;
  assign new_n2321 = new_n2317 & new_n2320;
  assign new_n2322 = new_n2314 & new_n2321;
  assign new_n2323 = new_n2307 & new_n2322;
  assign new_n2324 = ~pdata_26_ & ~new_n2323;
  assign new_n2325 = ~new_n522 & new_n2324;
  assign new_n2326 = pdata_26_ & new_n2323;
  assign new_n2327 = ~new_n522 & new_n2326;
  assign new_n2328 = pinreg_38_ & new_n522;
  assign new_n2329 = ~new_n2325 & ~new_n2327;
  assign pdata_new_58_ = new_n2328 | ~new_n2329;
  assign new_n2331 = ~pcount_0_ & pinreg_22_;
  assign new_n2332 = ~new_n522 & new_n2331;
  assign new_n2333 = pcount_0_ & pinreg_14_;
  assign new_n2334 = ~new_n522 & new_n2333;
  assign pinreg_new_22_ = new_n2332 | new_n2334;
  assign new_n2336 = ~pcount_0_ & pinreg_33_;
  assign new_n2337 = ~new_n522 & new_n2336;
  assign new_n2338 = pcount_0_ & pinreg_25_;
  assign new_n2339 = ~new_n522 & new_n2338;
  assign pinreg_new_33_ = new_n2337 | new_n2339;
  assign new_n2341 = ~pcount_0_ & pinreg_44_;
  assign new_n2342 = ~new_n522 & new_n2341;
  assign new_n2343 = pcount_0_ & pinreg_36_;
  assign new_n2344 = ~new_n522 & new_n2343;
  assign pinreg_new_44_ = new_n2342 | new_n2344;
  assign new_n2346 = ~pcount_0_ & pinreg_55_;
  assign new_n2347 = ~new_n522 & new_n2346;
  assign new_n2348 = pcount_0_ & pinreg_47_;
  assign new_n2349 = ~new_n522 & new_n2348;
  assign pinreg_new_55_ = new_n2347 | new_n2349;
  assign new_n2351 = new_n522 & new_n1016;
  assign new_n2352 = pcount_0_ & poutreg_9_;
  assign new_n2353 = ~new_n522 & new_n2352;
  assign new_n2354 = new_n522 & new_n1014;
  assign new_n2355 = ~pcount_0_ & poutreg_1_;
  assign new_n2356 = ~new_n522 & new_n2355;
  assign new_n2357 = ~new_n2351 & ~new_n2353;
  assign new_n2358 = ~new_n2354 & ~new_n2356;
  assign poutreg_new_1_ = ~new_n2357 | ~new_n2358;
  assign new_n2360 = new_n522 & new_n1500;
  assign new_n2361 = pcount_0_ & poutreg_33_;
  assign new_n2362 = ~new_n522 & new_n2361;
  assign new_n2363 = new_n522 & new_n1498;
  assign new_n2364 = ~pcount_0_ & poutreg_25_;
  assign new_n2365 = ~new_n522 & new_n2364;
  assign new_n2366 = ~new_n2360 & ~new_n2362;
  assign new_n2367 = ~new_n2363 & ~new_n2365;
  assign poutreg_new_25_ = ~new_n2366 | ~new_n2367;
  assign new_n2369 = ~pcount_0_ & poutreg_38_;
  assign new_n2370 = ~new_n522 & new_n2369;
  assign new_n2371 = pcount_0_ & poutreg_46_;
  assign new_n2372 = ~new_n522 & new_n2371;
  assign new_n2373 = pdata_59_ & new_n522;
  assign new_n2374 = ~new_n2370 & ~new_n2372;
  assign poutreg_new_38_ = new_n2373 | ~new_n2374;
  assign new_n2376 = new_n1744 & new_n1797;
  assign new_n2377 = new_n1747 & new_n2376;
  assign new_n2378 = new_n1747 & new_n1831;
  assign new_n2379 = new_n1744 & new_n1787;
  assign new_n2380 = new_n1747 & new_n2379;
  assign new_n2381 = ~new_n1747 & new_n1782;
  assign new_n2382 = new_n1747 & new_n1803;
  assign new_n2383 = ~new_n1747 & new_n1825;
  assign new_n2384 = ~new_n1747 & new_n1816;
  assign new_n2385 = ~new_n1744 & new_n1755;
  assign new_n2386 = new_n1747 & new_n2385;
  assign new_n2387 = ~new_n1747 & new_n1813;
  assign new_n2388 = new_n1747 & new_n1795;
  assign new_n2389 = new_n1747 & new_n1751;
  assign new_n2390 = new_n1747 & new_n1788;
  assign new_n2391 = ~new_n1747 & new_n1818;
  assign new_n2392 = ~new_n1747 & new_n2376;
  assign new_n2393 = new_n1744 & new_n1802;
  assign new_n2394 = ~new_n1747 & new_n2393;
  assign new_n2395 = new_n1744 & new_n1824;
  assign new_n2396 = ~new_n1747 & new_n2395;
  assign new_n2397 = ~new_n1830 & ~new_n2396;
  assign new_n2398 = new_n1855 & new_n2397;
  assign new_n2399 = ~new_n1829 & ~new_n2394;
  assign new_n2400 = ~new_n1789 & ~new_n2392;
  assign new_n2401 = new_n2399 & new_n2400;
  assign new_n2402 = new_n2398 & new_n2401;
  assign new_n2403 = ~new_n2390 & ~new_n2391;
  assign new_n2404 = ~new_n2388 & ~new_n2389;
  assign new_n2405 = new_n2403 & new_n2404;
  assign new_n2406 = ~new_n1826 & ~new_n2387;
  assign new_n2407 = ~new_n1811 & ~new_n2386;
  assign new_n2408 = new_n2406 & new_n2407;
  assign new_n2409 = new_n2405 & new_n2408;
  assign new_n2410 = new_n2402 & new_n2409;
  assign new_n2411 = ~new_n1823 & ~new_n1827;
  assign new_n2412 = ~new_n1783 & ~new_n1820;
  assign new_n2413 = new_n2411 & new_n2412;
  assign new_n2414 = ~new_n1814 & ~new_n2384;
  assign new_n2415 = ~new_n2382 & ~new_n2383;
  assign new_n2416 = new_n2414 & new_n2415;
  assign new_n2417 = new_n2413 & new_n2416;
  assign new_n2418 = ~new_n1766 & ~new_n1771;
  assign new_n2419 = ~new_n2377 & ~new_n2378;
  assign new_n2420 = new_n2418 & new_n2419;
  assign new_n2421 = ~new_n1808 & ~new_n2380;
  assign new_n2422 = ~new_n1806 & ~new_n2381;
  assign new_n2423 = new_n2421 & new_n2422;
  assign new_n2424 = new_n2420 & new_n2423;
  assign new_n2425 = new_n2417 & new_n2424;
  assign new_n2426 = new_n2410 & new_n2425;
  assign new_n2427 = ~pdata_16_ & ~new_n2426;
  assign new_n2428 = new_n522 & new_n2427;
  assign new_n2429 = pdata_16_ & new_n2426;
  assign new_n2430 = new_n522 & new_n2429;
  assign new_n2431 = ~pcount_0_ & poutreg_61_;
  assign new_n2432 = ~new_n522 & new_n2431;
  assign new_n2433 = ~new_n2428 & ~new_n2430;
  assign poutreg_new_61_ = new_n2432 | ~new_n2433;
  assign new_n2435 = pc_14_ & new_n535;
  assign new_n2436 = pencrypt_mode_0_ & new_n2435;
  assign new_n2437 = ~new_n529 & new_n2436;
  assign new_n2438 = ~preset_0_ & new_n2437;
  assign new_n2439 = pc_10_ & new_n535;
  assign new_n2440 = ~pencrypt_mode_0_ & new_n2439;
  assign new_n2441 = ~new_n529 & new_n2440;
  assign new_n2442 = ~preset_0_ & new_n2441;
  assign new_n2443 = pc_13_ & new_n530;
  assign new_n2444 = pencrypt_mode_0_ & new_n2443;
  assign new_n2445 = ~new_n529 & new_n2444;
  assign new_n2446 = ~preset_0_ & new_n2445;
  assign new_n2447 = pc_11_ & new_n530;
  assign new_n2448 = ~pencrypt_mode_0_ & new_n2447;
  assign new_n2449 = ~new_n529 & new_n2448;
  assign new_n2450 = ~preset_0_ & new_n2449;
  assign new_n2451 = ~preset_0_ & pc_12_;
  assign new_n2452 = ~new_n512 & new_n2451;
  assign new_n2453 = ~new_n529 & new_n2452;
  assign new_n2454 = pinreg_17_ & new_n554;
  assign new_n2455 = new_n529 & new_n2454;
  assign new_n2456 = pinreg_9_ & new_n582;
  assign new_n2457 = new_n529 & new_n2456;
  assign new_n2458 = ~new_n2453 & ~new_n2455;
  assign new_n2459 = ~new_n2457 & new_n2458;
  assign new_n2460 = ~new_n2438 & ~new_n2442;
  assign new_n2461 = ~new_n2446 & ~new_n2450;
  assign new_n2462 = new_n2460 & new_n2461;
  assign pc_new_12_ = ~new_n2459 | ~new_n2462;
  assign new_n2464 = pc_23_ & new_n535;
  assign new_n2465 = pencrypt_mode_0_ & new_n2464;
  assign new_n2466 = ~new_n529 & new_n2465;
  assign new_n2467 = ~preset_0_ & new_n2466;
  assign new_n2468 = pc_19_ & new_n535;
  assign new_n2469 = ~pencrypt_mode_0_ & new_n2468;
  assign new_n2470 = ~new_n529 & new_n2469;
  assign new_n2471 = ~preset_0_ & new_n2470;
  assign new_n2472 = pc_22_ & new_n530;
  assign new_n2473 = pencrypt_mode_0_ & new_n2472;
  assign new_n2474 = ~new_n529 & new_n2473;
  assign new_n2475 = ~preset_0_ & new_n2474;
  assign new_n2476 = ~pencrypt_mode_0_ & new_n571;
  assign new_n2477 = ~new_n529 & new_n2476;
  assign new_n2478 = ~preset_0_ & new_n2477;
  assign new_n2479 = ~preset_0_ & pc_21_;
  assign new_n2480 = ~new_n512 & new_n2479;
  assign new_n2481 = ~new_n529 & new_n2480;
  assign new_n2482 = pinreg_10_ & new_n554;
  assign new_n2483 = new_n529 & new_n2482;
  assign new_n2484 = pinreg_2_ & new_n582;
  assign new_n2485 = new_n529 & new_n2484;
  assign new_n2486 = ~new_n2481 & ~new_n2483;
  assign new_n2487 = ~new_n2485 & new_n2486;
  assign new_n2488 = ~new_n2467 & ~new_n2471;
  assign new_n2489 = ~new_n2475 & ~new_n2478;
  assign new_n2490 = new_n2488 & new_n2489;
  assign pc_new_21_ = ~new_n2487 | ~new_n2490;
  assign new_n2492 = pd_13_ & new_n535;
  assign new_n2493 = pencrypt_mode_0_ & new_n2492;
  assign new_n2494 = ~new_n529 & new_n2493;
  assign new_n2495 = ~preset_0_ & new_n2494;
  assign new_n2496 = pd_9_ & new_n535;
  assign new_n2497 = ~pencrypt_mode_0_ & new_n2496;
  assign new_n2498 = ~new_n529 & new_n2497;
  assign new_n2499 = ~preset_0_ & new_n2498;
  assign new_n2500 = pd_12_ & new_n530;
  assign new_n2501 = pencrypt_mode_0_ & new_n2500;
  assign new_n2502 = ~new_n529 & new_n2501;
  assign new_n2503 = ~preset_0_ & new_n2502;
  assign new_n2504 = pd_10_ & new_n530;
  assign new_n2505 = ~pencrypt_mode_0_ & new_n2504;
  assign new_n2506 = ~new_n529 & new_n2505;
  assign new_n2507 = ~preset_0_ & new_n2506;
  assign new_n2508 = ~preset_0_ & pd_11_;
  assign new_n2509 = ~new_n512 & new_n2508;
  assign new_n2510 = ~new_n529 & new_n2509;
  assign new_n2511 = pinreg_21_ & new_n582;
  assign new_n2512 = new_n529 & new_n2511;
  assign new_n2513 = pinreg_29_ & new_n554;
  assign new_n2514 = new_n529 & new_n2513;
  assign new_n2515 = ~new_n2510 & ~new_n2512;
  assign new_n2516 = ~new_n2514 & new_n2515;
  assign new_n2517 = ~new_n2495 & ~new_n2499;
  assign new_n2518 = ~new_n2503 & ~new_n2507;
  assign new_n2519 = new_n2517 & new_n2518;
  assign pd_new_11_ = ~new_n2516 | ~new_n2519;
  assign new_n2521 = pencrypt_mode_0_ & new_n1957;
  assign new_n2522 = ~new_n529 & new_n2521;
  assign new_n2523 = ~preset_0_ & new_n2522;
  assign new_n2524 = pd_22_ & new_n535;
  assign new_n2525 = ~pencrypt_mode_0_ & new_n2524;
  assign new_n2526 = ~new_n529 & new_n2525;
  assign new_n2527 = ~preset_0_ & new_n2526;
  assign new_n2528 = pd_25_ & new_n530;
  assign new_n2529 = pencrypt_mode_0_ & new_n2528;
  assign new_n2530 = ~new_n529 & new_n2529;
  assign new_n2531 = ~preset_0_ & new_n2530;
  assign new_n2532 = pd_23_ & new_n530;
  assign new_n2533 = ~pencrypt_mode_0_ & new_n2532;
  assign new_n2534 = ~new_n529 & new_n2533;
  assign new_n2535 = ~preset_0_ & new_n2534;
  assign new_n2536 = ~preset_0_ & pd_24_;
  assign new_n2537 = ~new_n512 & new_n2536;
  assign new_n2538 = ~new_n529 & new_n2537;
  assign new_n2539 = pinreg_11_ & new_n582;
  assign new_n2540 = new_n529 & new_n2539;
  assign new_n2541 = pinreg_19_ & new_n554;
  assign new_n2542 = new_n529 & new_n2541;
  assign new_n2543 = ~new_n2538 & ~new_n2540;
  assign new_n2544 = ~new_n2542 & new_n2543;
  assign new_n2545 = ~new_n2523 & ~new_n2527;
  assign new_n2546 = ~new_n2531 & ~new_n2535;
  assign new_n2547 = new_n2545 & new_n2546;
  assign pd_new_24_ = ~new_n2544 | ~new_n2547;
  assign new_n2549 = pinreg_17_ & new_n522;
  assign new_n2550 = pdata_36_ & ~new_n522;
  assign pdata_new_4_ = new_n2549 | new_n2550;
  assign new_n2552 = new_n1382 & new_n2281;
  assign new_n2553 = ~new_n1382 & new_n2285;
  assign new_n2554 = ~new_n1382 & new_n2292;
  assign new_n2555 = ~new_n1382 & new_n1456;
  assign new_n2556 = new_n1382 & new_n1429;
  assign new_n2557 = new_n1382 & new_n1462;
  assign new_n2558 = new_n1382 & new_n2275;
  assign new_n2559 = ~new_n1382 & new_n1395;
  assign new_n2560 = ~new_n1465 & ~new_n2293;
  assign new_n2561 = ~new_n1461 & ~new_n1463;
  assign new_n2562 = new_n2560 & new_n2561;
  assign new_n2563 = ~new_n2282 & ~new_n2559;
  assign new_n2564 = ~new_n2291 & ~new_n2558;
  assign new_n2565 = new_n2563 & new_n2564;
  assign new_n2566 = new_n2562 & new_n2565;
  assign new_n2567 = ~new_n1453 & ~new_n2557;
  assign new_n2568 = ~new_n1442 & ~new_n2556;
  assign new_n2569 = new_n2567 & new_n2568;
  assign new_n2570 = ~new_n1433 & ~new_n2555;
  assign new_n2571 = new_n2303 & new_n2570;
  assign new_n2572 = new_n2569 & new_n2571;
  assign new_n2573 = new_n2566 & new_n2572;
  assign new_n2574 = ~new_n1459 & ~new_n2284;
  assign new_n2575 = ~new_n1434 & ~new_n1457;
  assign new_n2576 = new_n2574 & new_n2575;
  assign new_n2577 = ~new_n1420 & ~new_n2554;
  assign new_n2578 = ~new_n2277 & ~new_n2553;
  assign new_n2579 = new_n2577 & new_n2578;
  assign new_n2580 = new_n2576 & new_n2579;
  assign new_n2581 = ~new_n1387 & ~new_n2552;
  assign new_n2582 = new_n1490 & new_n2581;
  assign new_n2583 = ~new_n1410 & ~new_n2272;
  assign new_n2584 = ~new_n1418 & ~new_n2274;
  assign new_n2585 = new_n2583 & new_n2584;
  assign new_n2586 = new_n2582 & new_n2585;
  assign new_n2587 = new_n2580 & new_n2586;
  assign new_n2588 = new_n2573 & new_n2587;
  assign new_n2589 = ~pdata_14_ & ~new_n2588;
  assign new_n2590 = ~new_n522 & new_n2589;
  assign new_n2591 = pdata_14_ & new_n2588;
  assign new_n2592 = ~new_n522 & new_n2591;
  assign new_n2593 = pinreg_2_ & new_n522;
  assign new_n2594 = ~new_n2590 & ~new_n2592;
  assign pdata_new_46_ = new_n2593 | ~new_n2594;
  assign new_n2596 = ~pdata_46_ & pc_19_;
  assign new_n2597 = pdata_46_ & ~pc_19_;
  assign new_n2598 = ~new_n2596 & ~new_n2597;
  assign new_n2599 = ~pdata_47_ & pc_12_;
  assign new_n2600 = pdata_47_ & ~pc_12_;
  assign new_n2601 = ~new_n2599 & ~new_n2600;
  assign new_n2602 = ~pdata_44_ & pc_6_;
  assign new_n2603 = pdata_44_ & ~pc_6_;
  assign new_n2604 = ~new_n2602 & ~new_n2603;
  assign new_n2605 = ~pdata_45_ & pc_26_;
  assign new_n2606 = pdata_45_ & ~pc_26_;
  assign new_n2607 = ~new_n2605 & ~new_n2606;
  assign new_n2608 = ~pdata_43_ & pc_15_;
  assign new_n2609 = pdata_43_ & ~pc_15_;
  assign new_n2610 = ~new_n2608 & ~new_n2609;
  assign new_n2611 = ~pdata_48_ & pc_1_;
  assign new_n2612 = pdata_48_ & ~pc_1_;
  assign new_n2613 = ~new_n2611 & ~new_n2612;
  assign new_n2614 = ~new_n2598 & ~new_n2601;
  assign new_n2615 = new_n2604 & new_n2614;
  assign new_n2616 = ~new_n2607 & new_n2615;
  assign new_n2617 = new_n2610 & new_n2616;
  assign new_n2618 = new_n2613 & new_n2617;
  assign new_n2619 = new_n2598 & new_n2601;
  assign new_n2620 = ~new_n2604 & new_n2619;
  assign new_n2621 = ~new_n2607 & new_n2620;
  assign new_n2622 = new_n2610 & new_n2621;
  assign new_n2623 = new_n2613 & new_n2622;
  assign new_n2624 = ~new_n2598 & new_n2601;
  assign new_n2625 = new_n2604 & new_n2624;
  assign new_n2626 = new_n2607 & new_n2625;
  assign new_n2627 = new_n2610 & new_n2626;
  assign new_n2628 = new_n2613 & new_n2627;
  assign new_n2629 = ~new_n2607 & new_n2625;
  assign new_n2630 = new_n2610 & new_n2629;
  assign new_n2631 = new_n2613 & new_n2630;
  assign new_n2632 = new_n2598 & ~new_n2601;
  assign new_n2633 = new_n2604 & new_n2632;
  assign new_n2634 = new_n2607 & new_n2633;
  assign new_n2635 = new_n2610 & new_n2634;
  assign new_n2636 = new_n2613 & new_n2635;
  assign new_n2637 = ~new_n2604 & new_n2614;
  assign new_n2638 = ~new_n2607 & new_n2637;
  assign new_n2639 = ~new_n2610 & new_n2638;
  assign new_n2640 = ~new_n2613 & new_n2639;
  assign new_n2641 = new_n2604 & new_n2619;
  assign new_n2642 = ~new_n2607 & new_n2641;
  assign new_n2643 = ~new_n2610 & new_n2642;
  assign new_n2644 = new_n2613 & new_n2643;
  assign new_n2645 = ~new_n2610 & new_n2621;
  assign new_n2646 = ~new_n2613 & new_n2645;
  assign new_n2647 = ~new_n2607 & new_n2633;
  assign new_n2648 = ~new_n2610 & new_n2647;
  assign new_n2649 = new_n2613 & new_n2648;
  assign new_n2650 = ~new_n2613 & new_n2635;
  assign new_n2651 = ~new_n2610 & new_n2616;
  assign new_n2652 = new_n2613 & new_n2651;
  assign new_n2653 = ~new_n2613 & new_n2651;
  assign new_n2654 = new_n2607 & new_n2620;
  assign new_n2655 = ~new_n2610 & new_n2654;
  assign new_n2656 = new_n2613 & new_n2655;
  assign new_n2657 = ~new_n2610 & new_n2629;
  assign new_n2658 = ~new_n2613 & new_n2657;
  assign new_n2659 = ~new_n2604 & new_n2624;
  assign new_n2660 = ~new_n2607 & new_n2659;
  assign new_n2661 = new_n2610 & new_n2660;
  assign new_n2662 = ~new_n2613 & new_n2661;
  assign new_n2663 = ~new_n2613 & new_n2643;
  assign new_n2664 = new_n2610 & new_n2638;
  assign new_n2665 = ~new_n2613 & new_n2664;
  assign new_n2666 = new_n2607 & new_n2637;
  assign new_n2667 = ~new_n2610 & new_n2666;
  assign new_n2668 = ~new_n2613 & new_n2667;
  assign new_n2669 = new_n2607 & new_n2641;
  assign new_n2670 = ~new_n2610 & new_n2669;
  assign new_n2671 = new_n2613 & new_n2670;
  assign new_n2672 = ~new_n2613 & new_n2655;
  assign new_n2673 = ~new_n2610 & new_n2626;
  assign new_n2674 = new_n2613 & new_n2673;
  assign new_n2675 = ~new_n2610 & new_n2660;
  assign new_n2676 = new_n2613 & new_n2675;
  assign new_n2677 = new_n2607 & new_n2659;
  assign new_n2678 = new_n2610 & new_n2677;
  assign new_n2679 = new_n2613 & new_n2678;
  assign new_n2680 = ~new_n2610 & new_n2634;
  assign new_n2681 = ~new_n2613 & new_n2680;
  assign new_n2682 = new_n2610 & new_n2666;
  assign new_n2683 = ~new_n2613 & new_n2682;
  assign new_n2684 = new_n2613 & new_n2667;
  assign new_n2685 = ~new_n2604 & new_n2632;
  assign new_n2686 = ~new_n2607 & new_n2685;
  assign new_n2687 = new_n2610 & new_n2686;
  assign new_n2688 = ~new_n2613 & new_n2687;
  assign new_n2689 = new_n2610 & new_n2647;
  assign new_n2690 = ~new_n2613 & new_n2689;
  assign new_n2691 = new_n2610 & new_n2669;
  assign new_n2692 = ~new_n2613 & new_n2691;
  assign new_n2693 = ~new_n2613 & new_n2627;
  assign new_n2694 = new_n2613 & new_n2687;
  assign new_n2695 = new_n2613 & new_n2664;
  assign new_n2696 = ~new_n2694 & ~new_n2695;
  assign new_n2697 = ~new_n2692 & ~new_n2693;
  assign new_n2698 = new_n2696 & new_n2697;
  assign new_n2699 = ~new_n2688 & ~new_n2690;
  assign new_n2700 = ~new_n2683 & ~new_n2684;
  assign new_n2701 = new_n2699 & new_n2700;
  assign new_n2702 = new_n2698 & new_n2701;
  assign new_n2703 = ~new_n2679 & ~new_n2681;
  assign new_n2704 = ~new_n2674 & ~new_n2676;
  assign new_n2705 = new_n2703 & new_n2704;
  assign new_n2706 = ~new_n2671 & ~new_n2672;
  assign new_n2707 = ~new_n2665 & ~new_n2668;
  assign new_n2708 = new_n2706 & new_n2707;
  assign new_n2709 = new_n2705 & new_n2708;
  assign new_n2710 = new_n2702 & new_n2709;
  assign new_n2711 = ~new_n2662 & ~new_n2663;
  assign new_n2712 = ~new_n2656 & ~new_n2658;
  assign new_n2713 = new_n2711 & new_n2712;
  assign new_n2714 = ~new_n2652 & ~new_n2653;
  assign new_n2715 = ~new_n2649 & ~new_n2650;
  assign new_n2716 = new_n2714 & new_n2715;
  assign new_n2717 = new_n2713 & new_n2716;
  assign new_n2718 = ~new_n2618 & ~new_n2623;
  assign new_n2719 = ~new_n2628 & ~new_n2631;
  assign new_n2720 = new_n2718 & new_n2719;
  assign new_n2721 = ~new_n2636 & ~new_n2640;
  assign new_n2722 = ~new_n2644 & ~new_n2646;
  assign new_n2723 = new_n2721 & new_n2722;
  assign new_n2724 = new_n2720 & new_n2723;
  assign new_n2725 = new_n2717 & new_n2724;
  assign new_n2726 = new_n2710 & new_n2725;
  assign new_n2727 = ~pdata_25_ & ~new_n2726;
  assign new_n2728 = ~new_n522 & new_n2727;
  assign new_n2729 = pdata_25_ & new_n2726;
  assign new_n2730 = ~new_n522 & new_n2729;
  assign new_n2731 = pinreg_46_ & new_n522;
  assign new_n2732 = ~new_n2728 & ~new_n2730;
  assign pdata_new_57_ = new_n2731 | ~new_n2732;
  assign new_n2734 = ~pcount_0_ & pinreg_23_;
  assign new_n2735 = ~new_n522 & new_n2734;
  assign new_n2736 = pcount_0_ & pinreg_15_;
  assign new_n2737 = ~new_n522 & new_n2736;
  assign pinreg_new_23_ = new_n2735 | new_n2737;
  assign new_n2739 = ~pcount_0_ & pinreg_32_;
  assign new_n2740 = ~new_n522 & new_n2739;
  assign new_n2741 = pcount_0_ & pinreg_24_;
  assign new_n2742 = ~new_n522 & new_n2741;
  assign pinreg_new_32_ = new_n2740 | new_n2742;
  assign new_n2744 = ~pcount_0_ & pinreg_45_;
  assign new_n2745 = ~new_n522 & new_n2744;
  assign new_n2746 = pcount_0_ & pinreg_37_;
  assign new_n2747 = ~new_n522 & new_n2746;
  assign pinreg_new_45_ = new_n2745 | new_n2747;
  assign new_n2749 = ~pcount_0_ & pinreg_54_;
  assign new_n2750 = ~new_n522 & new_n2749;
  assign new_n2751 = pcount_0_ & pinreg_46_;
  assign new_n2752 = ~new_n522 & new_n2751;
  assign pinreg_new_54_ = new_n2750 | new_n2752;
  assign new_n2754 = pcount_0_ & poutreg_10_;
  assign new_n2755 = ~new_n522 & new_n2754;
  assign new_n2756 = ~pcount_0_ & poutreg_2_;
  assign new_n2757 = ~new_n522 & new_n2756;
  assign new_n2758 = pdata_47_ & new_n522;
  assign new_n2759 = ~new_n2755 & ~new_n2757;
  assign poutreg_new_2_ = new_n2758 | ~new_n2759;
  assign new_n2761 = ~pcount_0_ & poutreg_26_;
  assign new_n2762 = ~new_n522 & new_n2761;
  assign new_n2763 = pcount_0_ & poutreg_34_;
  assign new_n2764 = ~new_n522 & new_n2763;
  assign new_n2765 = pdata_44_ & new_n522;
  assign new_n2766 = ~new_n2762 & ~new_n2764;
  assign poutreg_new_26_ = new_n2765 | ~new_n2766;
  assign new_n2768 = new_n2613 & new_n2689;
  assign new_n2769 = new_n2613 & new_n2682;
  assign new_n2770 = new_n2613 & new_n2691;
  assign new_n2771 = new_n2613 & new_n2657;
  assign new_n2772 = ~new_n2610 & new_n2686;
  assign new_n2773 = ~new_n2613 & new_n2772;
  assign new_n2774 = new_n2610 & new_n2654;
  assign new_n2775 = ~new_n2613 & new_n2774;
  assign new_n2776 = new_n2607 & new_n2685;
  assign new_n2777 = ~new_n2610 & new_n2776;
  assign new_n2778 = ~new_n2613 & new_n2777;
  assign new_n2779 = new_n2607 & new_n2615;
  assign new_n2780 = ~new_n2610 & new_n2779;
  assign new_n2781 = ~new_n2613 & new_n2780;
  assign new_n2782 = new_n2613 & new_n2680;
  assign new_n2783 = ~new_n2610 & new_n2677;
  assign new_n2784 = ~new_n2613 & new_n2783;
  assign new_n2785 = new_n2613 & new_n2639;
  assign new_n2786 = new_n2613 & new_n2661;
  assign new_n2787 = new_n2613 & new_n2645;
  assign new_n2788 = new_n2610 & new_n2776;
  assign new_n2789 = ~new_n2613 & new_n2788;
  assign new_n2790 = new_n2610 & new_n2642;
  assign new_n2791 = ~new_n2613 & new_n2790;
  assign new_n2792 = new_n2610 & new_n2779;
  assign new_n2793 = ~new_n2613 & new_n2792;
  assign new_n2794 = ~new_n2692 & ~new_n2793;
  assign new_n2795 = new_n2696 & new_n2794;
  assign new_n2796 = ~new_n2789 & ~new_n2791;
  assign new_n2797 = ~new_n2690 & ~new_n2787;
  assign new_n2798 = new_n2796 & new_n2797;
  assign new_n2799 = new_n2795 & new_n2798;
  assign new_n2800 = ~new_n2681 & ~new_n2786;
  assign new_n2801 = ~new_n2644 & ~new_n2785;
  assign new_n2802 = new_n2800 & new_n2801;
  assign new_n2803 = ~new_n2782 & ~new_n2784;
  assign new_n2804 = ~new_n2646 & ~new_n2662;
  assign new_n2805 = new_n2803 & new_n2804;
  assign new_n2806 = new_n2802 & new_n2805;
  assign new_n2807 = new_n2799 & new_n2806;
  assign new_n2808 = ~new_n2683 & ~new_n2781;
  assign new_n2809 = ~new_n2658 & ~new_n2684;
  assign new_n2810 = new_n2808 & new_n2809;
  assign new_n2811 = ~new_n2656 & ~new_n2778;
  assign new_n2812 = ~new_n2652 & ~new_n2775;
  assign new_n2813 = new_n2811 & new_n2812;
  assign new_n2814 = new_n2810 & new_n2813;
  assign new_n2815 = ~new_n2768 & ~new_n2769;
  assign new_n2816 = ~new_n2628 & ~new_n2636;
  assign new_n2817 = new_n2815 & new_n2816;
  assign new_n2818 = ~new_n2640 & ~new_n2770;
  assign new_n2819 = ~new_n2771 & ~new_n2773;
  assign new_n2820 = new_n2818 & new_n2819;
  assign new_n2821 = new_n2817 & new_n2820;
  assign new_n2822 = new_n2814 & new_n2821;
  assign new_n2823 = new_n2807 & new_n2822;
  assign new_n2824 = pdata_19_ & new_n2823;
  assign new_n2825 = new_n522 & new_n2824;
  assign new_n2826 = pcount_0_ & poutreg_45_;
  assign new_n2827 = ~new_n522 & new_n2826;
  assign new_n2828 = ~pdata_19_ & ~new_n2823;
  assign new_n2829 = new_n522 & new_n2828;
  assign new_n2830 = ~pcount_0_ & poutreg_37_;
  assign new_n2831 = ~new_n522 & new_n2830;
  assign new_n2832 = ~new_n2825 & ~new_n2827;
  assign new_n2833 = ~new_n2829 & ~new_n2831;
  assign poutreg_new_37_ = ~new_n2832 | ~new_n2833;
  assign new_n2835 = poutreg_62_ & ~pcount_0_;
  assign new_n2836 = ~new_n522 & new_n2835;
  assign new_n2837 = pdata_56_ & new_n522;
  assign poutreg_new_62_ = new_n2836 | new_n2837;
  assign new_n2839 = pc_15_ & new_n535;
  assign new_n2840 = pencrypt_mode_0_ & new_n2839;
  assign new_n2841 = ~new_n529 & new_n2840;
  assign new_n2842 = ~preset_0_ & new_n2841;
  assign new_n2843 = pc_11_ & new_n535;
  assign new_n2844 = ~pencrypt_mode_0_ & new_n2843;
  assign new_n2845 = ~new_n529 & new_n2844;
  assign new_n2846 = ~preset_0_ & new_n2845;
  assign new_n2847 = pc_14_ & new_n530;
  assign new_n2848 = pencrypt_mode_0_ & new_n2847;
  assign new_n2849 = ~new_n529 & new_n2848;
  assign new_n2850 = ~preset_0_ & new_n2849;
  assign new_n2851 = ~pencrypt_mode_0_ & new_n2151;
  assign new_n2852 = ~new_n529 & new_n2851;
  assign new_n2853 = ~preset_0_ & new_n2852;
  assign new_n2854 = ~preset_0_ & pc_13_;
  assign new_n2855 = ~new_n512 & new_n2854;
  assign new_n2856 = ~new_n529 & new_n2855;
  assign new_n2857 = pinreg_1_ & new_n582;
  assign new_n2858 = new_n529 & new_n2857;
  assign new_n2859 = pinreg_9_ & new_n554;
  assign new_n2860 = new_n529 & new_n2859;
  assign new_n2861 = ~new_n2856 & ~new_n2858;
  assign new_n2862 = ~new_n2860 & new_n2861;
  assign new_n2863 = ~new_n2842 & ~new_n2846;
  assign new_n2864 = ~new_n2850 & ~new_n2853;
  assign new_n2865 = new_n2863 & new_n2864;
  assign pc_new_13_ = ~new_n2862 | ~new_n2865;
  assign new_n2867 = pencrypt_mode_0_ & new_n1878;
  assign new_n2868 = ~new_n529 & new_n2867;
  assign new_n2869 = ~preset_0_ & new_n2868;
  assign new_n2870 = pc_22_ & new_n535;
  assign new_n2871 = ~pencrypt_mode_0_ & new_n2870;
  assign new_n2872 = ~new_n529 & new_n2871;
  assign new_n2873 = ~preset_0_ & new_n2872;
  assign new_n2874 = pc_25_ & new_n530;
  assign new_n2875 = pencrypt_mode_0_ & new_n2874;
  assign new_n2876 = ~new_n529 & new_n2875;
  assign new_n2877 = ~preset_0_ & new_n2876;
  assign new_n2878 = ~pencrypt_mode_0_ & new_n2183;
  assign new_n2879 = ~new_n529 & new_n2878;
  assign new_n2880 = ~preset_0_ & new_n2879;
  assign new_n2881 = ~preset_0_ & pc_24_;
  assign new_n2882 = ~new_n512 & new_n2881;
  assign new_n2883 = ~new_n529 & new_n2882;
  assign new_n2884 = pinreg_43_ & new_n582;
  assign new_n2885 = new_n529 & new_n2884;
  assign new_n2886 = pinreg_51_ & new_n554;
  assign new_n2887 = new_n529 & new_n2886;
  assign new_n2888 = ~new_n2883 & ~new_n2885;
  assign new_n2889 = ~new_n2887 & new_n2888;
  assign new_n2890 = ~new_n2869 & ~new_n2873;
  assign new_n2891 = ~new_n2877 & ~new_n2880;
  assign new_n2892 = new_n2890 & new_n2891;
  assign pc_new_24_ = ~new_n2889 | ~new_n2892;
  assign new_n2894 = ~pencrypt_mode_0_ & new_n2210;
  assign new_n2895 = ~new_n529 & new_n2894;
  assign new_n2896 = ~preset_0_ & new_n2895;
  assign new_n2897 = pd_16_ & new_n535;
  assign new_n2898 = pencrypt_mode_0_ & new_n2897;
  assign new_n2899 = ~new_n529 & new_n2898;
  assign new_n2900 = ~preset_0_ & new_n2899;
  assign new_n2901 = ~preset_0_ & pd_14_;
  assign new_n2902 = ~new_n512 & new_n2901;
  assign new_n2903 = ~new_n529 & new_n2902;
  assign new_n2904 = pd_15_ & new_n530;
  assign new_n2905 = pencrypt_mode_0_ & new_n2904;
  assign new_n2906 = ~new_n529 & new_n2905;
  assign new_n2907 = ~preset_0_ & new_n2906;
  assign new_n2908 = ~preset_0_ & pdata_in_5_;
  assign new_n2909 = pencrypt_0_ & new_n2908;
  assign new_n2910 = new_n529 & new_n2909;
  assign new_n2911 = pd_12_ & new_n535;
  assign new_n2912 = ~pencrypt_mode_0_ & new_n2911;
  assign new_n2913 = ~new_n529 & new_n2912;
  assign new_n2914 = ~preset_0_ & new_n2913;
  assign new_n2915 = pinreg_5_ & new_n554;
  assign new_n2916 = new_n529 & new_n2915;
  assign new_n2917 = ~new_n2910 & ~new_n2914;
  assign new_n2918 = ~new_n2916 & new_n2917;
  assign new_n2919 = ~new_n2896 & ~new_n2900;
  assign new_n2920 = ~new_n2903 & ~new_n2907;
  assign new_n2921 = new_n2919 & new_n2920;
  assign pd_new_14_ = ~new_n2918 | ~new_n2921;
  assign new_n2923 = pd_23_ & new_n535;
  assign new_n2924 = pencrypt_mode_0_ & new_n2923;
  assign new_n2925 = ~new_n529 & new_n2924;
  assign new_n2926 = ~preset_0_ & new_n2925;
  assign new_n2927 = pd_19_ & new_n535;
  assign new_n2928 = ~pencrypt_mode_0_ & new_n2927;
  assign new_n2929 = ~new_n529 & new_n2928;
  assign new_n2930 = ~preset_0_ & new_n2929;
  assign new_n2931 = pencrypt_mode_0_ & new_n2231;
  assign new_n2932 = ~new_n529 & new_n2931;
  assign new_n2933 = ~preset_0_ & new_n2932;
  assign new_n2934 = ~pencrypt_mode_0_ & new_n853;
  assign new_n2935 = ~new_n529 & new_n2934;
  assign new_n2936 = ~preset_0_ & new_n2935;
  assign new_n2937 = ~preset_0_ & pd_21_;
  assign new_n2938 = ~new_n512 & new_n2937;
  assign new_n2939 = ~new_n529 & new_n2938;
  assign new_n2940 = pinreg_12_ & new_n554;
  assign new_n2941 = new_n529 & new_n2940;
  assign new_n2942 = pinreg_4_ & new_n582;
  assign new_n2943 = new_n529 & new_n2942;
  assign new_n2944 = ~new_n2939 & ~new_n2941;
  assign new_n2945 = ~new_n2943 & new_n2944;
  assign new_n2946 = ~new_n2926 & ~new_n2930;
  assign new_n2947 = ~new_n2933 & ~new_n2936;
  assign new_n2948 = new_n2946 & new_n2947;
  assign pd_new_21_ = ~new_n2945 | ~new_n2948;
  assign new_n2950 = ~pcount_1_ & ~preset_0_;
  assign new_n2951 = pcount_2_ & new_n2950;
  assign new_n2952 = ~new_n529 & new_n2951;
  assign new_n2953 = pcount_1_ & pcount_0_;
  assign new_n2954 = ~preset_0_ & new_n2953;
  assign new_n2955 = ~pcount_2_ & new_n2954;
  assign new_n2956 = ~new_n529 & new_n2955;
  assign new_n2957 = pcount_2_ & new_n2260;
  assign new_n2958 = ~new_n529 & new_n2957;
  assign new_n2959 = ~new_n2952 & ~new_n2956;
  assign pcount_new_2_ = new_n2958 | ~new_n2959;
  assign new_n2961 = pinreg_41_ & new_n522;
  assign new_n2962 = pdata_33_ & ~new_n522;
  assign pdata_new_1_ = new_n2961 | new_n2962;
  assign new_n2964 = new_n1998 & new_n2069;
  assign new_n2965 = new_n1998 & new_n2076;
  assign new_n2966 = ~new_n1998 & new_n2071;
  assign new_n2967 = new_n1998 & new_n2055;
  assign new_n2968 = ~new_n1998 & new_n2038;
  assign new_n2969 = ~new_n1998 & new_n2011;
  assign new_n2970 = ~new_n1995 & new_n2051;
  assign new_n2971 = new_n1998 & new_n2970;
  assign new_n2972 = ~new_n1998 & new_n2085;
  assign new_n2973 = ~new_n1995 & new_n2068;
  assign new_n2974 = ~new_n1998 & new_n2973;
  assign new_n2975 = ~new_n1995 & new_n2073;
  assign new_n2976 = ~new_n1998 & new_n2975;
  assign new_n2977 = ~new_n1995 & new_n2080;
  assign new_n2978 = new_n1998 & new_n2977;
  assign new_n2979 = new_n1998 & new_n2047;
  assign new_n2980 = new_n1998 & new_n2066;
  assign new_n2981 = ~new_n1998 & new_n2083;
  assign new_n2982 = ~new_n1998 & new_n2016;
  assign new_n2983 = new_n1998 & new_n2074;
  assign new_n2984 = ~new_n2084 & ~new_n2983;
  assign new_n2985 = new_n2088 & new_n2984;
  assign new_n2986 = ~new_n2981 & ~new_n2982;
  assign new_n2987 = ~new_n2072 & ~new_n2075;
  assign new_n2988 = new_n2986 & new_n2987;
  assign new_n2989 = new_n2985 & new_n2988;
  assign new_n2990 = ~new_n2067 & ~new_n2980;
  assign new_n2991 = ~new_n2978 & ~new_n2979;
  assign new_n2992 = new_n2990 & new_n2991;
  assign new_n2993 = ~new_n2053 & ~new_n2976;
  assign new_n2994 = new_n2097 & new_n2993;
  assign new_n2995 = new_n2992 & new_n2994;
  assign new_n2996 = new_n2989 & new_n2995;
  assign new_n2997 = ~new_n2972 & ~new_n2974;
  assign new_n2998 = ~new_n2046 & ~new_n2971;
  assign new_n2999 = new_n2997 & new_n2998;
  assign new_n3000 = ~new_n2044 & ~new_n2969;
  assign new_n3001 = ~new_n2967 & ~new_n2968;
  assign new_n3002 = new_n3000 & new_n3001;
  assign new_n3003 = new_n2999 & new_n3002;
  assign new_n3004 = ~new_n2017 & ~new_n2964;
  assign new_n3005 = new_n2109 & new_n3004;
  assign new_n3006 = ~new_n2965 & ~new_n2966;
  assign new_n3007 = ~new_n2023 & ~new_n2025;
  assign new_n3008 = new_n3006 & new_n3007;
  assign new_n3009 = new_n3005 & new_n3008;
  assign new_n3010 = new_n3003 & new_n3009;
  assign new_n3011 = new_n2996 & new_n3010;
  assign new_n3012 = ~pdata_15_ & ~new_n3011;
  assign new_n3013 = ~new_n522 & new_n3012;
  assign new_n3014 = pdata_15_ & new_n3011;
  assign new_n3015 = ~new_n522 & new_n3014;
  assign new_n3016 = pdata_in_2_ & new_n522;
  assign new_n3017 = ~new_n3013 & ~new_n3015;
  assign pdata_new_47_ = new_n3016 | ~new_n3017;
  assign new_n3019 = new_n897 & new_n973;
  assign new_n3020 = ~new_n897 & new_n971;
  assign new_n3021 = ~new_n897 & new_n1049;
  assign new_n3022 = ~new_n897 & new_n1047;
  assign new_n3023 = new_n897 & new_n1041;
  assign new_n3024 = ~new_n897 & new_n906;
  assign new_n3025 = new_n897 & new_n938;
  assign new_n3026 = new_n897 & new_n977;
  assign new_n3027 = ~new_n902 & ~new_n980;
  assign new_n3028 = new_n984 & new_n3027;
  assign new_n3029 = ~new_n944 & ~new_n1053;
  assign new_n3030 = ~new_n972 & ~new_n974;
  assign new_n3031 = new_n3029 & new_n3030;
  assign new_n3032 = new_n3028 & new_n3031;
  assign new_n3033 = ~new_n968 & ~new_n3026;
  assign new_n3034 = ~new_n962 & ~new_n3025;
  assign new_n3035 = new_n3033 & new_n3034;
  assign new_n3036 = ~new_n955 & ~new_n1046;
  assign new_n3037 = ~new_n951 & ~new_n1045;
  assign new_n3038 = new_n3036 & new_n3037;
  assign new_n3039 = new_n3035 & new_n3038;
  assign new_n3040 = new_n3032 & new_n3039;
  assign new_n3041 = ~new_n1044 & ~new_n3024;
  assign new_n3042 = ~new_n943 & ~new_n3023;
  assign new_n3043 = new_n3041 & new_n3042;
  assign new_n3044 = ~new_n1043 & ~new_n3022;
  assign new_n3045 = ~new_n929 & ~new_n3021;
  assign new_n3046 = new_n3044 & new_n3045;
  assign new_n3047 = new_n3043 & new_n3046;
  assign new_n3048 = ~new_n1036 & ~new_n3019;
  assign new_n3049 = new_n1006 & new_n3048;
  assign new_n3050 = ~new_n1034 & ~new_n3020;
  assign new_n3051 = ~new_n922 & ~new_n1048;
  assign new_n3052 = new_n3050 & new_n3051;
  assign new_n3053 = new_n3049 & new_n3052;
  assign new_n3054 = new_n3047 & new_n3053;
  assign new_n3055 = new_n3040 & new_n3054;
  assign new_n3056 = ~pdata_24_ & ~new_n3055;
  assign new_n3057 = ~new_n522 & new_n3056;
  assign new_n3058 = pdata_24_ & new_n3055;
  assign new_n3059 = ~new_n522 & new_n3058;
  assign new_n3060 = pinreg_54_ & new_n522;
  assign new_n3061 = ~new_n3057 & ~new_n3059;
  assign pdata_new_56_ = new_n3060 | ~new_n3061;
  assign new_n3063 = pinreg_0_ & ~pcount_0_;
  assign new_n3064 = ~new_n522 & new_n3063;
  assign new_n3065 = pcount_0_ & pdata_in_0_;
  assign new_n3066 = ~new_n522 & new_n3065;
  assign pinreg_new_0_ = new_n3064 | new_n3066;
  assign new_n3068 = ~pcount_0_ & pinreg_24_;
  assign new_n3069 = ~new_n522 & new_n3068;
  assign new_n3070 = pcount_0_ & pinreg_16_;
  assign new_n3071 = ~new_n522 & new_n3070;
  assign pinreg_new_24_ = new_n3069 | new_n3071;
  assign new_n3073 = ~pcount_0_ & pinreg_35_;
  assign new_n3074 = ~new_n522 & new_n3073;
  assign new_n3075 = pcount_0_ & pinreg_27_;
  assign new_n3076 = ~new_n522 & new_n3075;
  assign pinreg_new_35_ = new_n3074 | new_n3076;
  assign new_n3078 = ~pcount_0_ & pinreg_42_;
  assign new_n3079 = ~new_n522 & new_n3078;
  assign new_n3080 = pcount_0_ & pinreg_34_;
  assign new_n3081 = ~new_n522 & new_n3080;
  assign pinreg_new_42_ = new_n3079 | new_n3081;
  assign new_n3083 = ~pcount_0_ & pinreg_53_;
  assign new_n3084 = ~new_n522 & new_n3083;
  assign new_n3085 = pcount_0_ & pinreg_45_;
  assign new_n3086 = ~new_n522 & new_n3085;
  assign pinreg_new_53_ = new_n3084 | new_n3086;
  assign new_n3088 = ~pdata_36_ & pc_27_;
  assign new_n3089 = pdata_36_ & ~pc_27_;
  assign new_n3090 = ~new_n3088 & ~new_n3089;
  assign new_n3091 = ~pdata_37_ & pc_14_;
  assign new_n3092 = pdata_37_ & ~pc_14_;
  assign new_n3093 = ~new_n3091 & ~new_n3092;
  assign new_n3094 = ~pdata_40_ & pc_9_;
  assign new_n3095 = pdata_40_ & ~pc_9_;
  assign new_n3096 = ~new_n3094 & ~new_n3095;
  assign new_n3097 = ~pdata_35_ & pc_2_;
  assign new_n3098 = pdata_35_ & ~pc_2_;
  assign new_n3099 = ~new_n3097 & ~new_n3098;
  assign new_n3100 = pc_20_ & ~pdata_39_;
  assign new_n3101 = ~pc_20_ & pdata_39_;
  assign new_n3102 = ~new_n3100 & ~new_n3101;
  assign new_n3103 = ~pdata_38_ & pc_5_;
  assign new_n3104 = pdata_38_ & ~pc_5_;
  assign new_n3105 = ~new_n3103 & ~new_n3104;
  assign new_n3106 = ~new_n3090 & new_n3093;
  assign new_n3107 = new_n3096 & new_n3106;
  assign new_n3108 = ~new_n3099 & new_n3107;
  assign new_n3109 = new_n3102 & new_n3108;
  assign new_n3110 = ~new_n3105 & new_n3109;
  assign new_n3111 = ~new_n3090 & ~new_n3093;
  assign new_n3112 = new_n3096 & new_n3111;
  assign new_n3113 = ~new_n3099 & new_n3112;
  assign new_n3114 = new_n3102 & new_n3113;
  assign new_n3115 = new_n3105 & new_n3114;
  assign new_n3116 = new_n3090 & ~new_n3093;
  assign new_n3117 = new_n3096 & new_n3116;
  assign new_n3118 = ~new_n3099 & new_n3117;
  assign new_n3119 = new_n3102 & new_n3118;
  assign new_n3120 = new_n3105 & new_n3119;
  assign new_n3121 = ~new_n3105 & new_n3119;
  assign new_n3122 = new_n3090 & new_n3093;
  assign new_n3123 = new_n3096 & new_n3122;
  assign new_n3124 = ~new_n3099 & new_n3123;
  assign new_n3125 = ~new_n3102 & new_n3124;
  assign new_n3126 = ~new_n3105 & new_n3125;
  assign new_n3127 = new_n3105 & new_n3125;
  assign new_n3128 = new_n3099 & new_n3107;
  assign new_n3129 = new_n3102 & new_n3128;
  assign new_n3130 = new_n3105 & new_n3129;
  assign new_n3131 = ~new_n3096 & new_n3111;
  assign new_n3132 = new_n3099 & new_n3131;
  assign new_n3133 = new_n3102 & new_n3132;
  assign new_n3134 = ~new_n3105 & new_n3133;
  assign new_n3135 = ~new_n3102 & new_n3128;
  assign new_n3136 = ~new_n3105 & new_n3135;
  assign new_n3137 = new_n3099 & new_n3123;
  assign new_n3138 = new_n3102 & new_n3137;
  assign new_n3139 = ~new_n3105 & new_n3138;
  assign new_n3140 = new_n3099 & new_n3112;
  assign new_n3141 = new_n3102 & new_n3140;
  assign new_n3142 = new_n3105 & new_n3141;
  assign new_n3143 = ~new_n3096 & new_n3116;
  assign new_n3144 = new_n3099 & new_n3143;
  assign new_n3145 = new_n3102 & new_n3144;
  assign new_n3146 = ~new_n3105 & new_n3145;
  assign new_n3147 = ~new_n3102 & new_n3140;
  assign new_n3148 = ~new_n3105 & new_n3147;
  assign new_n3149 = ~new_n3096 & new_n3106;
  assign new_n3150 = new_n3099 & new_n3149;
  assign new_n3151 = new_n3102 & new_n3150;
  assign new_n3152 = new_n3105 & new_n3151;
  assign new_n3153 = ~new_n3099 & new_n3131;
  assign new_n3154 = ~new_n3102 & new_n3153;
  assign new_n3155 = ~new_n3105 & new_n3154;
  assign new_n3156 = ~new_n3102 & new_n3144;
  assign new_n3157 = ~new_n3105 & new_n3156;
  assign new_n3158 = new_n3105 & new_n3138;
  assign new_n3159 = ~new_n3102 & new_n3132;
  assign new_n3160 = new_n3105 & new_n3159;
  assign new_n3161 = ~new_n3102 & new_n3137;
  assign new_n3162 = ~new_n3105 & new_n3161;
  assign new_n3163 = ~new_n3102 & new_n3150;
  assign new_n3164 = ~new_n3105 & new_n3163;
  assign new_n3165 = new_n3099 & new_n3117;
  assign new_n3166 = ~new_n3102 & new_n3165;
  assign new_n3167 = new_n3105 & new_n3166;
  assign new_n3168 = ~new_n3102 & new_n3108;
  assign new_n3169 = new_n3105 & new_n3168;
  assign new_n3170 = ~new_n3096 & new_n3122;
  assign new_n3171 = ~new_n3099 & new_n3170;
  assign new_n3172 = ~new_n3102 & new_n3171;
  assign new_n3173 = new_n3105 & new_n3172;
  assign new_n3174 = new_n3105 & new_n3145;
  assign new_n3175 = ~new_n3099 & new_n3149;
  assign new_n3176 = ~new_n3102 & new_n3175;
  assign new_n3177 = ~new_n3105 & new_n3176;
  assign new_n3178 = new_n3099 & new_n3170;
  assign new_n3179 = ~new_n3102 & new_n3178;
  assign new_n3180 = new_n3105 & new_n3179;
  assign new_n3181 = new_n3102 & new_n3153;
  assign new_n3182 = ~new_n3105 & new_n3181;
  assign new_n3183 = new_n3102 & new_n3175;
  assign new_n3184 = new_n3105 & new_n3183;
  assign new_n3185 = new_n3102 & new_n3171;
  assign new_n3186 = ~new_n3105 & new_n3185;
  assign new_n3187 = ~new_n3099 & new_n3143;
  assign new_n3188 = ~new_n3102 & new_n3187;
  assign new_n3189 = new_n3105 & new_n3188;
  assign new_n3190 = ~new_n3102 & new_n3113;
  assign new_n3191 = ~new_n3105 & new_n3190;
  assign new_n3192 = new_n3105 & new_n3185;
  assign new_n3193 = ~new_n3191 & ~new_n3192;
  assign new_n3194 = ~new_n3186 & ~new_n3189;
  assign new_n3195 = new_n3193 & new_n3194;
  assign new_n3196 = ~new_n3182 & ~new_n3184;
  assign new_n3197 = ~new_n3177 & ~new_n3180;
  assign new_n3198 = new_n3196 & new_n3197;
  assign new_n3199 = new_n3195 & new_n3198;
  assign new_n3200 = ~new_n3173 & ~new_n3174;
  assign new_n3201 = ~new_n3167 & ~new_n3169;
  assign new_n3202 = new_n3200 & new_n3201;
  assign new_n3203 = ~new_n3162 & ~new_n3164;
  assign new_n3204 = ~new_n3158 & ~new_n3160;
  assign new_n3205 = new_n3203 & new_n3204;
  assign new_n3206 = new_n3202 & new_n3205;
  assign new_n3207 = new_n3199 & new_n3206;
  assign new_n3208 = ~new_n3155 & ~new_n3157;
  assign new_n3209 = ~new_n3148 & ~new_n3152;
  assign new_n3210 = new_n3208 & new_n3209;
  assign new_n3211 = ~new_n3142 & ~new_n3146;
  assign new_n3212 = ~new_n3136 & ~new_n3139;
  assign new_n3213 = new_n3211 & new_n3212;
  assign new_n3214 = new_n3210 & new_n3213;
  assign new_n3215 = ~new_n3110 & ~new_n3115;
  assign new_n3216 = ~new_n3120 & ~new_n3121;
  assign new_n3217 = new_n3215 & new_n3216;
  assign new_n3218 = ~new_n3126 & ~new_n3127;
  assign new_n3219 = ~new_n3130 & ~new_n3134;
  assign new_n3220 = new_n3218 & new_n3219;
  assign new_n3221 = new_n3217 & new_n3220;
  assign new_n3222 = new_n3214 & new_n3221;
  assign new_n3223 = new_n3207 & new_n3222;
  assign new_n3224 = pdata_12_ & new_n3223;
  assign new_n3225 = new_n522 & new_n3224;
  assign new_n3226 = pcount_0_ & poutreg_35_;
  assign new_n3227 = ~new_n522 & new_n3226;
  assign new_n3228 = ~pdata_12_ & ~new_n3223;
  assign new_n3229 = new_n522 & new_n3228;
  assign new_n3230 = ~pcount_0_ & poutreg_27_;
  assign new_n3231 = ~new_n522 & new_n3230;
  assign new_n3232 = ~new_n3225 & ~new_n3227;
  assign new_n3233 = ~new_n3229 & ~new_n3231;
  assign poutreg_new_27_ = ~new_n3232 | ~new_n3233;
  assign new_n3235 = ~pcount_0_ & poutreg_36_;
  assign new_n3236 = ~new_n522 & new_n3235;
  assign new_n3237 = pcount_0_ & poutreg_44_;
  assign new_n3238 = ~new_n522 & new_n3237;
  assign new_n3239 = pdata_51_ & new_n522;
  assign new_n3240 = ~new_n3236 & ~new_n3238;
  assign poutreg_new_36_ = new_n3239 | ~new_n3240;
  assign new_n3242 = new_n3105 & new_n3190;
  assign new_n3243 = ~new_n3105 & new_n3168;
  assign new_n3244 = new_n3102 & new_n3124;
  assign new_n3245 = ~new_n3105 & new_n3244;
  assign new_n3246 = new_n3102 & new_n3165;
  assign new_n3247 = ~new_n3105 & new_n3246;
  assign new_n3248 = new_n3105 & new_n3135;
  assign new_n3249 = ~new_n3105 & new_n3188;
  assign new_n3250 = ~new_n3105 & new_n3114;
  assign new_n3251 = new_n3102 & new_n3178;
  assign new_n3252 = new_n3105 & new_n3251;
  assign new_n3253 = new_n3105 & new_n3246;
  assign new_n3254 = new_n3105 & new_n3133;
  assign new_n3255 = ~new_n3105 & new_n3129;
  assign new_n3256 = new_n3105 & new_n3156;
  assign new_n3257 = ~new_n3105 & new_n3183;
  assign new_n3258 = ~new_n3105 & new_n3179;
  assign new_n3259 = new_n3105 & new_n3176;
  assign new_n3260 = new_n3102 & new_n3187;
  assign new_n3261 = new_n3105 & new_n3260;
  assign new_n3262 = ~new_n3186 & ~new_n3261;
  assign new_n3263 = ~new_n3184 & ~new_n3189;
  assign new_n3264 = new_n3262 & new_n3263;
  assign new_n3265 = ~new_n3182 & ~new_n3259;
  assign new_n3266 = ~new_n3257 & ~new_n3258;
  assign new_n3267 = new_n3265 & new_n3266;
  assign new_n3268 = new_n3264 & new_n3267;
  assign new_n3269 = ~new_n3174 & ~new_n3256;
  assign new_n3270 = ~new_n3167 & ~new_n3255;
  assign new_n3271 = new_n3269 & new_n3270;
  assign new_n3272 = ~new_n3253 & ~new_n3254;
  assign new_n3273 = ~new_n3134 & ~new_n3162;
  assign new_n3274 = new_n3272 & new_n3273;
  assign new_n3275 = new_n3271 & new_n3274;
  assign new_n3276 = new_n3268 & new_n3275;
  assign new_n3277 = ~new_n3157 & ~new_n3158;
  assign new_n3278 = ~new_n3164 & ~new_n3252;
  assign new_n3279 = new_n3277 & new_n3278;
  assign new_n3280 = ~new_n3148 & ~new_n3250;
  assign new_n3281 = ~new_n3248 & ~new_n3249;
  assign new_n3282 = new_n3280 & new_n3281;
  assign new_n3283 = new_n3279 & new_n3282;
  assign new_n3284 = ~new_n3191 & ~new_n3242;
  assign new_n3285 = ~new_n3120 & ~new_n3243;
  assign new_n3286 = new_n3284 & new_n3285;
  assign new_n3287 = ~new_n3126 & ~new_n3245;
  assign new_n3288 = ~new_n3127 & ~new_n3247;
  assign new_n3289 = new_n3287 & new_n3288;
  assign new_n3290 = new_n3286 & new_n3289;
  assign new_n3291 = new_n3283 & new_n3290;
  assign new_n3292 = new_n3276 & new_n3291;
  assign new_n3293 = pdata_1_ & new_n3292;
  assign new_n3294 = new_n522 & new_n3293;
  assign new_n3295 = pcount_0_ & poutreg_57_;
  assign new_n3296 = ~new_n522 & new_n3295;
  assign new_n3297 = ~pdata_1_ & ~new_n3292;
  assign new_n3298 = new_n522 & new_n3297;
  assign new_n3299 = ~pcount_0_ & poutreg_49_;
  assign new_n3300 = ~new_n522 & new_n3299;
  assign new_n3301 = ~new_n3294 & ~new_n3296;
  assign new_n3302 = ~new_n3298 & ~new_n3300;
  assign poutreg_new_49_ = ~new_n3301 | ~new_n3302;
  assign new_n3304 = ~pcount_0_ & poutreg_50_;
  assign new_n3305 = ~new_n522 & new_n3304;
  assign new_n3306 = pcount_0_ & poutreg_58_;
  assign new_n3307 = ~new_n522 & new_n3306;
  assign new_n3308 = pdata_41_ & new_n522;
  assign new_n3309 = ~new_n3305 & ~new_n3307;
  assign poutreg_new_50_ = new_n3308 | ~new_n3309;
  assign new_n3311 = new_n522 & new_n3056;
  assign new_n3312 = new_n522 & new_n3058;
  assign new_n3313 = poutreg_63_ & ~pcount_0_;
  assign new_n3314 = ~new_n522 & new_n3313;
  assign new_n3315 = ~new_n3311 & ~new_n3312;
  assign poutreg_new_63_ = new_n3314 | ~new_n3315;
  assign new_n3317 = ~pencrypt_mode_0_ & new_n2443;
  assign new_n3318 = ~new_n529 & new_n3317;
  assign new_n3319 = ~preset_0_ & new_n3318;
  assign new_n3320 = pc_16_ & new_n535;
  assign new_n3321 = pencrypt_mode_0_ & new_n3320;
  assign new_n3322 = ~new_n529 & new_n3321;
  assign new_n3323 = ~preset_0_ & new_n3322;
  assign new_n3324 = ~preset_0_ & pc_14_;
  assign new_n3325 = ~new_n512 & new_n3324;
  assign new_n3326 = ~new_n529 & new_n3325;
  assign new_n3327 = pc_15_ & new_n530;
  assign new_n3328 = pencrypt_mode_0_ & new_n3327;
  assign new_n3329 = ~new_n529 & new_n3328;
  assign new_n3330 = ~preset_0_ & new_n3329;
  assign new_n3331 = ~preset_0_ & pdata_in_1_;
  assign new_n3332 = pencrypt_0_ & new_n3331;
  assign new_n3333 = new_n529 & new_n3332;
  assign new_n3334 = pc_12_ & new_n535;
  assign new_n3335 = ~pencrypt_mode_0_ & new_n3334;
  assign new_n3336 = ~new_n529 & new_n3335;
  assign new_n3337 = ~preset_0_ & new_n3336;
  assign new_n3338 = pinreg_1_ & new_n554;
  assign new_n3339 = new_n529 & new_n3338;
  assign new_n3340 = ~new_n3333 & ~new_n3337;
  assign new_n3341 = ~new_n3339 & new_n3340;
  assign new_n3342 = ~new_n3319 & ~new_n3323;
  assign new_n3343 = ~new_n3326 & ~new_n3330;
  assign new_n3344 = new_n3342 & new_n3343;
  assign pc_new_14_ = ~new_n3341 | ~new_n3344;
  assign new_n3346 = ~pencrypt_mode_0_ & new_n2472;
  assign new_n3347 = ~new_n529 & new_n3346;
  assign new_n3348 = ~preset_0_ & new_n3347;
  assign new_n3349 = pc_25_ & new_n535;
  assign new_n3350 = pencrypt_mode_0_ & new_n3349;
  assign new_n3351 = ~new_n529 & new_n3350;
  assign new_n3352 = ~preset_0_ & new_n3351;
  assign new_n3353 = ~preset_0_ & pc_23_;
  assign new_n3354 = ~new_n512 & new_n3353;
  assign new_n3355 = ~new_n529 & new_n3354;
  assign new_n3356 = pc_24_ & new_n530;
  assign new_n3357 = pencrypt_mode_0_ & new_n3356;
  assign new_n3358 = ~new_n529 & new_n3357;
  assign new_n3359 = ~preset_0_ & new_n3358;
  assign new_n3360 = ~pencrypt_0_ & new_n2187;
  assign new_n3361 = new_n529 & new_n3360;
  assign new_n3362 = ~pencrypt_mode_0_ & new_n563;
  assign new_n3363 = ~new_n529 & new_n3362;
  assign new_n3364 = ~preset_0_ & new_n3363;
  assign new_n3365 = pinreg_51_ & new_n582;
  assign new_n3366 = new_n529 & new_n3365;
  assign new_n3367 = ~new_n3361 & ~new_n3364;
  assign new_n3368 = ~new_n3366 & new_n3367;
  assign new_n3369 = ~new_n3348 & ~new_n3352;
  assign new_n3370 = ~new_n3355 & ~new_n3359;
  assign new_n3371 = new_n3369 & new_n3370;
  assign pc_new_23_ = ~new_n3368 | ~new_n3371;
  assign new_n3373 = pd_15_ & new_n535;
  assign new_n3374 = pencrypt_mode_0_ & new_n3373;
  assign new_n3375 = ~new_n529 & new_n3374;
  assign new_n3376 = ~preset_0_ & new_n3375;
  assign new_n3377 = pd_11_ & new_n535;
  assign new_n3378 = ~pencrypt_mode_0_ & new_n3377;
  assign new_n3379 = ~new_n529 & new_n3378;
  assign new_n3380 = ~preset_0_ & new_n3379;
  assign new_n3381 = pd_14_ & new_n530;
  assign new_n3382 = pencrypt_mode_0_ & new_n3381;
  assign new_n3383 = ~new_n529 & new_n3382;
  assign new_n3384 = ~preset_0_ & new_n3383;
  assign new_n3385 = ~pencrypt_mode_0_ & new_n2500;
  assign new_n3386 = ~new_n529 & new_n3385;
  assign new_n3387 = ~preset_0_ & new_n3386;
  assign new_n3388 = ~preset_0_ & pd_13_;
  assign new_n3389 = ~new_n512 & new_n3388;
  assign new_n3390 = ~new_n529 & new_n3389;
  assign new_n3391 = pinreg_13_ & new_n554;
  assign new_n3392 = new_n529 & new_n3391;
  assign new_n3393 = pinreg_5_ & new_n582;
  assign new_n3394 = new_n529 & new_n3393;
  assign new_n3395 = ~new_n3390 & ~new_n3392;
  assign new_n3396 = ~new_n3394 & new_n3395;
  assign new_n3397 = ~new_n3376 & ~new_n3380;
  assign new_n3398 = ~new_n3384 & ~new_n3387;
  assign new_n3399 = new_n3397 & new_n3398;
  assign pd_new_13_ = ~new_n3396 | ~new_n3399;
  assign new_n3401 = pd_21_ & new_n530;
  assign new_n3402 = ~pencrypt_mode_0_ & new_n3401;
  assign new_n3403 = ~new_n529 & new_n3402;
  assign new_n3404 = ~preset_0_ & new_n3403;
  assign new_n3405 = pd_24_ & new_n535;
  assign new_n3406 = pencrypt_mode_0_ & new_n3405;
  assign new_n3407 = ~new_n529 & new_n3406;
  assign new_n3408 = ~preset_0_ & new_n3407;
  assign new_n3409 = ~preset_0_ & pd_22_;
  assign new_n3410 = ~new_n512 & new_n3409;
  assign new_n3411 = ~new_n529 & new_n3410;
  assign new_n3412 = pencrypt_mode_0_ & new_n2532;
  assign new_n3413 = ~new_n529 & new_n3412;
  assign new_n3414 = ~preset_0_ & new_n3413;
  assign new_n3415 = pencrypt_0_ & new_n2246;
  assign new_n3416 = new_n529 & new_n3415;
  assign new_n3417 = pd_20_ & new_n535;
  assign new_n3418 = ~pencrypt_mode_0_ & new_n3417;
  assign new_n3419 = ~new_n529 & new_n3418;
  assign new_n3420 = ~preset_0_ & new_n3419;
  assign new_n3421 = pinreg_4_ & new_n554;
  assign new_n3422 = new_n529 & new_n3421;
  assign new_n3423 = ~new_n3416 & ~new_n3420;
  assign new_n3424 = ~new_n3422 & new_n3423;
  assign new_n3425 = ~new_n3404 & ~new_n3408;
  assign new_n3426 = ~new_n3411 & ~new_n3414;
  assign new_n3427 = new_n3425 & new_n3426;
  assign pd_new_22_ = ~new_n3424 | ~new_n3427;
  assign new_n3429 = pcount_0_ & new_n2950;
  assign new_n3430 = ~new_n529 & new_n3429;
  assign new_n3431 = pcount_1_ & ~preset_0_;
  assign new_n3432 = ~pcount_0_ & new_n3431;
  assign new_n3433 = ~new_n529 & new_n3432;
  assign pcount_new_1_ = new_n3430 | new_n3433;
  assign new_n3435 = pinreg_33_ & new_n522;
  assign new_n3436 = pdata_34_ & ~new_n522;
  assign pdata_new_2_ = new_n3435 | new_n3436;
  assign new_n3438 = ~new_n522 & new_n2427;
  assign new_n3439 = ~new_n522 & new_n2429;
  assign new_n3440 = pinreg_52_ & new_n522;
  assign new_n3441 = ~new_n3438 & ~new_n3439;
  assign pdata_new_48_ = new_n3440 | ~new_n3441;
  assign new_n3443 = new_n1998 & new_n2078;
  assign new_n3444 = ~new_n1998 & new_n2031;
  assign new_n3445 = ~new_n1998 & new_n2007;
  assign new_n3446 = new_n1998 & new_n2022;
  assign new_n3447 = new_n1998 & new_n2042;
  assign new_n3448 = new_n1998 & new_n2973;
  assign new_n3449 = ~new_n1998 & new_n2977;
  assign new_n3450 = ~new_n1998 & new_n2002;
  assign new_n3451 = ~new_n2086 & ~new_n2983;
  assign new_n3452 = ~new_n2077 & ~new_n2079;
  assign new_n3453 = new_n3451 & new_n3452;
  assign new_n3454 = ~new_n2972 & ~new_n3450;
  assign new_n3455 = ~new_n2971 & ~new_n2981;
  assign new_n3456 = new_n3454 & new_n3455;
  assign new_n3457 = new_n3453 & new_n3456;
  assign new_n3458 = ~new_n3448 & ~new_n3449;
  assign new_n3459 = ~new_n2062 & ~new_n3447;
  assign new_n3460 = new_n3458 & new_n3459;
  assign new_n3461 = new_n2994 & new_n3460;
  assign new_n3462 = new_n3457 & new_n3461;
  assign new_n3463 = ~new_n2048 & ~new_n2067;
  assign new_n3464 = ~new_n2049 & ~new_n3446;
  assign new_n3465 = new_n3463 & new_n3464;
  assign new_n3466 = ~new_n2967 & ~new_n3445;
  assign new_n3467 = ~new_n2039 & ~new_n3444;
  assign new_n3468 = new_n3466 & new_n3467;
  assign new_n3469 = new_n3465 & new_n3468;
  assign new_n3470 = ~new_n2008 & ~new_n2017;
  assign new_n3471 = ~new_n2020 & ~new_n2965;
  assign new_n3472 = new_n3470 & new_n3471;
  assign new_n3473 = ~new_n2966 & ~new_n3443;
  assign new_n3474 = new_n2113 & new_n3473;
  assign new_n3475 = new_n3472 & new_n3474;
  assign new_n3476 = new_n3469 & new_n3475;
  assign new_n3477 = new_n3462 & new_n3476;
  assign new_n3478 = ~pdata_23_ & ~new_n3477;
  assign new_n3479 = ~new_n522 & new_n3478;
  assign new_n3480 = pdata_23_ & new_n3477;
  assign new_n3481 = ~new_n522 & new_n3480;
  assign new_n3482 = pdata_in_4_ & new_n522;
  assign new_n3483 = ~new_n3479 & ~new_n3481;
  assign pdata_new_55_ = new_n3482 | ~new_n3483;
  assign new_n3485 = ~pcount_0_ & pinreg_25_;
  assign new_n3486 = ~new_n522 & new_n3485;
  assign new_n3487 = pcount_0_ & pinreg_17_;
  assign new_n3488 = ~new_n522 & new_n3487;
  assign pinreg_new_25_ = new_n3486 | new_n3488;
  assign new_n3490 = ~pcount_0_ & pinreg_34_;
  assign new_n3491 = ~new_n522 & new_n3490;
  assign new_n3492 = pcount_0_ & pinreg_26_;
  assign new_n3493 = ~new_n522 & new_n3492;
  assign pinreg_new_34_ = new_n3491 | new_n3493;
  assign new_n3495 = ~pcount_0_ & pinreg_43_;
  assign new_n3496 = ~new_n522 & new_n3495;
  assign new_n3497 = pcount_0_ & pinreg_35_;
  assign new_n3498 = ~new_n522 & new_n3497;
  assign pinreg_new_43_ = new_n3496 | new_n3498;
  assign new_n3500 = ~pcount_0_ & pinreg_52_;
  assign new_n3501 = ~new_n522 & new_n3500;
  assign new_n3502 = pcount_0_ & pinreg_44_;
  assign new_n3503 = ~new_n522 & new_n3502;
  assign pinreg_new_52_ = new_n3501 | new_n3503;
  assign new_n3505 = ~pcount_0_ & poutreg_0_;
  assign new_n3506 = ~new_n522 & new_n3505;
  assign new_n3507 = pcount_0_ & poutreg_8_;
  assign new_n3508 = ~new_n522 & new_n3507;
  assign new_n3509 = pdata_39_ & new_n522;
  assign new_n3510 = ~new_n3506 & ~new_n3508;
  assign poutreg_new_0_ = new_n3509 | ~new_n3510;
  assign new_n3512 = ~pcount_0_ & poutreg_28_;
  assign new_n3513 = ~new_n522 & new_n3512;
  assign new_n3514 = pcount_0_ & poutreg_36_;
  assign new_n3515 = ~new_n522 & new_n3514;
  assign new_n3516 = pdata_52_ & new_n522;
  assign new_n3517 = ~new_n3513 & ~new_n3515;
  assign poutreg_new_28_ = new_n3516 | ~new_n3517;
  assign new_n3519 = ~new_n655 & new_n668;
  assign new_n3520 = ~new_n655 & new_n684;
  assign new_n3521 = ~new_n652 & new_n663;
  assign new_n3522 = new_n655 & new_n3521;
  assign new_n3523 = ~new_n655 & new_n721;
  assign new_n3524 = new_n655 & new_n726;
  assign new_n3525 = new_n655 & new_n735;
  assign new_n3526 = ~new_n655 & new_n724;
  assign new_n3527 = new_n655 & new_n1178;
  assign new_n3528 = ~new_n743 & ~new_n3527;
  assign new_n3529 = ~new_n734 & ~new_n736;
  assign new_n3530 = new_n3528 & new_n3529;
  assign new_n3531 = ~new_n1183 & ~new_n1187;
  assign new_n3532 = ~new_n704 & ~new_n707;
  assign new_n3533 = new_n3531 & new_n3532;
  assign new_n3534 = new_n3530 & new_n3533;
  assign new_n3535 = ~new_n3525 & ~new_n3526;
  assign new_n3536 = ~new_n1174 & ~new_n3524;
  assign new_n3537 = new_n3535 & new_n3536;
  assign new_n3538 = ~new_n713 & ~new_n719;
  assign new_n3539 = ~new_n689 & ~new_n3523;
  assign new_n3540 = new_n3538 & new_n3539;
  assign new_n3541 = new_n3537 & new_n3540;
  assign new_n3542 = new_n3534 & new_n3541;
  assign new_n3543 = ~new_n710 & ~new_n712;
  assign new_n3544 = ~new_n706 & ~new_n3522;
  assign new_n3545 = new_n3543 & new_n3544;
  assign new_n3546 = ~new_n699 & ~new_n3520;
  assign new_n3547 = ~new_n1177 & ~new_n3519;
  assign new_n3548 = new_n3546 & new_n3547;
  assign new_n3549 = new_n3545 & new_n3548;
  assign new_n3550 = ~new_n740 & ~new_n1170;
  assign new_n3551 = new_n767 & new_n3550;
  assign new_n3552 = ~new_n1171 & ~new_n1173;
  assign new_n3553 = ~new_n693 & ~new_n1176;
  assign new_n3554 = new_n3552 & new_n3553;
  assign new_n3555 = new_n3551 & new_n3554;
  assign new_n3556 = new_n3549 & new_n3555;
  assign new_n3557 = new_n3542 & new_n3556;
  assign new_n3558 = pdata_11_ & new_n3557;
  assign new_n3559 = new_n522 & new_n3558;
  assign new_n3560 = pcount_0_ & poutreg_43_;
  assign new_n3561 = ~new_n522 & new_n3560;
  assign new_n3562 = ~pdata_11_ & ~new_n3557;
  assign new_n3563 = new_n522 & new_n3562;
  assign new_n3564 = ~pcount_0_ & poutreg_35_;
  assign new_n3565 = ~new_n522 & new_n3564;
  assign new_n3566 = ~new_n3559 & ~new_n3561;
  assign new_n3567 = ~new_n3563 & ~new_n3565;
  assign poutreg_new_35_ = ~new_n3566 | ~new_n3567;
  assign new_n3569 = ~pencrypt_mode_0_ & new_n2847;
  assign new_n3570 = ~new_n529 & new_n3569;
  assign new_n3571 = ~preset_0_ & new_n3570;
  assign new_n3572 = pencrypt_mode_0_ & new_n567;
  assign new_n3573 = ~new_n529 & new_n3572;
  assign new_n3574 = ~preset_0_ & new_n3573;
  assign new_n3575 = ~preset_0_ & pc_15_;
  assign new_n3576 = ~new_n512 & new_n3575;
  assign new_n3577 = ~new_n529 & new_n3576;
  assign new_n3578 = pc_16_ & new_n530;
  assign new_n3579 = pencrypt_mode_0_ & new_n3578;
  assign new_n3580 = ~new_n529 & new_n3579;
  assign new_n3581 = ~preset_0_ & new_n3580;
  assign new_n3582 = ~pencrypt_0_ & new_n3331;
  assign new_n3583 = new_n529 & new_n3582;
  assign new_n3584 = ~pencrypt_mode_0_ & new_n2144;
  assign new_n3585 = ~new_n529 & new_n3584;
  assign new_n3586 = ~preset_0_ & new_n3585;
  assign new_n3587 = pinreg_50_ & new_n582;
  assign new_n3588 = new_n529 & new_n3587;
  assign new_n3589 = ~new_n3583 & ~new_n3586;
  assign new_n3590 = ~new_n3588 & new_n3589;
  assign new_n3591 = ~new_n3571 & ~new_n3574;
  assign new_n3592 = ~new_n3577 & ~new_n3581;
  assign new_n3593 = new_n3591 & new_n3592;
  assign pc_new_15_ = ~new_n3590 | ~new_n3593;
  assign new_n3595 = pencrypt_mode_0_ & new_n1311;
  assign new_n3596 = ~new_n529 & new_n3595;
  assign new_n3597 = ~preset_0_ & new_n3596;
  assign new_n3598 = ~pencrypt_mode_0_ & new_n2176;
  assign new_n3599 = ~new_n529 & new_n3598;
  assign new_n3600 = ~preset_0_ & new_n3599;
  assign new_n3601 = pencrypt_mode_0_ & new_n1885;
  assign new_n3602 = ~new_n529 & new_n3601;
  assign new_n3603 = ~preset_0_ & new_n3602;
  assign new_n3604 = ~pencrypt_mode_0_ & new_n2874;
  assign new_n3605 = ~new_n529 & new_n3604;
  assign new_n3606 = ~preset_0_ & new_n3605;
  assign new_n3607 = ~preset_0_ & pc_26_;
  assign new_n3608 = ~new_n512 & new_n3607;
  assign new_n3609 = ~new_n529 & new_n3608;
  assign new_n3610 = pinreg_27_ & new_n582;
  assign new_n3611 = new_n529 & new_n3610;
  assign new_n3612 = pinreg_35_ & new_n554;
  assign new_n3613 = new_n529 & new_n3612;
  assign new_n3614 = ~new_n3609 & ~new_n3611;
  assign new_n3615 = ~new_n3613 & new_n3614;
  assign new_n3616 = ~new_n3597 & ~new_n3600;
  assign new_n3617 = ~new_n3603 & ~new_n3606;
  assign new_n3618 = new_n3616 & new_n3617;
  assign pc_new_26_ = ~new_n3615 | ~new_n3618;
  assign new_n3620 = pd_18_ & new_n535;
  assign new_n3621 = pencrypt_mode_0_ & new_n3620;
  assign new_n3622 = ~new_n529 & new_n3621;
  assign new_n3623 = ~preset_0_ & new_n3622;
  assign new_n3624 = ~pencrypt_mode_0_ & new_n2202;
  assign new_n3625 = ~new_n529 & new_n3624;
  assign new_n3626 = ~preset_0_ & new_n3625;
  assign new_n3627 = pd_17_ & new_n530;
  assign new_n3628 = pencrypt_mode_0_ & new_n3627;
  assign new_n3629 = ~new_n529 & new_n3628;
  assign new_n3630 = ~preset_0_ & new_n3629;
  assign new_n3631 = ~pencrypt_mode_0_ & new_n2904;
  assign new_n3632 = ~new_n529 & new_n3631;
  assign new_n3633 = ~preset_0_ & new_n3632;
  assign new_n3634 = ~preset_0_ & pd_16_;
  assign new_n3635 = ~new_n512 & new_n3634;
  assign new_n3636 = ~new_n529 & new_n3635;
  assign new_n3637 = pinreg_44_ & new_n582;
  assign new_n3638 = new_n529 & new_n3637;
  assign new_n3639 = pinreg_52_ & new_n554;
  assign new_n3640 = new_n529 & new_n3639;
  assign new_n3641 = ~new_n3636 & ~new_n3638;
  assign new_n3642 = ~new_n3640 & new_n3641;
  assign new_n3643 = ~new_n3623 & ~new_n3626;
  assign new_n3644 = ~new_n3630 & ~new_n3633;
  assign new_n3645 = new_n3643 & new_n3644;
  assign pd_new_16_ = ~new_n3642 | ~new_n3645;
  assign new_n3647 = pd_26_ & new_n530;
  assign new_n3648 = ~pencrypt_mode_0_ & new_n3647;
  assign new_n3649 = ~new_n529 & new_n3648;
  assign new_n3650 = ~preset_0_ & new_n3649;
  assign new_n3651 = pencrypt_mode_0_ & new_n1127;
  assign new_n3652 = ~new_n529 & new_n3651;
  assign new_n3653 = ~preset_0_ & new_n3652;
  assign new_n3654 = ~preset_0_ & pd_27_;
  assign new_n3655 = ~new_n512 & new_n3654;
  assign new_n3656 = ~new_n529 & new_n3655;
  assign new_n3657 = pencrypt_mode_0_ & new_n1345;
  assign new_n3658 = ~new_n529 & new_n3657;
  assign new_n3659 = ~preset_0_ & new_n3658;
  assign new_n3660 = ~preset_0_ & pdata_in_3_;
  assign new_n3661 = ~pencrypt_0_ & new_n3660;
  assign new_n3662 = new_n529 & new_n3661;
  assign new_n3663 = ~pencrypt_mode_0_ & new_n2235;
  assign new_n3664 = ~new_n529 & new_n3663;
  assign new_n3665 = ~preset_0_ & new_n3664;
  assign new_n3666 = pinreg_54_ & new_n582;
  assign new_n3667 = new_n529 & new_n3666;
  assign new_n3668 = ~new_n3662 & ~new_n3665;
  assign new_n3669 = ~new_n3667 & new_n3668;
  assign new_n3670 = ~new_n3650 & ~new_n3653;
  assign new_n3671 = ~new_n3656 & ~new_n3659;
  assign new_n3672 = new_n3670 & new_n3671;
  assign pd_new_27_ = ~new_n3669 | ~new_n3672;
  assign new_n3674 = pdata_in_1_ & new_n522;
  assign new_n3675 = pdata_39_ & ~new_n522;
  assign pdata_new_7_ = new_n3674 | new_n3675;
  assign new_n3677 = new_n3105 & new_n3109;
  assign new_n3678 = ~new_n3105 & new_n3159;
  assign new_n3679 = ~new_n3105 & new_n3151;
  assign new_n3680 = ~new_n3102 & new_n3118;
  assign new_n3681 = ~new_n3105 & new_n3680;
  assign new_n3682 = ~new_n3105 & new_n3141;
  assign new_n3683 = ~new_n3105 & new_n3172;
  assign new_n3684 = new_n3105 & new_n3161;
  assign new_n3685 = new_n3105 & new_n3154;
  assign new_n3686 = ~new_n3189 & ~new_n3261;
  assign new_n3687 = new_n3193 & new_n3686;
  assign new_n3688 = ~new_n3184 & ~new_n3685;
  assign new_n3689 = ~new_n3252 & ~new_n3257;
  assign new_n3690 = new_n3688 & new_n3689;
  assign new_n3691 = new_n3687 & new_n3690;
  assign new_n3692 = ~new_n3180 & ~new_n3684;
  assign new_n3693 = ~new_n3247 & ~new_n3683;
  assign new_n3694 = new_n3692 & new_n3693;
  assign new_n3695 = ~new_n3160 & ~new_n3167;
  assign new_n3696 = ~new_n3134 & ~new_n3158;
  assign new_n3697 = new_n3695 & new_n3696;
  assign new_n3698 = new_n3694 & new_n3697;
  assign new_n3699 = new_n3691 & new_n3698;
  assign new_n3700 = ~new_n3155 & ~new_n3258;
  assign new_n3701 = ~new_n3174 & ~new_n3682;
  assign new_n3702 = new_n3700 & new_n3701;
  assign new_n3703 = ~new_n3136 & ~new_n3681;
  assign new_n3704 = ~new_n3248 & ~new_n3679;
  assign new_n3705 = new_n3703 & new_n3704;
  assign new_n3706 = new_n3702 & new_n3705;
  assign new_n3707 = ~new_n3115 & ~new_n3242;
  assign new_n3708 = ~new_n3121 & ~new_n3677;
  assign new_n3709 = new_n3707 & new_n3708;
  assign new_n3710 = ~new_n3130 & ~new_n3678;
  assign new_n3711 = new_n3287 & new_n3710;
  assign new_n3712 = new_n3709 & new_n3711;
  assign new_n3713 = new_n3706 & new_n3712;
  assign new_n3714 = new_n3699 & new_n3713;
  assign new_n3715 = ~pdata_17_ & ~new_n3714;
  assign new_n3716 = ~new_n522 & new_n3715;
  assign new_n3717 = pdata_17_ & new_n3714;
  assign new_n3718 = ~new_n522 & new_n3717;
  assign new_n3719 = pinreg_44_ & new_n522;
  assign new_n3720 = ~new_n3716 & ~new_n3718;
  assign pdata_new_49_ = new_n3719 | ~new_n3720;
  assign new_n3722 = ~pcount_0_ & pinreg_26_;
  assign new_n3723 = ~new_n522 & new_n3722;
  assign new_n3724 = pcount_0_ & pinreg_18_;
  assign new_n3725 = ~new_n522 & new_n3724;
  assign pinreg_new_26_ = new_n3723 | new_n3725;
  assign new_n3727 = ~pcount_0_ & pinreg_37_;
  assign new_n3728 = ~new_n522 & new_n3727;
  assign new_n3729 = pcount_0_ & pinreg_29_;
  assign new_n3730 = ~new_n522 & new_n3729;
  assign pinreg_new_37_ = new_n3728 | new_n3730;
  assign new_n3732 = ~pcount_0_ & pinreg_48_;
  assign new_n3733 = ~new_n522 & new_n3732;
  assign new_n3734 = pcount_0_ & pinreg_40_;
  assign new_n3735 = ~new_n522 & new_n3734;
  assign pinreg_new_48_ = new_n3733 | new_n3735;
  assign new_n3737 = new_n522 & new_n3480;
  assign new_n3738 = ~pcount_0_ & poutreg_5_;
  assign new_n3739 = ~new_n522 & new_n3738;
  assign new_n3740 = new_n522 & new_n3478;
  assign new_n3741 = pcount_0_ & poutreg_13_;
  assign new_n3742 = ~new_n522 & new_n3741;
  assign new_n3743 = ~new_n3737 & ~new_n3739;
  assign new_n3744 = ~new_n3740 & ~new_n3742;
  assign poutreg_new_5_ = ~new_n3743 | ~new_n3744;
  assign new_n3746 = ~new_n1382 & new_n1404;
  assign new_n3747 = ~new_n1382 & new_n1441;
  assign new_n3748 = new_n1382 & new_n2279;
  assign new_n3749 = new_n1382 & new_n2283;
  assign new_n3750 = ~new_n2271 & ~new_n2293;
  assign new_n3751 = new_n1468 & new_n3750;
  assign new_n3752 = ~new_n2290 & ~new_n2559;
  assign new_n3753 = ~new_n2289 & ~new_n2291;
  assign new_n3754 = new_n3752 & new_n3753;
  assign new_n3755 = new_n3751 & new_n3754;
  assign new_n3756 = ~new_n2284 & ~new_n3749;
  assign new_n3757 = ~new_n1442 & ~new_n3748;
  assign new_n3758 = new_n3756 & new_n3757;
  assign new_n3759 = ~new_n1416 & ~new_n2286;
  assign new_n3760 = ~new_n1437 & ~new_n2555;
  assign new_n3761 = new_n3759 & new_n3760;
  assign new_n3762 = new_n3758 & new_n3761;
  assign new_n3763 = new_n3755 & new_n3762;
  assign new_n3764 = ~new_n1430 & ~new_n1459;
  assign new_n3765 = ~new_n1444 & ~new_n2558;
  assign new_n3766 = new_n3764 & new_n3765;
  assign new_n3767 = ~new_n1457 & ~new_n3747;
  assign new_n3768 = ~new_n1427 & ~new_n3746;
  assign new_n3769 = new_n3767 & new_n3768;
  assign new_n3770 = new_n3766 & new_n3769;
  assign new_n3771 = ~new_n1392 & ~new_n2552;
  assign new_n3772 = new_n1490 & new_n3771;
  assign new_n3773 = ~new_n1447 & ~new_n2276;
  assign new_n3774 = new_n1492 & new_n3773;
  assign new_n3775 = new_n3772 & new_n3774;
  assign new_n3776 = new_n3770 & new_n3775;
  assign new_n3777 = new_n3763 & new_n3776;
  assign new_n3778 = pdata_20_ & new_n3777;
  assign new_n3779 = new_n522 & new_n3778;
  assign new_n3780 = pcount_0_ & poutreg_37_;
  assign new_n3781 = ~new_n522 & new_n3780;
  assign new_n3782 = ~pdata_20_ & ~new_n3777;
  assign new_n3783 = new_n522 & new_n3782;
  assign new_n3784 = ~pcount_0_ & poutreg_29_;
  assign new_n3785 = ~new_n522 & new_n3784;
  assign new_n3786 = ~new_n3779 & ~new_n3781;
  assign new_n3787 = ~new_n3783 & ~new_n3785;
  assign poutreg_new_29_ = ~new_n3786 | ~new_n3787;
  assign new_n3789 = new_n522 & new_n2326;
  assign new_n3790 = pcount_0_ & poutreg_55_;
  assign new_n3791 = ~new_n522 & new_n3790;
  assign new_n3792 = new_n522 & new_n2324;
  assign new_n3793 = ~pcount_0_ & poutreg_47_;
  assign new_n3794 = ~new_n522 & new_n3793;
  assign new_n3795 = ~new_n3789 & ~new_n3791;
  assign new_n3796 = ~new_n3792 & ~new_n3794;
  assign poutreg_new_47_ = ~new_n3795 | ~new_n3796;
  assign new_n3798 = poutreg_52_ & ~pcount_0_;
  assign new_n3799 = ~new_n522 & new_n3798;
  assign new_n3800 = pcount_0_ & poutreg_60_;
  assign new_n3801 = ~new_n522 & new_n3800;
  assign new_n3802 = pdata_49_ & new_n522;
  assign new_n3803 = ~new_n3799 & ~new_n3801;
  assign poutreg_new_52_ = new_n3802 | ~new_n3803;
  assign new_n3805 = pc_18_ & new_n535;
  assign new_n3806 = pencrypt_mode_0_ & new_n3805;
  assign new_n3807 = ~new_n529 & new_n3806;
  assign new_n3808 = ~preset_0_ & new_n3807;
  assign new_n3809 = ~pencrypt_mode_0_ & new_n2435;
  assign new_n3810 = ~new_n529 & new_n3809;
  assign new_n3811 = ~preset_0_ & new_n3810;
  assign new_n3812 = pc_17_ & new_n530;
  assign new_n3813 = pencrypt_mode_0_ & new_n3812;
  assign new_n3814 = ~new_n529 & new_n3813;
  assign new_n3815 = ~preset_0_ & new_n3814;
  assign new_n3816 = ~pencrypt_mode_0_ & new_n3327;
  assign new_n3817 = ~new_n529 & new_n3816;
  assign new_n3818 = ~preset_0_ & new_n3817;
  assign new_n3819 = ~preset_0_ & pc_16_;
  assign new_n3820 = ~new_n512 & new_n3819;
  assign new_n3821 = ~new_n529 & new_n3820;
  assign new_n3822 = pinreg_42_ & new_n582;
  assign new_n3823 = new_n529 & new_n3822;
  assign new_n3824 = pinreg_50_ & new_n554;
  assign new_n3825 = new_n529 & new_n3824;
  assign new_n3826 = ~new_n3821 & ~new_n3823;
  assign new_n3827 = ~new_n3825 & new_n3826;
  assign new_n3828 = ~new_n3808 & ~new_n3811;
  assign new_n3829 = ~new_n3815 & ~new_n3818;
  assign new_n3830 = new_n3828 & new_n3829;
  assign pc_new_16_ = ~new_n3827 | ~new_n3830;
  assign new_n3832 = pencrypt_mode_0_ & new_n1930;
  assign new_n3833 = ~new_n529 & new_n3832;
  assign new_n3834 = ~preset_0_ & new_n3833;
  assign new_n3835 = ~pencrypt_mode_0_ & new_n2464;
  assign new_n3836 = ~new_n529 & new_n3835;
  assign new_n3837 = ~preset_0_ & new_n3836;
  assign new_n3838 = pc_26_ & new_n530;
  assign new_n3839 = pencrypt_mode_0_ & new_n3838;
  assign new_n3840 = ~new_n529 & new_n3839;
  assign new_n3841 = ~preset_0_ & new_n3840;
  assign new_n3842 = ~pencrypt_mode_0_ & new_n3356;
  assign new_n3843 = ~new_n529 & new_n3842;
  assign new_n3844 = ~preset_0_ & new_n3843;
  assign new_n3845 = ~preset_0_ & pc_25_;
  assign new_n3846 = ~new_n512 & new_n3845;
  assign new_n3847 = ~new_n529 & new_n3846;
  assign new_n3848 = pinreg_35_ & new_n582;
  assign new_n3849 = new_n529 & new_n3848;
  assign new_n3850 = pinreg_43_ & new_n554;
  assign new_n3851 = new_n529 & new_n3850;
  assign new_n3852 = ~new_n3847 & ~new_n3849;
  assign new_n3853 = ~new_n3851 & new_n3852;
  assign new_n3854 = ~new_n3834 & ~new_n3837;
  assign new_n3855 = ~new_n3841 & ~new_n3844;
  assign new_n3856 = new_n3854 & new_n3855;
  assign pc_new_25_ = ~new_n3853 | ~new_n3856;
  assign new_n3858 = ~pencrypt_mode_0_ & new_n3381;
  assign new_n3859 = ~new_n529 & new_n3858;
  assign new_n3860 = ~preset_0_ & new_n3859;
  assign new_n3861 = pencrypt_mode_0_ & new_n849;
  assign new_n3862 = ~new_n529 & new_n3861;
  assign new_n3863 = ~preset_0_ & new_n3862;
  assign new_n3864 = ~preset_0_ & pd_15_;
  assign new_n3865 = ~new_n512 & new_n3864;
  assign new_n3866 = ~new_n529 & new_n3865;
  assign new_n3867 = pd_16_ & new_n530;
  assign new_n3868 = pencrypt_mode_0_ & new_n3867;
  assign new_n3869 = ~new_n529 & new_n3868;
  assign new_n3870 = ~preset_0_ & new_n3869;
  assign new_n3871 = ~pencrypt_0_ & new_n2908;
  assign new_n3872 = new_n529 & new_n3871;
  assign new_n3873 = ~pencrypt_mode_0_ & new_n2492;
  assign new_n3874 = ~new_n529 & new_n3873;
  assign new_n3875 = ~preset_0_ & new_n3874;
  assign new_n3876 = pinreg_52_ & new_n582;
  assign new_n3877 = new_n529 & new_n3876;
  assign new_n3878 = ~new_n3872 & ~new_n3875;
  assign new_n3879 = ~new_n3877 & new_n3878;
  assign new_n3880 = ~new_n3860 & ~new_n3863;
  assign new_n3881 = ~new_n3866 & ~new_n3870;
  assign new_n3882 = new_n3880 & new_n3881;
  assign pd_new_15_ = ~new_n3879 | ~new_n3882;
  assign new_n3884 = pcount_2_ & pcount_0_;
  assign new_n3885 = ~preset_0_ & new_n3884;
  assign new_n3886 = ~pcount_3_ & new_n3885;
  assign new_n3887 = ~new_n529 & new_n3886;
  assign new_n3888 = pcount_1_ & new_n3887;
  assign new_n3889 = pcount_3_ & new_n2260;
  assign new_n3890 = ~new_n529 & new_n3889;
  assign new_n3891 = pcount_3_ & new_n2950;
  assign new_n3892 = ~new_n529 & new_n3891;
  assign new_n3893 = ~pcount_2_ & ~preset_0_;
  assign new_n3894 = pcount_3_ & new_n3893;
  assign new_n3895 = ~new_n529 & new_n3894;
  assign new_n3896 = ~new_n3888 & ~new_n3890;
  assign new_n3897 = ~new_n3892 & ~new_n3895;
  assign pcount_new_3_ = ~new_n3896 | ~new_n3897;
  assign new_n3899 = pinreg_51_ & new_n522;
  assign new_n3900 = pdata_40_ & ~new_n522;
  assign pdata_new_8_ = new_n3899 | new_n3900;
  assign new_n3902 = ~pcount_0_ & pinreg_27_;
  assign new_n3903 = ~new_n522 & new_n3902;
  assign new_n3904 = pcount_0_ & pinreg_19_;
  assign new_n3905 = ~new_n522 & new_n3904;
  assign pinreg_new_27_ = new_n3903 | new_n3905;
  assign new_n3907 = ~pcount_0_ & pinreg_36_;
  assign new_n3908 = ~new_n522 & new_n3907;
  assign new_n3909 = pcount_0_ & pinreg_28_;
  assign new_n3910 = ~new_n522 & new_n3909;
  assign pinreg_new_36_ = new_n3908 | new_n3910;
  assign new_n3912 = ~pcount_0_ & pinreg_49_;
  assign new_n3913 = ~new_n522 & new_n3912;
  assign new_n3914 = pcount_0_ & pinreg_41_;
  assign new_n3915 = ~new_n522 & new_n3914;
  assign pinreg_new_49_ = new_n3913 | new_n3915;
  assign new_n3917 = pcount_0_ & poutreg_14_;
  assign new_n3918 = ~new_n522 & new_n3917;
  assign new_n3919 = ~pcount_0_ & poutreg_6_;
  assign new_n3920 = ~new_n522 & new_n3919;
  assign new_n3921 = pdata_63_ & new_n522;
  assign new_n3922 = ~new_n3918 & ~new_n3920;
  assign poutreg_new_6_ = new_n3921 | ~new_n3922;
  assign new_n3924 = ~pcount_0_ & poutreg_48_;
  assign new_n3925 = ~new_n522 & new_n3924;
  assign new_n3926 = pcount_0_ & poutreg_56_;
  assign new_n3927 = ~new_n522 & new_n3926;
  assign new_n3928 = pdata_33_ & new_n522;
  assign new_n3929 = ~new_n3925 & ~new_n3927;
  assign poutreg_new_48_ = new_n3928 | ~new_n3929;
  assign new_n3931 = new_n2613 & new_n2792;
  assign new_n3932 = ~new_n2613 & new_n2678;
  assign new_n3933 = ~new_n2613 & new_n2675;
  assign new_n3934 = new_n2613 & new_n2783;
  assign new_n3935 = new_n2613 & new_n2772;
  assign new_n3936 = new_n2613 & new_n2788;
  assign new_n3937 = ~new_n2613 & new_n2670;
  assign new_n3938 = ~new_n2613 & new_n2617;
  assign new_n3939 = ~new_n2623 & ~new_n2695;
  assign new_n3940 = ~new_n2693 & ~new_n2791;
  assign new_n3941 = new_n3939 & new_n3940;
  assign new_n3942 = ~new_n2690 & ~new_n2789;
  assign new_n3943 = ~new_n2684 & ~new_n3938;
  assign new_n3944 = new_n3942 & new_n3943;
  assign new_n3945 = new_n3941 & new_n3944;
  assign new_n3946 = ~new_n3936 & ~new_n3937;
  assign new_n3947 = ~new_n2782 & ~new_n3935;
  assign new_n3948 = new_n3946 & new_n3947;
  assign new_n3949 = ~new_n2663 & ~new_n2671;
  assign new_n3950 = ~new_n2662 & ~new_n2668;
  assign new_n3951 = new_n3949 & new_n3950;
  assign new_n3952 = new_n3948 & new_n3951;
  assign new_n3953 = new_n3945 & new_n3952;
  assign new_n3954 = ~new_n2681 & ~new_n2688;
  assign new_n3955 = ~new_n2781 & ~new_n3934;
  assign new_n3956 = new_n3954 & new_n3955;
  assign new_n3957 = ~new_n2656 & ~new_n3933;
  assign new_n3958 = ~new_n2771 & ~new_n3932;
  assign new_n3959 = new_n3957 & new_n3958;
  assign new_n3960 = new_n3956 & new_n3959;
  assign new_n3961 = ~new_n2618 & ~new_n2768;
  assign new_n3962 = ~new_n2628 & ~new_n3931;
  assign new_n3963 = new_n3961 & new_n3962;
  assign new_n3964 = ~new_n2649 & ~new_n2773;
  assign new_n3965 = new_n2818 & new_n3964;
  assign new_n3966 = new_n3963 & new_n3965;
  assign new_n3967 = new_n3960 & new_n3966;
  assign new_n3968 = new_n3953 & new_n3967;
  assign new_n3969 = pdata_9_ & new_n3968;
  assign new_n3970 = new_n522 & new_n3969;
  assign new_n3971 = pcount_0_ & poutreg_59_;
  assign new_n3972 = ~new_n522 & new_n3971;
  assign new_n3973 = ~pdata_9_ & ~new_n3968;
  assign new_n3974 = new_n522 & new_n3973;
  assign new_n3975 = poutreg_51_ & ~pcount_0_;
  assign new_n3976 = ~new_n522 & new_n3975;
  assign new_n3977 = ~new_n3970 & ~new_n3972;
  assign new_n3978 = ~new_n3974 & ~new_n3976;
  assign poutreg_new_51_ = ~new_n3977 | ~new_n3978;
  assign new_n3980 = pencrypt_mode_0_ & new_n2468;
  assign new_n3981 = ~new_n529 & new_n3980;
  assign new_n3982 = ~preset_0_ & new_n3981;
  assign new_n3983 = ~pencrypt_mode_0_ & new_n2839;
  assign new_n3984 = ~new_n529 & new_n3983;
  assign new_n3985 = ~preset_0_ & new_n3984;
  assign new_n3986 = pencrypt_mode_0_ & new_n575;
  assign new_n3987 = ~new_n529 & new_n3986;
  assign new_n3988 = ~preset_0_ & new_n3987;
  assign new_n3989 = ~pencrypt_mode_0_ & new_n3578;
  assign new_n3990 = ~new_n529 & new_n3989;
  assign new_n3991 = ~preset_0_ & new_n3990;
  assign new_n3992 = ~preset_0_ & pc_17_;
  assign new_n3993 = ~new_n512 & new_n3992;
  assign new_n3994 = ~new_n529 & new_n3993;
  assign new_n3995 = pinreg_34_ & new_n582;
  assign new_n3996 = new_n529 & new_n3995;
  assign new_n3997 = pinreg_42_ & new_n554;
  assign new_n3998 = new_n529 & new_n3997;
  assign new_n3999 = ~new_n3994 & ~new_n3996;
  assign new_n4000 = ~new_n3998 & new_n3999;
  assign new_n4001 = ~new_n3982 & ~new_n3985;
  assign new_n4002 = ~new_n3988 & ~new_n3991;
  assign new_n4003 = new_n4001 & new_n4002;
  assign pc_new_17_ = ~new_n4000 | ~new_n4003;
  assign new_n4005 = pencrypt_mode_0_ & new_n3417;
  assign new_n4006 = ~new_n529 & new_n4005;
  assign new_n4007 = ~preset_0_ & new_n4006;
  assign new_n4008 = ~pencrypt_mode_0_ & new_n2897;
  assign new_n4009 = ~new_n529 & new_n4008;
  assign new_n4010 = ~preset_0_ & new_n4009;
  assign new_n4011 = pd_19_ & new_n530;
  assign new_n4012 = pencrypt_mode_0_ & new_n4011;
  assign new_n4013 = ~new_n529 & new_n4012;
  assign new_n4014 = ~preset_0_ & new_n4013;
  assign new_n4015 = ~pencrypt_mode_0_ & new_n3627;
  assign new_n4016 = ~new_n529 & new_n4015;
  assign new_n4017 = ~preset_0_ & new_n4016;
  assign new_n4018 = ~preset_0_ & pd_18_;
  assign new_n4019 = ~new_n512 & new_n4018;
  assign new_n4020 = ~new_n529 & new_n4019;
  assign new_n4021 = pinreg_28_ & new_n582;
  assign new_n4022 = new_n529 & new_n4021;
  assign new_n4023 = pinreg_36_ & new_n554;
  assign new_n4024 = new_n529 & new_n4023;
  assign new_n4025 = ~new_n4020 & ~new_n4022;
  assign new_n4026 = ~new_n4024 & new_n4025;
  assign new_n4027 = ~new_n4007 & ~new_n4010;
  assign new_n4028 = ~new_n4014 & ~new_n4017;
  assign new_n4029 = new_n4027 & new_n4028;
  assign pd_new_18_ = ~new_n4026 | ~new_n4029;
  assign new_n4031 = pencrypt_mode_0_ & new_n1338;
  assign new_n4032 = ~new_n529 & new_n4031;
  assign new_n4033 = ~preset_0_ & new_n4032;
  assign new_n4034 = ~pencrypt_mode_0_ & new_n2923;
  assign new_n4035 = ~new_n529 & new_n4034;
  assign new_n4036 = ~preset_0_ & new_n4035;
  assign new_n4037 = pencrypt_mode_0_ & new_n3647;
  assign new_n4038 = ~new_n529 & new_n4037;
  assign new_n4039 = ~preset_0_ & new_n4038;
  assign new_n4040 = ~pencrypt_mode_0_ & new_n2242;
  assign new_n4041 = ~new_n529 & new_n4040;
  assign new_n4042 = ~preset_0_ & new_n4041;
  assign new_n4043 = ~preset_0_ & pd_25_;
  assign new_n4044 = ~new_n512 & new_n4043;
  assign new_n4045 = ~new_n529 & new_n4044;
  assign new_n4046 = pinreg_11_ & new_n554;
  assign new_n4047 = new_n529 & new_n4046;
  assign new_n4048 = pinreg_3_ & new_n582;
  assign new_n4049 = new_n529 & new_n4048;
  assign new_n4050 = ~new_n4045 & ~new_n4047;
  assign new_n4051 = ~new_n4049 & new_n4050;
  assign new_n4052 = ~new_n4033 & ~new_n4036;
  assign new_n4053 = ~new_n4039 & ~new_n4042;
  assign new_n4054 = new_n4052 & new_n4053;
  assign pd_new_25_ = ~new_n4051 | ~new_n4054;
  assign new_n4056 = pinreg_9_ & new_n522;
  assign new_n4057 = pdata_37_ & ~new_n522;
  assign pdata_new_5_ = new_n4056 | new_n4057;
  assign new_n4059 = ~pcount_0_ & pinreg_28_;
  assign new_n4060 = ~new_n522 & new_n4059;
  assign new_n4061 = pcount_0_ & pinreg_20_;
  assign new_n4062 = ~new_n522 & new_n4061;
  assign pinreg_new_28_ = new_n4060 | new_n4062;
  assign new_n4064 = ~pcount_0_ & pinreg_39_;
  assign new_n4065 = ~new_n522 & new_n4064;
  assign new_n4066 = pcount_0_ & pinreg_31_;
  assign new_n4067 = ~new_n522 & new_n4066;
  assign pinreg_new_39_ = new_n4065 | new_n4067;
  assign new_n4069 = ~pcount_0_ & pinreg_46_;
  assign new_n4070 = ~new_n522 & new_n4069;
  assign new_n4071 = pcount_0_ & pinreg_38_;
  assign new_n4072 = ~new_n522 & new_n4071;
  assign pinreg_new_46_ = new_n4070 | new_n4072;
  assign new_n4074 = new_n522 & new_n3014;
  assign new_n4075 = ~pcount_0_ & poutreg_3_;
  assign new_n4076 = ~new_n522 & new_n4075;
  assign new_n4077 = new_n522 & new_n3012;
  assign new_n4078 = pcount_0_ & poutreg_11_;
  assign new_n4079 = ~new_n522 & new_n4078;
  assign new_n4080 = ~new_n4074 & ~new_n4076;
  assign new_n4081 = ~new_n4077 & ~new_n4079;
  assign poutreg_new_3_ = ~new_n4080 | ~new_n4081;
  assign new_n4083 = new_n1593 & new_n1671;
  assign new_n4084 = new_n1593 & new_n1645;
  assign new_n4085 = new_n1593 & new_n1665;
  assign new_n4086 = ~new_n1593 & new_n1633;
  assign new_n4087 = new_n1593 & new_n1654;
  assign new_n4088 = ~new_n1590 & new_n1670;
  assign new_n4089 = ~new_n1593 & new_n4088;
  assign new_n4090 = new_n1593 & new_n1649;
  assign new_n4091 = ~new_n1593 & new_n1602;
  assign new_n4092 = ~new_n1593 & new_n1663;
  assign new_n4093 = new_n1590 & new_n1629;
  assign new_n4094 = ~new_n1593 & new_n4093;
  assign new_n4095 = new_n1593 & new_n1676;
  assign new_n4096 = ~new_n1590 & new_n1678;
  assign new_n4097 = new_n1593 & new_n4096;
  assign new_n4098 = ~new_n1593 & new_n1658;
  assign new_n4099 = ~new_n1593 & new_n1660;
  assign new_n4100 = ~new_n1593 & new_n1597;
  assign new_n4101 = new_n1593 & new_n4093;
  assign new_n4102 = ~new_n1681 & ~new_n4101;
  assign new_n4103 = ~new_n1677 & ~new_n4100;
  assign new_n4104 = new_n4102 & new_n4103;
  assign new_n4105 = ~new_n1668 & ~new_n1672;
  assign new_n4106 = ~new_n1669 & ~new_n4099;
  assign new_n4107 = new_n4105 & new_n4106;
  assign new_n4108 = new_n4104 & new_n4107;
  assign new_n4109 = ~new_n4097 & ~new_n4098;
  assign new_n4110 = ~new_n1622 & ~new_n4095;
  assign new_n4111 = new_n4109 & new_n4110;
  assign new_n4112 = ~new_n1640 & ~new_n1652;
  assign new_n4113 = ~new_n1650 & ~new_n4094;
  assign new_n4114 = new_n4112 & new_n4113;
  assign new_n4115 = new_n4111 & new_n4114;
  assign new_n4116 = new_n4108 & new_n4115;
  assign new_n4117 = ~new_n1644 & ~new_n1646;
  assign new_n4118 = ~new_n1639 & ~new_n4092;
  assign new_n4119 = new_n4117 & new_n4118;
  assign new_n4120 = ~new_n4090 & ~new_n4091;
  assign new_n4121 = ~new_n4087 & ~new_n4089;
  assign new_n4122 = new_n4120 & new_n4121;
  assign new_n4123 = new_n4119 & new_n4122;
  assign new_n4124 = ~new_n4083 & ~new_n4084;
  assign new_n4125 = new_n1704 & new_n4124;
  assign new_n4126 = ~new_n1613 & ~new_n1620;
  assign new_n4127 = ~new_n4085 & ~new_n4086;
  assign new_n4128 = new_n4126 & new_n4127;
  assign new_n4129 = new_n4125 & new_n4128;
  assign new_n4130 = new_n4123 & new_n4129;
  assign new_n4131 = new_n4116 & new_n4130;
  assign new_n4132 = pdata_18_ & new_n4131;
  assign new_n4133 = new_n522 & new_n4132;
  assign new_n4134 = poutreg_53_ & pcount_0_;
  assign new_n4135 = ~new_n522 & new_n4134;
  assign new_n4136 = ~pdata_18_ & ~new_n4131;
  assign new_n4137 = new_n522 & new_n4136;
  assign new_n4138 = ~pcount_0_ & poutreg_45_;
  assign new_n4139 = ~new_n522 & new_n4138;
  assign new_n4140 = ~new_n4133 & ~new_n4135;
  assign new_n4141 = ~new_n4137 & ~new_n4139;
  assign poutreg_new_45_ = ~new_n4140 | ~new_n4141;
  assign new_n4143 = ~pcount_0_ & poutreg_54_;
  assign new_n4144 = ~new_n522 & new_n4143;
  assign new_n4145 = poutreg_62_ & pcount_0_;
  assign new_n4146 = ~new_n522 & new_n4145;
  assign new_n4147 = pdata_57_ & new_n522;
  assign new_n4148 = ~new_n4144 & ~new_n4146;
  assign poutreg_new_54_ = new_n4147 | ~new_n4148;
  assign new_n4150 = pencrypt_mode_0_ & new_n2190;
  assign new_n4151 = ~new_n529 & new_n4150;
  assign new_n4152 = ~preset_0_ & new_n4151;
  assign new_n4153 = ~pencrypt_mode_0_ & new_n3320;
  assign new_n4154 = ~new_n529 & new_n4153;
  assign new_n4155 = ~preset_0_ & new_n4154;
  assign new_n4156 = pc_19_ & new_n530;
  assign new_n4157 = pencrypt_mode_0_ & new_n4156;
  assign new_n4158 = ~new_n529 & new_n4157;
  assign new_n4159 = ~preset_0_ & new_n4158;
  assign new_n4160 = ~pencrypt_mode_0_ & new_n3812;
  assign new_n4161 = ~new_n529 & new_n4160;
  assign new_n4162 = ~preset_0_ & new_n4161;
  assign new_n4163 = ~preset_0_ & pc_18_;
  assign new_n4164 = ~new_n512 & new_n4163;
  assign new_n4165 = ~new_n529 & new_n4164;
  assign new_n4166 = pinreg_26_ & new_n582;
  assign new_n4167 = new_n529 & new_n4166;
  assign new_n4168 = pinreg_34_ & new_n554;
  assign new_n4169 = new_n529 & new_n4168;
  assign new_n4170 = ~new_n4165 & ~new_n4167;
  assign new_n4171 = ~new_n4169 & new_n4170;
  assign new_n4172 = ~new_n4152 & ~new_n4155;
  assign new_n4173 = ~new_n4159 & ~new_n4162;
  assign new_n4174 = new_n4172 & new_n4173;
  assign pc_new_18_ = ~new_n4171 | ~new_n4174;
  assign new_n4176 = pencrypt_mode_0_ & new_n1525;
  assign new_n4177 = ~new_n529 & new_n4176;
  assign new_n4178 = ~preset_0_ & new_n4177;
  assign new_n4179 = ~pencrypt_mode_0_ & new_n3349;
  assign new_n4180 = ~new_n529 & new_n4179;
  assign new_n4181 = ~preset_0_ & new_n4180;
  assign new_n4182 = pencrypt_mode_0_ & new_n1937;
  assign new_n4183 = ~new_n529 & new_n4182;
  assign new_n4184 = ~preset_0_ & new_n4183;
  assign new_n4185 = ~pencrypt_mode_0_ & new_n3838;
  assign new_n4186 = ~new_n529 & new_n4185;
  assign new_n4187 = ~preset_0_ & new_n4186;
  assign new_n4188 = ~preset_0_ & pc_27_;
  assign new_n4189 = ~new_n512 & new_n4188;
  assign new_n4190 = ~new_n529 & new_n4189;
  assign new_n4191 = pinreg_27_ & new_n554;
  assign new_n4192 = new_n529 & new_n4191;
  assign new_n4193 = pinreg_48_ & new_n582;
  assign new_n4194 = new_n529 & new_n4193;
  assign new_n4195 = ~new_n4190 & ~new_n4192;
  assign new_n4196 = ~new_n4194 & new_n4195;
  assign new_n4197 = ~new_n4178 & ~new_n4181;
  assign new_n4198 = ~new_n4184 & ~new_n4187;
  assign new_n4199 = new_n4197 & new_n4198;
  assign pc_new_27_ = ~new_n4196 | ~new_n4199;
  assign new_n4201 = pencrypt_mode_0_ & new_n2927;
  assign new_n4202 = ~new_n529 & new_n4201;
  assign new_n4203 = ~preset_0_ & new_n4202;
  assign new_n4204 = ~pencrypt_mode_0_ & new_n3373;
  assign new_n4205 = ~new_n529 & new_n4204;
  assign new_n4206 = ~preset_0_ & new_n4205;
  assign new_n4207 = pencrypt_mode_0_ & new_n857;
  assign new_n4208 = ~new_n529 & new_n4207;
  assign new_n4209 = ~preset_0_ & new_n4208;
  assign new_n4210 = ~pencrypt_mode_0_ & new_n3867;
  assign new_n4211 = ~new_n529 & new_n4210;
  assign new_n4212 = ~preset_0_ & new_n4211;
  assign new_n4213 = ~preset_0_ & pd_17_;
  assign new_n4214 = ~new_n512 & new_n4213;
  assign new_n4215 = ~new_n529 & new_n4214;
  assign new_n4216 = pinreg_36_ & new_n582;
  assign new_n4217 = new_n529 & new_n4216;
  assign new_n4218 = pinreg_44_ & new_n554;
  assign new_n4219 = new_n529 & new_n4218;
  assign new_n4220 = ~new_n4215 & ~new_n4217;
  assign new_n4221 = ~new_n4219 & new_n4220;
  assign new_n4222 = ~new_n4203 & ~new_n4206;
  assign new_n4223 = ~new_n4209 & ~new_n4212;
  assign new_n4224 = new_n4222 & new_n4223;
  assign pd_new_17_ = ~new_n4221 | ~new_n4224;
  assign new_n4226 = ~pencrypt_mode_0_ & new_n2528;
  assign new_n4227 = ~new_n529 & new_n4226;
  assign new_n4228 = ~preset_0_ & new_n4227;
  assign new_n4229 = pencrypt_mode_0_ & new_n1552;
  assign new_n4230 = ~new_n529 & new_n4229;
  assign new_n4231 = ~preset_0_ & new_n4230;
  assign new_n4232 = ~preset_0_ & pd_26_;
  assign new_n4233 = ~new_n512 & new_n4232;
  assign new_n4234 = ~new_n529 & new_n4233;
  assign new_n4235 = pencrypt_mode_0_ & new_n1964;
  assign new_n4236 = ~new_n529 & new_n4235;
  assign new_n4237 = ~preset_0_ & new_n4236;
  assign new_n4238 = pencrypt_0_ & new_n3660;
  assign new_n4239 = new_n529 & new_n4238;
  assign new_n4240 = ~pencrypt_mode_0_ & new_n3405;
  assign new_n4241 = ~new_n529 & new_n4240;
  assign new_n4242 = ~preset_0_ & new_n4241;
  assign new_n4243 = pinreg_3_ & new_n554;
  assign new_n4244 = new_n529 & new_n4243;
  assign new_n4245 = ~new_n4239 & ~new_n4242;
  assign new_n4246 = ~new_n4244 & new_n4245;
  assign new_n4247 = ~new_n4228 & ~new_n4231;
  assign new_n4248 = ~new_n4234 & ~new_n4237;
  assign new_n4249 = new_n4247 & new_n4248;
  assign pd_new_26_ = ~new_n4246 | ~new_n4249;
  assign new_n4251 = pinreg_1_ & new_n522;
  assign new_n4252 = pdata_38_ & ~new_n522;
  assign pdata_new_6_ = new_n4251 | new_n4252;
  assign new_n4254 = ~new_n3105 & new_n3166;
  assign new_n4255 = ~new_n3105 & new_n3260;
  assign new_n4256 = ~new_n3105 & new_n3251;
  assign new_n4257 = new_n3105 & new_n3680;
  assign new_n4258 = ~new_n3189 & ~new_n3192;
  assign new_n4259 = ~new_n3257 & ~new_n3259;
  assign new_n4260 = new_n4258 & new_n4259;
  assign new_n4261 = ~new_n3177 & ~new_n3182;
  assign new_n4262 = ~new_n3258 & ~new_n3685;
  assign new_n4263 = new_n4261 & new_n4262;
  assign new_n4264 = new_n4260 & new_n4263;
  assign new_n4265 = ~new_n3174 & ~new_n4257;
  assign new_n4266 = ~new_n3248 & ~new_n4256;
  assign new_n4267 = new_n4265 & new_n4266;
  assign new_n4268 = ~new_n3162 & ~new_n3678;
  assign new_n4269 = new_n3272 & new_n4268;
  assign new_n4270 = new_n4267 & new_n4269;
  assign new_n4271 = new_n4264 & new_n4270;
  assign new_n4272 = ~new_n3152 & ~new_n3180;
  assign new_n4273 = new_n3277 & new_n4272;
  assign new_n4274 = ~new_n3682 & ~new_n4255;
  assign new_n4275 = ~new_n3142 & ~new_n4254;
  assign new_n4276 = new_n4274 & new_n4275;
  assign new_n4277 = new_n4273 & new_n4276;
  assign new_n4278 = ~new_n3191 & ~new_n3243;
  assign new_n4279 = ~new_n3110 & ~new_n3677;
  assign new_n4280 = new_n4278 & new_n4279;
  assign new_n4281 = ~new_n3121 & ~new_n3245;
  assign new_n4282 = ~new_n3127 & ~new_n3136;
  assign new_n4283 = new_n4281 & new_n4282;
  assign new_n4284 = new_n4280 & new_n4283;
  assign new_n4285 = new_n4277 & new_n4284;
  assign new_n4286 = new_n4271 & new_n4285;
  assign new_n4287 = ~pdata_27_ & ~new_n4286;
  assign new_n4288 = ~new_n522 & new_n4287;
  assign new_n4289 = pdata_27_ & new_n4286;
  assign new_n4290 = ~new_n522 & new_n4289;
  assign new_n4291 = pinreg_30_ & new_n522;
  assign new_n4292 = ~new_n4288 & ~new_n4290;
  assign pdata_new_59_ = new_n4291 | ~new_n4292;
  assign new_n4294 = ~pcount_0_ & pinreg_29_;
  assign new_n4295 = ~new_n522 & new_n4294;
  assign new_n4296 = pcount_0_ & pinreg_21_;
  assign new_n4297 = ~new_n522 & new_n4296;
  assign pinreg_new_29_ = new_n4295 | new_n4297;
  assign new_n4299 = ~pcount_0_ & pinreg_38_;
  assign new_n4300 = ~new_n522 & new_n4299;
  assign new_n4301 = pcount_0_ & pinreg_30_;
  assign new_n4302 = ~new_n522 & new_n4301;
  assign pinreg_new_38_ = new_n4300 | new_n4302;
  assign new_n4304 = ~pcount_0_ & pinreg_47_;
  assign new_n4305 = ~new_n522 & new_n4304;
  assign new_n4306 = pcount_0_ & pinreg_39_;
  assign new_n4307 = ~new_n522 & new_n4306;
  assign pinreg_new_47_ = new_n4305 | new_n4307;
  assign new_n4309 = pcount_0_ & poutreg_12_;
  assign new_n4310 = ~new_n522 & new_n4309;
  assign new_n4311 = ~pcount_0_ & poutreg_4_;
  assign new_n4312 = ~new_n522 & new_n4311;
  assign new_n4313 = pdata_55_ & new_n522;
  assign new_n4314 = ~new_n4310 & ~new_n4312;
  assign poutreg_new_4_ = new_n4313 | ~new_n4314;
  assign new_n4316 = new_n522 & new_n4289;
  assign new_n4317 = pcount_0_ & poutreg_47_;
  assign new_n4318 = ~new_n522 & new_n4317;
  assign new_n4319 = new_n522 & new_n4287;
  assign new_n4320 = ~pcount_0_ & poutreg_39_;
  assign new_n4321 = ~new_n522 & new_n4320;
  assign new_n4322 = ~new_n4316 & ~new_n4318;
  assign new_n4323 = ~new_n4319 & ~new_n4321;
  assign poutreg_new_39_ = ~new_n4322 | ~new_n4323;
  assign new_n4325 = ~pcount_0_ & poutreg_46_;
  assign new_n4326 = ~new_n522 & new_n4325;
  assign new_n4327 = pcount_0_ & poutreg_54_;
  assign new_n4328 = ~new_n522 & new_n4327;
  assign new_n4329 = pdata_58_ & new_n522;
  assign new_n4330 = ~new_n4326 & ~new_n4328;
  assign poutreg_new_46_ = new_n4329 | ~new_n4330;
  assign new_n4332 = new_n522 & new_n3717;
  assign new_n4333 = pcount_0_ & poutreg_61_;
  assign new_n4334 = ~new_n522 & new_n4333;
  assign new_n4335 = new_n522 & new_n3715;
  assign new_n4336 = poutreg_53_ & ~pcount_0_;
  assign new_n4337 = ~new_n522 & new_n4336;
  assign new_n4338 = ~new_n4332 & ~new_n4334;
  assign new_n4339 = ~new_n4335 & ~new_n4337;
  assign poutreg_new_53_ = ~new_n4338 | ~new_n4339;
  assign new_n4341 = ~pcount_0_ & poutreg_60_;
  assign new_n4342 = ~new_n522 & new_n4341;
  assign new_n4343 = pdata_48_ & new_n522;
  assign poutreg_new_60_ = new_n4342 | new_n4343;
  assign new_n4345 = ~new_n522 & new_n4136;
  assign new_n4346 = ~new_n522 & new_n4132;
  assign new_n4347 = pinreg_36_ & new_n522;
  assign new_n4348 = ~new_n4345 & ~new_n4346;
  assign pdata_new_50_ = new_n4347 | ~new_n4348;
  assign new_n4350 = ~new_n522 & new_n1222;
  assign new_n4351 = ~new_n522 & new_n1218;
  assign new_n4352 = pdata_in_6_ & new_n522;
  assign new_n4353 = ~new_n4350 & ~new_n4351;
  assign pdata_new_63_ = new_n4352 | ~new_n4353;
  assign new_n4355 = ~pcount_0_ & poutreg_30_;
  assign new_n4356 = ~new_n522 & new_n4355;
  assign new_n4357 = pcount_0_ & poutreg_38_;
  assign new_n4358 = ~new_n522 & new_n4357;
  assign new_n4359 = pdata_60_ & new_n522;
  assign new_n4360 = ~new_n4356 & ~new_n4358;
  assign poutreg_new_30_ = new_n4359 | ~new_n4360;
  assign new_n4362 = new_n1593 & new_n1667;
  assign new_n4363 = ~new_n1593 & new_n4096;
  assign new_n4364 = ~new_n1593 & new_n1621;
  assign new_n4365 = ~new_n1593 & new_n1612;
  assign new_n4366 = new_n1593 & new_n1673;
  assign new_n4367 = new_n1593 & new_n1643;
  assign new_n4368 = new_n1590 & new_n1648;
  assign new_n4369 = ~new_n1593 & new_n4368;
  assign new_n4370 = new_n1593 & new_n1619;
  assign new_n4371 = ~new_n1681 & ~new_n4084;
  assign new_n4372 = new_n1683 & new_n4371;
  assign new_n4373 = ~new_n1642 & ~new_n4100;
  assign new_n4374 = ~new_n4369 & ~new_n4370;
  assign new_n4375 = new_n4373 & new_n4374;
  assign new_n4376 = new_n4372 & new_n4375;
  assign new_n4377 = ~new_n4098 & ~new_n4367;
  assign new_n4378 = ~new_n1622 & ~new_n4366;
  assign new_n4379 = new_n4377 & new_n4378;
  assign new_n4380 = ~new_n1650 & ~new_n1659;
  assign new_n4381 = ~new_n1624 & ~new_n4094;
  assign new_n4382 = new_n4380 & new_n4381;
  assign new_n4383 = new_n4379 & new_n4382;
  assign new_n4384 = new_n4376 & new_n4383;
  assign new_n4385 = ~new_n1640 & ~new_n1646;
  assign new_n4386 = ~new_n1655 & ~new_n1669;
  assign new_n4387 = new_n4385 & new_n4386;
  assign new_n4388 = ~new_n1634 & ~new_n4365;
  assign new_n4389 = ~new_n4090 & ~new_n4364;
  assign new_n4390 = new_n4388 & new_n4389;
  assign new_n4391 = new_n4387 & new_n4390;
  assign new_n4392 = ~new_n1680 & ~new_n4083;
  assign new_n4393 = ~new_n1613 & ~new_n4362;
  assign new_n4394 = new_n4392 & new_n4393;
  assign new_n4395 = ~new_n1608 & ~new_n4363;
  assign new_n4396 = ~new_n4086 & ~new_n4087;
  assign new_n4397 = new_n4395 & new_n4396;
  assign new_n4398 = new_n4394 & new_n4397;
  assign new_n4399 = new_n4391 & new_n4398;
  assign new_n4400 = new_n4384 & new_n4399;
  assign new_n4401 = pdata_10_ & new_n4400;
  assign new_n4402 = new_n522 & new_n4401;
  assign new_n4403 = poutreg_51_ & pcount_0_;
  assign new_n4404 = ~new_n522 & new_n4403;
  assign new_n4405 = ~pdata_10_ & ~new_n4400;
  assign new_n4406 = new_n522 & new_n4405;
  assign new_n4407 = ~pcount_0_ & poutreg_43_;
  assign new_n4408 = ~new_n522 & new_n4407;
  assign new_n4409 = ~new_n4402 & ~new_n4404;
  assign new_n4410 = ~new_n4406 & ~new_n4408;
  assign poutreg_new_43_ = ~new_n4409 | ~new_n4410;
  assign new_n4412 = ~pcount_0_ & poutreg_56_;
  assign new_n4413 = ~new_n522 & new_n4412;
  assign new_n4414 = pdata_32_ & new_n522;
  assign poutreg_new_56_ = new_n4413 | new_n4414;
  assign new_n4416 = ~pcount_0_ & poutreg_44_;
  assign new_n4417 = ~new_n522 & new_n4416;
  assign new_n4418 = poutreg_52_ & pcount_0_;
  assign new_n4419 = ~new_n522 & new_n4418;
  assign new_n4420 = pdata_50_ & new_n522;
  assign new_n4421 = ~new_n4417 & ~new_n4419;
  assign poutreg_new_44_ = new_n4420 | ~new_n4421;
  assign new_n4423 = new_n522 & new_n2729;
  assign new_n4424 = poutreg_63_ & pcount_0_;
  assign new_n4425 = ~new_n522 & new_n4424;
  assign new_n4426 = new_n522 & new_n2727;
  assign new_n4427 = ~pcount_0_ & poutreg_55_;
  assign new_n4428 = ~new_n522 & new_n4427;
  assign new_n4429 = ~new_n4423 & ~new_n4425;
  assign new_n4430 = ~new_n4426 & ~new_n4428;
  assign poutreg_new_55_ = ~new_n4429 | ~new_n4430;
  assign new_n4432 = ~new_n1998 & new_n2064;
  assign new_n4433 = ~new_n1998 & new_n2970;
  assign new_n4434 = new_n1998 & new_n2052;
  assign new_n4435 = new_n1998 & new_n2975;
  assign new_n4436 = ~new_n2070 & ~new_n2082;
  assign new_n4437 = new_n2087 & new_n4436;
  assign new_n4438 = ~new_n2072 & ~new_n3450;
  assign new_n4439 = new_n2986 & new_n4438;
  assign new_n4440 = new_n4437 & new_n4439;
  assign new_n4441 = ~new_n3449 & ~new_n4435;
  assign new_n4442 = ~new_n2025 & ~new_n4434;
  assign new_n4443 = new_n4441 & new_n4442;
  assign new_n4444 = ~new_n2059 & ~new_n2978;
  assign new_n4445 = new_n2993 & new_n4444;
  assign new_n4446 = new_n4443 & new_n4445;
  assign new_n4447 = new_n4440 & new_n4446;
  assign new_n4448 = ~new_n2048 & ~new_n2974;
  assign new_n4449 = new_n2998 & new_n4448;
  assign new_n4450 = ~new_n3446 & ~new_n4433;
  assign new_n4451 = ~new_n2039 & ~new_n4432;
  assign new_n4452 = new_n4450 & new_n4451;
  assign new_n4453 = new_n4449 & new_n4452;
  assign new_n4454 = ~new_n2964 & ~new_n2965;
  assign new_n4455 = new_n2110 & new_n4454;
  assign new_n4456 = ~new_n2030 & ~new_n3443;
  assign new_n4457 = ~new_n2032 & ~new_n2056;
  assign new_n4458 = new_n4456 & new_n4457;
  assign new_n4459 = new_n4455 & new_n4458;
  assign new_n4460 = new_n4453 & new_n4459;
  assign new_n4461 = new_n4447 & new_n4460;
  assign new_n4462 = ~pdata_29_ & ~new_n4461;
  assign new_n4463 = ~new_n522 & new_n4462;
  assign new_n4464 = pdata_29_ & new_n4461;
  assign new_n4465 = ~new_n522 & new_n4464;
  assign new_n4466 = pinreg_14_ & new_n522;
  assign new_n4467 = ~new_n4463 & ~new_n4465;
  assign pdata_new_61_ = new_n4466 | ~new_n4467;
  assign new_n4469 = ~pcount_3_ & pencrypt_mode_0_;
  assign new_n4470 = pcount_3_ & pcount_2_;
  assign new_n4471 = pcount_0_ & new_n4470;
  assign new_n4472 = pcount_1_ & new_n4471;
  assign new_n4473 = pencrypt_0_ & new_n4472;
  assign new_n4474 = ~pcount_1_ & pencrypt_mode_0_;
  assign new_n4475 = ~pcount_2_ & pencrypt_mode_0_;
  assign new_n4476 = ~pcount_0_ & pencrypt_mode_0_;
  assign new_n4477 = ~new_n4469 & ~new_n4473;
  assign new_n4478 = ~new_n4474 & new_n4477;
  assign new_n4479 = ~new_n4475 & ~new_n4476;
  assign pencrypt_mode_new_0_ = ~new_n4478 | ~new_n4479;
  assign new_n4481 = ~new_n897 & new_n961;
  assign new_n4482 = ~new_n897 & new_n1035;
  assign new_n4483 = new_n897 & new_n975;
  assign new_n4484 = new_n897 & new_n946;
  assign new_n4485 = ~new_n907 & ~new_n982;
  assign new_n4486 = ~new_n979 & ~new_n1053;
  assign new_n4487 = new_n4485 & new_n4486;
  assign new_n4488 = ~new_n969 & ~new_n974;
  assign new_n4489 = ~new_n1052 & ~new_n3023;
  assign new_n4490 = new_n4488 & new_n4489;
  assign new_n4491 = new_n4487 & new_n4490;
  assign new_n4492 = ~new_n968 & ~new_n4484;
  assign new_n4493 = ~new_n924 & ~new_n4483;
  assign new_n4494 = new_n4492 & new_n4493;
  assign new_n4495 = ~new_n951 & ~new_n955;
  assign new_n4496 = ~new_n926 & ~new_n950;
  assign new_n4497 = new_n4495 & new_n4496;
  assign new_n4498 = new_n4494 & new_n4497;
  assign new_n4499 = new_n4491 & new_n4498;
  assign new_n4500 = ~new_n958 & ~new_n1040;
  assign new_n4501 = new_n3041 & new_n4500;
  assign new_n4502 = ~new_n937 & ~new_n4482;
  assign new_n4503 = ~new_n929 & ~new_n4481;
  assign new_n4504 = new_n4502 & new_n4503;
  assign new_n4505 = new_n4501 & new_n4504;
  assign new_n4506 = ~new_n902 & ~new_n3019;
  assign new_n4507 = ~new_n917 & ~new_n1032;
  assign new_n4508 = new_n4506 & new_n4507;
  assign new_n4509 = ~new_n1038 & ~new_n1048;
  assign new_n4510 = new_n3050 & new_n4509;
  assign new_n4511 = new_n4508 & new_n4510;
  assign new_n4512 = new_n4505 & new_n4511;
  assign new_n4513 = new_n4499 & new_n4512;
  assign new_n4514 = pdata_2_ & new_n4513;
  assign new_n4515 = new_n522 & new_n4514;
  assign new_n4516 = pcount_0_ & poutreg_49_;
  assign new_n4517 = ~new_n522 & new_n4516;
  assign new_n4518 = ~pdata_2_ & ~new_n4513;
  assign new_n4519 = new_n522 & new_n4518;
  assign new_n4520 = ~pcount_0_ & poutreg_41_;
  assign new_n4521 = ~new_n522 & new_n4520;
  assign new_n4522 = ~new_n4515 & ~new_n4517;
  assign new_n4523 = ~new_n4519 & ~new_n4521;
  assign poutreg_new_41_ = ~new_n4522 | ~new_n4523;
  assign new_n4525 = ~pcount_0_ & poutreg_58_;
  assign new_n4526 = ~new_n522 & new_n4525;
  assign new_n4527 = pdata_40_ & new_n522;
  assign poutreg_new_58_ = new_n4526 | new_n4527;
  assign new_n4529 = new_n1747 & new_n2393;
  assign new_n4530 = ~new_n1744 & new_n1759;
  assign new_n4531 = new_n1747 & new_n4530;
  assign new_n4532 = ~new_n1747 & new_n2385;
  assign new_n4533 = ~new_n1747 & new_n1765;
  assign new_n4534 = ~new_n1747 & new_n1775;
  assign new_n4535 = new_n1747 & new_n1792;
  assign new_n4536 = ~new_n1744 & new_n1815;
  assign new_n4537 = new_n1747 & new_n4536;
  assign new_n4538 = ~new_n1747 & new_n1773;
  assign new_n4539 = ~new_n1830 & ~new_n4538;
  assign new_n4540 = ~new_n1832 & ~new_n2392;
  assign new_n4541 = new_n4539 & new_n4540;
  assign new_n4542 = ~new_n1828 & ~new_n2386;
  assign new_n4543 = ~new_n1796 & ~new_n1827;
  assign new_n4544 = new_n4542 & new_n4543;
  assign new_n4545 = new_n4541 & new_n4544;
  assign new_n4546 = ~new_n1804 & ~new_n4537;
  assign new_n4547 = ~new_n2382 & ~new_n4535;
  assign new_n4548 = new_n4546 & new_n4547;
  assign new_n4549 = ~new_n1806 & ~new_n4534;
  assign new_n4550 = ~new_n1801 & ~new_n1808;
  assign new_n4551 = new_n4549 & new_n4550;
  assign new_n4552 = new_n4548 & new_n4551;
  assign new_n4553 = new_n4545 & new_n4552;
  assign new_n4554 = ~new_n1811 & ~new_n2391;
  assign new_n4555 = new_n2406 & new_n4554;
  assign new_n4556 = ~new_n1789 & ~new_n4533;
  assign new_n4557 = ~new_n4531 & ~new_n4532;
  assign new_n4558 = new_n4556 & new_n4557;
  assign new_n4559 = new_n4555 & new_n4558;
  assign new_n4560 = ~new_n1752 & ~new_n2396;
  assign new_n4561 = ~new_n1761 & ~new_n2378;
  assign new_n4562 = new_n4560 & new_n4561;
  assign new_n4563 = ~new_n2380 & ~new_n4529;
  assign new_n4564 = ~new_n1779 & ~new_n1809;
  assign new_n4565 = new_n4563 & new_n4564;
  assign new_n4566 = new_n4562 & new_n4565;
  assign new_n4567 = new_n4559 & new_n4566;
  assign new_n4568 = new_n4553 & new_n4567;
  assign new_n4569 = ~pdata_8_ & ~new_n4568;
  assign new_n4570 = ~new_n522 & new_n4569;
  assign new_n4571 = pdata_8_ & new_n4568;
  assign new_n4572 = ~new_n522 & new_n4571;
  assign new_n4573 = pinreg_50_ & new_n522;
  assign new_n4574 = ~new_n4570 & ~new_n4572;
  assign pdata_new_40_ = new_n4573 | ~new_n4574;
  assign new_n4576 = ~new_n522 & new_n1868;
  assign new_n4577 = ~new_n522 & new_n1864;
  assign new_n4578 = pinreg_6_ & new_n522;
  assign new_n4579 = ~new_n4576 & ~new_n4577;
  assign pdata_new_62_ = new_n4578 | ~new_n4579;
  assign new_n4581 = ~pcount_0_ & poutreg_20_;
  assign new_n4582 = ~new_n522 & new_n4581;
  assign new_n4583 = pcount_0_ & poutreg_28_;
  assign new_n4584 = ~new_n522 & new_n4583;
  assign new_n4585 = pdata_53_ & new_n522;
  assign new_n4586 = ~new_n4582 & ~new_n4584;
  assign poutreg_new_20_ = new_n4585 | ~new_n4586;
  assign new_n4588 = ~pcount_0_ & poutreg_42_;
  assign new_n4589 = ~new_n522 & new_n4588;
  assign new_n4590 = pcount_0_ & poutreg_50_;
  assign new_n4591 = ~new_n522 & new_n4590;
  assign new_n4592 = pdata_42_ & new_n522;
  assign new_n4593 = ~new_n4589 & ~new_n4591;
  assign poutreg_new_42_ = new_n4592 | ~new_n4593;
  assign new_n4595 = ~new_n2613 & new_n2622;
  assign new_n4596 = ~new_n2613 & new_n2648;
  assign new_n4597 = new_n2613 & new_n2777;
  assign new_n4598 = new_n2613 & new_n2774;
  assign new_n4599 = new_n2697 & new_n3939;
  assign new_n4600 = ~new_n2793 & ~new_n3938;
  assign new_n4601 = new_n2797 & new_n4600;
  assign new_n4602 = new_n4599 & new_n4601;
  assign new_n4603 = ~new_n3937 & ~new_n4598;
  assign new_n4604 = ~new_n2649 & ~new_n4597;
  assign new_n4605 = new_n4603 & new_n4604;
  assign new_n4606 = ~new_n2672 & ~new_n2674;
  assign new_n4607 = ~new_n2665 & ~new_n2784;
  assign new_n4608 = new_n4606 & new_n4607;
  assign new_n4609 = new_n4605 & new_n4608;
  assign new_n4610 = new_n4602 & new_n4609;
  assign new_n4611 = ~new_n2681 & ~new_n2789;
  assign new_n4612 = ~new_n2658 & ~new_n3934;
  assign new_n4613 = new_n4611 & new_n4612;
  assign new_n4614 = ~new_n2656 & ~new_n4596;
  assign new_n4615 = ~new_n2652 & ~new_n4595;
  assign new_n4616 = new_n4614 & new_n4615;
  assign new_n4617 = new_n4613 & new_n4616;
  assign new_n4618 = ~new_n2631 & ~new_n2769;
  assign new_n4619 = ~new_n2636 & ~new_n3931;
  assign new_n4620 = new_n4618 & new_n4619;
  assign new_n4621 = ~new_n2770 & ~new_n2773;
  assign new_n4622 = ~new_n2668 & ~new_n2771;
  assign new_n4623 = new_n4621 & new_n4622;
  assign new_n4624 = new_n4620 & new_n4623;
  assign new_n4625 = new_n4617 & new_n4624;
  assign new_n4626 = new_n4610 & new_n4625;
  assign new_n4627 = ~pdata_0_ & ~new_n4626;
  assign new_n4628 = new_n522 & new_n4627;
  assign new_n4629 = pdata_0_ & new_n4626;
  assign new_n4630 = new_n522 & new_n4629;
  assign new_n4631 = ~pcount_0_ & poutreg_57_;
  assign new_n4632 = ~new_n522 & new_n4631;
  assign new_n4633 = ~new_n4628 & ~new_n4630;
  assign poutreg_new_57_ = new_n4632 | ~new_n4633;
  assign new_n4635 = ~new_n522 & new_n3973;
  assign new_n4636 = ~new_n522 & new_n3969;
  assign new_n4637 = pinreg_42_ & new_n522;
  assign new_n4638 = ~new_n4635 & ~new_n4636;
  assign pdata_new_41_ = new_n4637 | ~new_n4638;
  assign new_n4640 = ~new_n1747 & new_n1810;
  assign new_n4641 = ~new_n1747 & new_n4536;
  assign new_n4642 = new_n1747 & new_n1784;
  assign new_n4643 = new_n1747 & new_n2395;
  assign new_n4644 = ~new_n2396 & ~new_n4538;
  assign new_n4645 = ~new_n1832 & ~new_n2394;
  assign new_n4646 = new_n4644 & new_n4645;
  assign new_n4647 = ~new_n1822 & ~new_n2388;
  assign new_n4648 = ~new_n1799 & ~new_n2386;
  assign new_n4649 = new_n4647 & new_n4648;
  assign new_n4650 = new_n4646 & new_n4649;
  assign new_n4651 = ~new_n2387 & ~new_n4643;
  assign new_n4652 = ~new_n1776 & ~new_n4642;
  assign new_n4653 = new_n4651 & new_n4652;
  assign new_n4654 = ~new_n1814 & ~new_n2381;
  assign new_n4655 = ~new_n1779 & ~new_n1806;
  assign new_n4656 = new_n4654 & new_n4655;
  assign new_n4657 = new_n4653 & new_n4656;
  assign new_n4658 = new_n4650 & new_n4657;
  assign new_n4659 = ~new_n1801 & ~new_n1811;
  assign new_n4660 = ~new_n1804 & ~new_n4534;
  assign new_n4661 = new_n4659 & new_n4660;
  assign new_n4662 = ~new_n1823 & ~new_n4641;
  assign new_n4663 = ~new_n1789 & ~new_n4640;
  assign new_n4664 = new_n4662 & new_n4663;
  assign new_n4665 = new_n4661 & new_n4664;
  assign new_n4666 = ~new_n1766 & ~new_n2377;
  assign new_n4667 = new_n1855 & new_n4666;
  assign new_n4668 = ~new_n1774 & ~new_n4531;
  assign new_n4669 = new_n4563 & new_n4668;
  assign new_n4670 = new_n4667 & new_n4669;
  assign new_n4671 = new_n4665 & new_n4670;
  assign new_n4672 = new_n4658 & new_n4671;
  assign new_n4673 = ~pdata_22_ & ~new_n4672;
  assign new_n4674 = ~new_n522 & new_n4673;
  assign new_n4675 = pdata_22_ & new_n4672;
  assign new_n4676 = ~new_n522 & new_n4675;
  assign new_n4677 = pinreg_4_ & new_n522;
  assign new_n4678 = ~new_n4674 & ~new_n4676;
  assign pdata_new_54_ = new_n4677 | ~new_n4678;
  assign new_n4680 = ~pcount_0_ & pinreg_40_;
  assign new_n4681 = ~new_n522 & new_n4680;
  assign new_n4682 = pcount_0_ & pinreg_32_;
  assign new_n4683 = ~new_n522 & new_n4682;
  assign pinreg_new_40_ = new_n4681 | new_n4683;
  assign new_n4685 = ~pcount_0_ & pinreg_51_;
  assign new_n4686 = ~new_n522 & new_n4685;
  assign new_n4687 = pcount_0_ & pinreg_43_;
  assign new_n4688 = ~new_n522 & new_n4687;
  assign pinreg_new_51_ = new_n4686 | new_n4688;
  assign new_n4690 = ~new_n655 & new_n742;
  assign new_n4691 = ~new_n655 & new_n703;
  assign new_n4692 = new_n655 & new_n1172;
  assign new_n4693 = new_n655 & new_n737;
  assign new_n4694 = ~new_n1188 & ~new_n3527;
  assign new_n4695 = ~new_n734 & ~new_n738;
  assign new_n4696 = new_n4694 & new_n4695;
  assign new_n4697 = ~new_n732 & ~new_n1186;
  assign new_n4698 = ~new_n1187 & ~new_n3522;
  assign new_n4699 = new_n4697 & new_n4698;
  assign new_n4700 = new_n4696 & new_n4699;
  assign new_n4701 = ~new_n3526 & ~new_n4693;
  assign new_n4702 = ~new_n685 & ~new_n4692;
  assign new_n4703 = new_n4701 & new_n4702;
  assign new_n4704 = ~new_n706 & ~new_n714;
  assign new_n4705 = new_n3539 & new_n4704;
  assign new_n4706 = new_n4703 & new_n4705;
  assign new_n4707 = new_n4700 & new_n4706;
  assign new_n4708 = ~new_n712 & ~new_n727;
  assign new_n4709 = new_n1203 & new_n4708;
  assign new_n4710 = ~new_n1180 & ~new_n4691;
  assign new_n4711 = ~new_n1177 & ~new_n4690;
  assign new_n4712 = new_n4710 & new_n4711;
  assign new_n4713 = new_n4709 & new_n4712;
  assign new_n4714 = ~new_n660 & ~new_n740;
  assign new_n4715 = new_n1210 & new_n4714;
  assign new_n4716 = new_n769 & new_n3553;
  assign new_n4717 = new_n4715 & new_n4716;
  assign new_n4718 = new_n4713 & new_n4717;
  assign new_n4719 = new_n4707 & new_n4718;
  assign new_n4720 = pdata_21_ & new_n4719;
  assign new_n4721 = new_n522 & new_n4720;
  assign new_n4722 = pcount_0_ & poutreg_29_;
  assign new_n4723 = ~new_n522 & new_n4722;
  assign new_n4724 = ~pdata_21_ & ~new_n4719;
  assign new_n4725 = new_n522 & new_n4724;
  assign new_n4726 = ~pcount_0_ & poutreg_21_;
  assign new_n4727 = ~new_n522 & new_n4726;
  assign new_n4728 = ~new_n4721 & ~new_n4723;
  assign new_n4729 = ~new_n4725 & ~new_n4727;
  assign poutreg_new_21_ = ~new_n4728 | ~new_n4729;
  assign new_n4731 = ~pcount_0_ & poutreg_34_;
  assign new_n4732 = ~new_n522 & new_n4731;
  assign new_n4733 = pcount_0_ & poutreg_42_;
  assign new_n4734 = ~new_n522 & new_n4733;
  assign new_n4735 = pdata_43_ & new_n522;
  assign new_n4736 = ~new_n4732 & ~new_n4734;
  assign poutreg_new_34_ = new_n4735 | ~new_n4736;
  assign new_n4738 = pencrypt_mode_0_ & new_n2524;
  assign new_n4739 = ~new_n529 & new_n4738;
  assign new_n4740 = ~preset_0_ & new_n4739;
  assign new_n4741 = ~pencrypt_mode_0_ & new_n3620;
  assign new_n4742 = ~new_n529 & new_n4741;
  assign new_n4743 = ~preset_0_ & new_n4742;
  assign new_n4744 = pencrypt_mode_0_ & new_n3401;
  assign new_n4745 = ~new_n529 & new_n4744;
  assign new_n4746 = ~preset_0_ & new_n4745;
  assign new_n4747 = ~pencrypt_mode_0_ & new_n4011;
  assign new_n4748 = ~new_n529 & new_n4747;
  assign new_n4749 = ~preset_0_ & new_n4748;
  assign new_n4750 = pd_20_ & ~preset_0_;
  assign new_n4751 = ~new_n512 & new_n4750;
  assign new_n4752 = ~new_n529 & new_n4751;
  assign new_n4753 = pinreg_12_ & new_n582;
  assign new_n4754 = new_n529 & new_n4753;
  assign new_n4755 = pinreg_20_ & new_n554;
  assign new_n4756 = new_n529 & new_n4755;
  assign new_n4757 = ~new_n4752 & ~new_n4754;
  assign new_n4758 = ~new_n4756 & new_n4757;
  assign new_n4759 = ~new_n4740 & ~new_n4743;
  assign new_n4760 = ~new_n4746 & ~new_n4749;
  assign new_n4761 = new_n4759 & new_n4760;
  assign pd_new_20_ = ~new_n4758 | ~new_n4761;
  assign new_n4763 = pinreg_49_ & new_n522;
  assign new_n4764 = pdata_32_ & ~new_n522;
  assign pdata_new_0_ = new_n4763 | new_n4764;
  assign new_n4766 = ~new_n522 & new_n4405;
  assign new_n4767 = ~new_n522 & new_n4401;
  assign new_n4768 = pinreg_34_ & new_n522;
  assign new_n4769 = ~new_n4766 & ~new_n4767;
  assign pdata_new_42_ = new_n4768 | ~new_n4769;
  assign new_n4771 = ~new_n522 & new_n4724;
  assign new_n4772 = ~new_n522 & new_n4720;
  assign new_n4773 = pinreg_12_ & new_n522;
  assign new_n4774 = ~new_n4771 & ~new_n4772;
  assign pdata_new_53_ = new_n4773 | ~new_n4774;
  assign new_n4776 = ~new_n1593 & new_n1651;
  assign new_n4777 = ~new_n1593 & new_n1607;
  assign new_n4778 = new_n1593 & new_n1641;
  assign new_n4779 = new_n1593 & new_n4088;
  assign new_n4780 = ~new_n4084 & ~new_n4101;
  assign new_n4781 = new_n4103 & new_n4780;
  assign new_n4782 = ~new_n1674 & ~new_n4369;
  assign new_n4783 = ~new_n4099 & ~new_n4370;
  assign new_n4784 = new_n4782 & new_n4783;
  assign new_n4785 = new_n4781 & new_n4784;
  assign new_n4786 = ~new_n1666 & ~new_n4779;
  assign new_n4787 = ~new_n1622 & ~new_n4778;
  assign new_n4788 = new_n4786 & new_n4787;
  assign new_n4789 = ~new_n1624 & ~new_n1659;
  assign new_n4790 = ~new_n1642 & ~new_n4086;
  assign new_n4791 = new_n4789 & new_n4790;
  assign new_n4792 = new_n4788 & new_n4791;
  assign new_n4793 = new_n4785 & new_n4792;
  assign new_n4794 = ~new_n1672 & ~new_n4092;
  assign new_n4795 = new_n1698 & new_n4794;
  assign new_n4796 = ~new_n4090 & ~new_n4777;
  assign new_n4797 = ~new_n1627 & ~new_n4776;
  assign new_n4798 = new_n4796 & new_n4797;
  assign new_n4799 = new_n4795 & new_n4798;
  assign new_n4800 = ~new_n1603 & ~new_n1680;
  assign new_n4801 = new_n4393 & new_n4800;
  assign new_n4802 = ~new_n4085 & ~new_n4363;
  assign new_n4803 = new_n1707 & new_n4802;
  assign new_n4804 = new_n4801 & new_n4803;
  assign new_n4805 = new_n4799 & new_n4804;
  assign new_n4806 = new_n4793 & new_n4805;
  assign new_n4807 = ~pdata_28_ & ~new_n4806;
  assign new_n4808 = ~new_n522 & new_n4807;
  assign new_n4809 = pdata_28_ & new_n4806;
  assign new_n4810 = ~new_n522 & new_n4809;
  assign new_n4811 = pinreg_22_ & new_n522;
  assign new_n4812 = ~new_n4808 & ~new_n4810;
  assign pdata_new_60_ = new_n4811 | ~new_n4812;
  assign new_n4814 = ~pcount_0_ & pinreg_41_;
  assign new_n4815 = ~new_n522 & new_n4814;
  assign new_n4816 = pcount_0_ & pinreg_33_;
  assign new_n4817 = ~new_n522 & new_n4816;
  assign pinreg_new_41_ = new_n4815 | new_n4817;
  assign new_n4819 = ~pcount_0_ & pinreg_50_;
  assign new_n4820 = ~new_n522 & new_n4819;
  assign new_n4821 = pcount_0_ & pinreg_42_;
  assign new_n4822 = ~new_n522 & new_n4821;
  assign pinreg_new_50_ = new_n4820 | new_n4822;
  assign new_n4824 = ~pcount_0_ & poutreg_22_;
  assign new_n4825 = ~new_n522 & new_n4824;
  assign new_n4826 = pcount_0_ & poutreg_30_;
  assign new_n4827 = ~new_n522 & new_n4826;
  assign new_n4828 = pdata_61_ & new_n522;
  assign new_n4829 = ~new_n4825 & ~new_n4827;
  assign poutreg_new_22_ = new_n4828 | ~new_n4829;
  assign new_n4831 = new_n522 & new_n1715;
  assign new_n4832 = pcount_0_ & poutreg_41_;
  assign new_n4833 = ~new_n522 & new_n4832;
  assign new_n4834 = new_n522 & new_n1713;
  assign new_n4835 = ~pcount_0_ & poutreg_33_;
  assign new_n4836 = ~new_n522 & new_n4835;
  assign new_n4837 = ~new_n4831 & ~new_n4833;
  assign new_n4838 = ~new_n4834 & ~new_n4836;
  assign poutreg_new_33_ = ~new_n4837 | ~new_n4838;
  assign new_n4840 = poutreg_40_ & ~pcount_0_;
  assign new_n4841 = ~new_n522 & new_n4840;
  assign new_n4842 = pcount_0_ & poutreg_48_;
  assign new_n4843 = ~new_n522 & new_n4842;
  assign new_n4844 = pdata_34_ & new_n522;
  assign new_n4845 = ~new_n4841 & ~new_n4843;
  assign poutreg_new_40_ = new_n4844 | ~new_n4845;
  assign new_n4847 = new_n522 & new_n4569;
  assign new_n4848 = new_n522 & new_n4571;
  assign new_n4849 = ~pcount_0_ & poutreg_59_;
  assign new_n4850 = ~new_n522 & new_n4849;
  assign new_n4851 = ~new_n4847 & ~new_n4848;
  assign poutreg_new_59_ = new_n4850 | ~new_n4851;
  assign new_n4853 = pencrypt_mode_0_ & new_n2870;
  assign new_n4854 = ~new_n529 & new_n4853;
  assign new_n4855 = ~preset_0_ & new_n4854;
  assign new_n4856 = ~pencrypt_mode_0_ & new_n3805;
  assign new_n4857 = ~new_n529 & new_n4856;
  assign new_n4858 = ~preset_0_ & new_n4857;
  assign new_n4859 = pencrypt_mode_0_ & new_n2172;
  assign new_n4860 = ~new_n529 & new_n4859;
  assign new_n4861 = ~preset_0_ & new_n4860;
  assign new_n4862 = ~pencrypt_mode_0_ & new_n4156;
  assign new_n4863 = ~new_n529 & new_n4862;
  assign new_n4864 = ~preset_0_ & new_n4863;
  assign new_n4865 = pc_20_ & ~preset_0_;
  assign new_n4866 = ~new_n512 & new_n4865;
  assign new_n4867 = ~new_n529 & new_n4866;
  assign new_n4868 = pinreg_10_ & new_n582;
  assign new_n4869 = new_n529 & new_n4868;
  assign new_n4870 = pinreg_18_ & new_n554;
  assign new_n4871 = new_n529 & new_n4870;
  assign new_n4872 = ~new_n4867 & ~new_n4869;
  assign new_n4873 = ~new_n4871 & new_n4872;
  assign new_n4874 = ~new_n4855 & ~new_n4858;
  assign new_n4875 = ~new_n4861 & ~new_n4864;
  assign new_n4876 = new_n4874 & new_n4875;
  assign pc_new_20_ = ~new_n4873 | ~new_n4876;
  assign new_n4878 = pencrypt_mode_0_ & new_n2911;
  assign new_n4879 = ~new_n529 & new_n4878;
  assign new_n4880 = ~preset_0_ & new_n4879;
  assign new_n4881 = ~pencrypt_mode_0_ & new_n819;
  assign new_n4882 = ~new_n529 & new_n4881;
  assign new_n4883 = ~preset_0_ & new_n4882;
  assign new_n4884 = pencrypt_mode_0_ & new_n2214;
  assign new_n4885 = ~new_n529 & new_n4884;
  assign new_n4886 = ~preset_0_ & new_n4885;
  assign new_n4887 = pd_9_ & new_n530;
  assign new_n4888 = ~pencrypt_mode_0_ & new_n4887;
  assign new_n4889 = ~new_n529 & new_n4888;
  assign new_n4890 = ~preset_0_ & new_n4889;
  assign new_n4891 = pd_10_ & ~preset_0_;
  assign new_n4892 = ~new_n512 & new_n4891;
  assign new_n4893 = ~new_n529 & new_n4892;
  assign new_n4894 = pinreg_29_ & new_n582;
  assign new_n4895 = new_n529 & new_n4894;
  assign new_n4896 = pinreg_37_ & new_n554;
  assign new_n4897 = new_n529 & new_n4896;
  assign new_n4898 = ~new_n4893 & ~new_n4895;
  assign new_n4899 = ~new_n4897 & new_n4898;
  assign new_n4900 = ~new_n4880 & ~new_n4883;
  assign new_n4901 = ~new_n4886 & ~new_n4890;
  assign new_n4902 = new_n4900 & new_n4901;
  assign pd_new_10_ = ~new_n4899 | ~new_n4902;
  assign new_n4904 = ~new_n522 & new_n3562;
  assign new_n4905 = ~new_n522 & new_n3558;
  assign new_n4906 = pinreg_26_ & new_n522;
  assign new_n4907 = ~new_n4904 & ~new_n4905;
  assign pdata_new_43_ = new_n4906 | ~new_n4907;
  assign new_n4909 = ~new_n522 & new_n3782;
  assign new_n4910 = ~new_n522 & new_n3778;
  assign new_n4911 = pinreg_20_ & new_n522;
  assign new_n4912 = ~new_n4909 & ~new_n4910;
  assign pdata_new_52_ = new_n4911 | ~new_n4912;
  assign new_n4914 = ~pcount_0_ & pinreg_20_;
  assign new_n4915 = ~new_n522 & new_n4914;
  assign new_n4916 = pcount_0_ & pinreg_12_;
  assign new_n4917 = ~new_n522 & new_n4916;
  assign pinreg_new_20_ = new_n4915 | new_n4917;
  assign new_n4919 = ~pcount_0_ & pinreg_31_;
  assign new_n4920 = ~new_n522 & new_n4919;
  assign new_n4921 = pcount_0_ & pinreg_23_;
  assign new_n4922 = ~new_n522 & new_n4921;
  assign pinreg_new_31_ = new_n4920 | new_n4922;
  assign new_n4924 = new_n522 & new_n4464;
  assign new_n4925 = pcount_0_ & poutreg_31_;
  assign new_n4926 = ~new_n522 & new_n4925;
  assign new_n4927 = new_n522 & new_n4462;
  assign new_n4928 = ~pcount_0_ & poutreg_23_;
  assign new_n4929 = ~new_n522 & new_n4928;
  assign new_n4930 = ~new_n4924 & ~new_n4926;
  assign new_n4931 = ~new_n4927 & ~new_n4929;
  assign poutreg_new_23_ = ~new_n4930 | ~new_n4931;
  assign new_n4933 = ~pcount_0_ & poutreg_32_;
  assign new_n4934 = ~new_n522 & new_n4933;
  assign new_n4935 = poutreg_40_ & pcount_0_;
  assign new_n4936 = ~new_n522 & new_n4935;
  assign new_n4937 = pdata_35_ & new_n522;
  assign new_n4938 = ~new_n4934 & ~new_n4936;
  assign poutreg_new_32_ = new_n4937 | ~new_n4938;
  assign new_n4940 = pencrypt_mode_0_ & new_n3334;
  assign new_n4941 = ~new_n529 & new_n4940;
  assign new_n4942 = ~preset_0_ & new_n4941;
  assign new_n4943 = ~pencrypt_mode_0_ & new_n536;
  assign new_n4944 = ~new_n529 & new_n4943;
  assign new_n4945 = ~preset_0_ & new_n4944;
  assign new_n4946 = pencrypt_mode_0_ & new_n2447;
  assign new_n4947 = ~new_n529 & new_n4946;
  assign new_n4948 = ~preset_0_ & new_n4947;
  assign new_n4949 = pc_9_ & new_n530;
  assign new_n4950 = ~pencrypt_mode_0_ & new_n4949;
  assign new_n4951 = ~new_n529 & new_n4950;
  assign new_n4952 = ~preset_0_ & new_n4951;
  assign new_n4953 = ~preset_0_ & pc_10_;
  assign new_n4954 = ~new_n512 & new_n4953;
  assign new_n4955 = ~new_n529 & new_n4954;
  assign new_n4956 = pinreg_25_ & new_n582;
  assign new_n4957 = new_n529 & new_n4956;
  assign new_n4958 = pinreg_33_ & new_n554;
  assign new_n4959 = new_n529 & new_n4958;
  assign new_n4960 = ~new_n4955 & ~new_n4957;
  assign new_n4961 = ~new_n4959 & new_n4960;
  assign new_n4962 = ~new_n4942 & ~new_n4945;
  assign new_n4963 = ~new_n4948 & ~new_n4952;
  assign new_n4964 = new_n4962 & new_n4963;
  assign pc_new_10_ = ~new_n4961 | ~new_n4964;
  assign new_n4966 = ~new_n522 & new_n3228;
  assign new_n4967 = ~new_n522 & new_n3224;
  assign new_n4968 = pinreg_18_ & new_n522;
  assign new_n4969 = ~new_n4966 & ~new_n4967;
  assign pdata_new_44_ = new_n4968 | ~new_n4969;
  assign new_n4971 = ~new_n522 & new_n2828;
  assign new_n4972 = ~new_n522 & new_n2824;
  assign new_n4973 = pinreg_28_ & new_n522;
  assign new_n4974 = ~new_n4971 & ~new_n4972;
  assign pdata_new_51_ = new_n4973 | ~new_n4974;
  assign new_n4976 = ~pcount_0_ & pinreg_21_;
  assign new_n4977 = ~new_n522 & new_n4976;
  assign new_n4978 = pcount_0_ & pinreg_13_;
  assign new_n4979 = ~new_n522 & new_n4978;
  assign pinreg_new_21_ = new_n4977 | new_n4979;
  assign new_n4981 = ~pcount_0_ & pinreg_30_;
  assign new_n4982 = ~new_n522 & new_n4981;
  assign new_n4983 = pcount_0_ & pinreg_22_;
  assign new_n4984 = ~new_n522 & new_n4983;
  assign pinreg_new_30_ = new_n4982 | new_n4984;
  assign new_n4986 = ~pcount_0_ & poutreg_24_;
  assign new_n4987 = ~new_n522 & new_n4986;
  assign new_n4988 = pcount_0_ & poutreg_32_;
  assign new_n4989 = ~new_n522 & new_n4988;
  assign new_n4990 = pdata_36_ & new_n522;
  assign new_n4991 = ~new_n4987 & ~new_n4989;
  assign poutreg_new_24_ = new_n4990 | ~new_n4991;
  assign new_n4993 = new_n522 & new_n4809;
  assign new_n4994 = pcount_0_ & poutreg_39_;
  assign new_n4995 = ~new_n522 & new_n4994;
  assign new_n4996 = new_n522 & new_n4807;
  assign new_n4997 = ~pcount_0_ & poutreg_31_;
  assign new_n4998 = ~new_n522 & new_n4997;
  assign new_n4999 = ~new_n4993 & ~new_n4995;
  assign new_n5000 = ~new_n4996 & ~new_n4998;
  assign poutreg_new_31_ = ~new_n4999 | ~new_n5000;
  assign new_n5002 = ~new_n522 & new_n4627;
  assign new_n5003 = ~new_n522 & new_n4629;
  assign new_n5004 = pinreg_48_ & new_n522;
  assign new_n5005 = ~new_n5002 & ~new_n5003;
  assign pdata_new_32_ = new_n5004 | ~new_n5005;
  assign new_n5007 = pcount_0_ & pinreg_3_;
  assign new_n5008 = ~new_n522 & new_n5007;
  assign new_n5009 = ~pcount_0_ & pinreg_11_;
  assign new_n5010 = ~new_n522 & new_n5009;
  assign pinreg_new_11_ = new_n5008 | new_n5010;
  assign new_n5012 = ~pcount_0_ & poutreg_12_;
  assign new_n5013 = ~new_n522 & new_n5012;
  assign new_n5014 = pcount_0_ & poutreg_20_;
  assign new_n5015 = ~new_n522 & new_n5014;
  assign new_n5016 = pdata_54_ & new_n522;
  assign new_n5017 = ~new_n5013 & ~new_n5015;
  assign poutreg_new_12_ = new_n5016 | ~new_n5017;
  assign new_n5019 = pinreg_21_ & new_n522;
  assign new_n5020 = pdata_52_ & ~new_n522;
  assign pdata_new_20_ = new_n5019 | new_n5020;
  assign new_n5022 = pdata_in_7_ & new_n522;
  assign new_n5023 = pdata_63_ & ~new_n522;
  assign pdata_new_31_ = new_n5022 | new_n5023;
  assign new_n5025 = pcount_0_ & pinreg_2_;
  assign new_n5026 = ~new_n522 & new_n5025;
  assign new_n5027 = ~pcount_0_ & pinreg_10_;
  assign new_n5028 = ~new_n522 & new_n5027;
  assign pinreg_new_10_ = new_n5026 | new_n5028;
  assign new_n5030 = new_n522 & new_n2591;
  assign new_n5031 = pcount_0_ & poutreg_19_;
  assign new_n5032 = ~new_n522 & new_n5031;
  assign new_n5033 = new_n522 & new_n2589;
  assign new_n5034 = ~pcount_0_ & poutreg_11_;
  assign new_n5035 = ~new_n522 & new_n5034;
  assign new_n5036 = ~new_n5030 & ~new_n5032;
  assign new_n5037 = ~new_n5033 & ~new_n5035;
  assign poutreg_new_11_ = ~new_n5036 | ~new_n5037;
  assign new_n5039 = ~new_n522 & new_n4518;
  assign new_n5040 = ~new_n522 & new_n4514;
  assign new_n5041 = pinreg_32_ & new_n522;
  assign new_n5042 = ~new_n5039 & ~new_n5040;
  assign pdata_new_34_ = new_n5041 | ~new_n5042;
  assign new_n5044 = ~pcount_0_ & poutreg_14_;
  assign new_n5045 = ~new_n522 & new_n5044;
  assign new_n5046 = pcount_0_ & poutreg_22_;
  assign new_n5047 = ~new_n522 & new_n5046;
  assign new_n5048 = pdata_62_ & new_n522;
  assign new_n5049 = ~new_n5045 & ~new_n5047;
  assign poutreg_new_14_ = new_n5048 | ~new_n5049;
  assign new_n5051 = pinreg_29_ & new_n522;
  assign new_n5052 = pdata_51_ & ~new_n522;
  assign pdata_new_19_ = new_n5051 | new_n5052;
  assign new_n5054 = ~new_n522 & new_n3297;
  assign new_n5055 = ~new_n522 & new_n3293;
  assign new_n5056 = pinreg_40_ & new_n522;
  assign new_n5057 = ~new_n5054 & ~new_n5055;
  assign pdata_new_33_ = new_n5056 | ~new_n5057;
  assign new_n5059 = new_n522 & new_n4675;
  assign new_n5060 = pcount_0_ & poutreg_21_;
  assign new_n5061 = ~new_n522 & new_n5060;
  assign new_n5062 = new_n522 & new_n4673;
  assign new_n5063 = ~pcount_0_ & poutreg_13_;
  assign new_n5064 = ~new_n522 & new_n5063;
  assign new_n5065 = ~new_n5059 & ~new_n5061;
  assign new_n5066 = ~new_n5062 & ~new_n5064;
  assign poutreg_new_13_ = ~new_n5065 | ~new_n5066;
  assign new_n5068 = pencrypt_mode_0_ & new_n3377;
  assign new_n5069 = ~new_n529 & new_n5068;
  assign new_n5070 = ~preset_0_ & new_n5069;
  assign new_n5071 = ~pencrypt_mode_0_ & new_n593;
  assign new_n5072 = ~new_n529 & new_n5071;
  assign new_n5073 = ~preset_0_ & new_n5072;
  assign new_n5074 = pencrypt_mode_0_ & new_n2504;
  assign new_n5075 = ~new_n529 & new_n5074;
  assign new_n5076 = ~preset_0_ & new_n5075;
  assign new_n5077 = pd_8_ & new_n530;
  assign new_n5078 = ~pencrypt_mode_0_ & new_n5077;
  assign new_n5079 = ~new_n529 & new_n5078;
  assign new_n5080 = ~preset_0_ & new_n5079;
  assign new_n5081 = ~preset_0_ & pd_9_;
  assign new_n5082 = ~new_n512 & new_n5081;
  assign new_n5083 = ~new_n529 & new_n5082;
  assign new_n5084 = pinreg_37_ & new_n582;
  assign new_n5085 = new_n529 & new_n5084;
  assign new_n5086 = pinreg_45_ & new_n554;
  assign new_n5087 = new_n529 & new_n5086;
  assign new_n5088 = ~new_n5083 & ~new_n5085;
  assign new_n5089 = ~new_n5087 & new_n5088;
  assign new_n5090 = ~new_n5070 & ~new_n5073;
  assign new_n5091 = ~new_n5076 & ~new_n5080;
  assign new_n5092 = new_n5090 & new_n5091;
  assign pd_new_9_ = ~new_n5089 | ~new_n5092;
  assign new_n5094 = pinreg_37_ & new_n522;
  assign new_n5095 = pdata_50_ & ~new_n522;
  assign pdata_new_18_ = new_n5094 | new_n5095;
  assign new_n5097 = pdata_in_5_ & new_n522;
  assign new_n5098 = pdata_55_ & ~new_n522;
  assign pdata_new_23_ = new_n5097 | new_n5098;
  assign new_n5100 = pinreg_45_ & new_n522;
  assign new_n5101 = pdata_49_ & ~new_n522;
  assign pdata_new_17_ = new_n5100 | new_n5101;
  assign new_n5103 = pinreg_55_ & new_n522;
  assign new_n5104 = pdata_56_ & ~new_n522;
  assign pdata_new_24_ = new_n5103 | new_n5104;
  assign new_n5106 = ~pcount_0_ & pinreg_9_;
  assign new_n5107 = ~new_n522 & new_n5106;
  assign new_n5108 = pinreg_1_ & pcount_0_;
  assign new_n5109 = ~new_n522 & new_n5108;
  assign pinreg_new_9_ = new_n5107 | new_n5109;
  assign new_n5111 = pencrypt_mode_0_ & new_n2439;
  assign new_n5112 = ~new_n529 & new_n5111;
  assign new_n5113 = ~preset_0_ & new_n5112;
  assign new_n5114 = ~pencrypt_mode_0_ & new_n1095;
  assign new_n5115 = ~new_n529 & new_n5114;
  assign new_n5116 = ~preset_0_ & new_n5115;
  assign new_n5117 = pencrypt_mode_0_ & new_n4949;
  assign new_n5118 = ~new_n529 & new_n5117;
  assign new_n5119 = ~preset_0_ & new_n5118;
  assign new_n5120 = ~pencrypt_mode_0_ & new_n543;
  assign new_n5121 = ~new_n529 & new_n5120;
  assign new_n5122 = ~preset_0_ & new_n5121;
  assign new_n5123 = ~preset_0_ & pc_8_;
  assign new_n5124 = ~new_n512 & new_n5123;
  assign new_n5125 = ~new_n529 & new_n5124;
  assign new_n5126 = pinreg_41_ & new_n582;
  assign new_n5127 = new_n529 & new_n5126;
  assign new_n5128 = pinreg_49_ & new_n554;
  assign new_n5129 = new_n529 & new_n5128;
  assign new_n5130 = ~new_n5125 & ~new_n5127;
  assign new_n5131 = ~new_n5129 & new_n5130;
  assign new_n5132 = ~new_n5113 & ~new_n5116;
  assign new_n5133 = ~new_n5119 & ~new_n5122;
  assign new_n5134 = new_n5132 & new_n5133;
  assign pc_new_8_ = ~new_n5131 | ~new_n5134;
  assign new_n5136 = ~pencrypt_mode_0_ & new_n601;
  assign new_n5137 = ~new_n529 & new_n5136;
  assign new_n5138 = ~preset_0_ & new_n5137;
  assign new_n5139 = pencrypt_mode_0_ & new_n2496;
  assign new_n5140 = ~new_n529 & new_n5139;
  assign new_n5141 = ~preset_0_ & new_n5140;
  assign new_n5142 = ~preset_0_ & pd_7_;
  assign new_n5143 = ~new_n512 & new_n5142;
  assign new_n5144 = ~new_n529 & new_n5143;
  assign new_n5145 = pencrypt_mode_0_ & new_n5077;
  assign new_n5146 = ~new_n529 & new_n5145;
  assign new_n5147 = ~preset_0_ & new_n5146;
  assign new_n5148 = ~pencrypt_0_ & new_n830;
  assign new_n5149 = new_n529 & new_n5148;
  assign new_n5150 = ~pencrypt_mode_0_ & new_n1123;
  assign new_n5151 = ~new_n529 & new_n5150;
  assign new_n5152 = ~preset_0_ & new_n5151;
  assign new_n5153 = pinreg_53_ & new_n582;
  assign new_n5154 = new_n529 & new_n5153;
  assign new_n5155 = ~new_n5149 & ~new_n5152;
  assign new_n5156 = ~new_n5154 & new_n5155;
  assign new_n5157 = ~new_n5138 & ~new_n5141;
  assign new_n5158 = ~new_n5144 & ~new_n5147;
  assign new_n5159 = new_n5157 & new_n5158;
  assign pd_new_7_ = ~new_n5156 | ~new_n5159;
  assign new_n5161 = pinreg_53_ & new_n522;
  assign new_n5162 = pdata_48_ & ~new_n522;
  assign pdata_new_16_ = new_n5161 | new_n5162;
  assign new_n5164 = pinreg_13_ & new_n522;
  assign new_n5165 = pdata_53_ & ~new_n522;
  assign pdata_new_21_ = new_n5164 | new_n5165;
  assign new_n5167 = pinreg_7_ & new_n522;
  assign new_n5168 = pdata_62_ & ~new_n522;
  assign pdata_new_30_ = new_n5167 | new_n5168;
  assign new_n5170 = ~pcount_0_ & poutreg_10_;
  assign new_n5171 = ~new_n522 & new_n5170;
  assign new_n5172 = pcount_0_ & poutreg_18_;
  assign new_n5173 = ~new_n522 & new_n5172;
  assign new_n5174 = pdata_46_ & new_n522;
  assign new_n5175 = ~new_n5171 & ~new_n5173;
  assign poutreg_new_10_ = new_n5174 | ~new_n5175;
  assign new_n5177 = pencrypt_mode_0_ & new_n2843;
  assign new_n5178 = ~new_n529 & new_n5177;
  assign new_n5179 = ~preset_0_ & new_n5178;
  assign new_n5180 = ~pencrypt_mode_0_ & new_n1229;
  assign new_n5181 = ~new_n529 & new_n5180;
  assign new_n5182 = ~preset_0_ & new_n5181;
  assign new_n5183 = pencrypt_mode_0_ & new_n2155;
  assign new_n5184 = ~new_n529 & new_n5183;
  assign new_n5185 = ~preset_0_ & new_n5184;
  assign new_n5186 = ~pencrypt_mode_0_ & new_n797;
  assign new_n5187 = ~new_n529 & new_n5186;
  assign new_n5188 = ~preset_0_ & new_n5187;
  assign new_n5189 = ~preset_0_ & pc_9_;
  assign new_n5190 = ~new_n512 & new_n5189;
  assign new_n5191 = ~new_n529 & new_n5190;
  assign new_n5192 = pinreg_33_ & new_n582;
  assign new_n5193 = new_n529 & new_n5192;
  assign new_n5194 = pinreg_41_ & new_n554;
  assign new_n5195 = new_n529 & new_n5194;
  assign new_n5196 = ~new_n5191 & ~new_n5193;
  assign new_n5197 = ~new_n5195 & new_n5196;
  assign new_n5198 = ~new_n5179 & ~new_n5182;
  assign new_n5199 = ~new_n5185 & ~new_n5188;
  assign new_n5200 = new_n5198 & new_n5199;
  assign pc_new_9_ = ~new_n5197 | ~new_n5200;
  assign new_n5202 = pencrypt_mode_0_ & new_n2206;
  assign new_n5203 = ~new_n529 & new_n5202;
  assign new_n5204 = ~preset_0_ & new_n5203;
  assign new_n5205 = ~pencrypt_mode_0_ & new_n1257;
  assign new_n5206 = ~new_n529 & new_n5205;
  assign new_n5207 = ~preset_0_ & new_n5206;
  assign new_n5208 = pencrypt_mode_0_ & new_n4887;
  assign new_n5209 = ~new_n529 & new_n5208;
  assign new_n5210 = ~preset_0_ & new_n5209;
  assign new_n5211 = ~pencrypt_mode_0_ & new_n826;
  assign new_n5212 = ~new_n529 & new_n5211;
  assign new_n5213 = ~preset_0_ & new_n5212;
  assign new_n5214 = ~preset_0_ & pd_8_;
  assign new_n5215 = ~new_n512 & new_n5214;
  assign new_n5216 = ~new_n529 & new_n5215;
  assign new_n5217 = pinreg_45_ & new_n582;
  assign new_n5218 = new_n529 & new_n5217;
  assign new_n5219 = pinreg_53_ & new_n554;
  assign new_n5220 = new_n529 & new_n5219;
  assign new_n5221 = ~new_n5216 & ~new_n5218;
  assign new_n5222 = ~new_n5220 & new_n5221;
  assign new_n5223 = ~new_n5204 & ~new_n5207;
  assign new_n5224 = ~new_n5210 & ~new_n5213;
  assign new_n5225 = new_n5223 & new_n5224;
  assign pd_new_8_ = ~new_n5222 | ~new_n5225;
  assign new_n5227 = pdata_in_3_ & new_n522;
  assign new_n5228 = pdata_47_ & ~new_n522;
  assign pdata_new_15_ = new_n5227 | new_n5228;
  assign new_n5230 = pinreg_5_ & new_n522;
  assign new_n5231 = pdata_54_ & ~new_n522;
  assign pdata_new_22_ = new_n5230 | new_n5231;
endmodule


