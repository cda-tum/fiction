// Benchmark "c1196" written by ABC on Mon Sep 23 09:57:39 2019

module c1196 ( 
    G0, G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46,
    G546, G539, G550, G551, G552, G547, G548, G549, G530, G542, G532, G535,
    G537, G502, G503, G504, G505, G506, G507, G508, G509, G510, G511, G512,
    G513, G514, G515, G516, G517, G518, G519  );
  input  G0, G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G29,
    G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43,
    G44, G45, G46;
  output G546, G539, G550, G551, G552, G547, G548, G549, G530, G542, G532,
    G535, G537, G502, G503, G504, G505, G506, G507, G508, G509, G510, G511,
    G512, G513, G514, G515, G516, G517, G518, G519;
  wire new_G520_, new_G521_, new_G522_, new_G524_, new_II156_, new_G334_,
    new_G527_, new_G528_, new_G529_, new_G531_, new_G533_, new_G536_,
    new_G538_, new_G540_, new_G541_, new_G543_, new_G476_, new_G484_,
    new_G125_, new_G140_, new_G132_, new_G70_, new_G67_, new_G99_,
    new_G475_, new_G59_, new_G228_, new_G272_, new_G98_, new_G135_,
    new_II218_, new_G333_, new_G55_, new_G165_, new_G72_, new_G236_,
    new_G275_, new_II249_, new_G370_, new_G75_, new_G490_, new_G482_,
    new_G153_, new_G192_, new_G123_, new_II272_, new_G458_, new_II276_,
    new_G332_, new_II280_, new_G309_, new_II287_, new_G347_, new_G498_,
    new_G78_, new_II295_, new_G459_, new_G199_, new_G90_, new_G221_,
    new_G223_, new_II316_, new_G369_, new_G234_, new_II327_, new_G435_,
    new_II330_, new_G441_, new_G50_, new_G130_, new_G501_, new_G477_,
    new_G485_, new_II352_, new_G299_, new_G497_, new_II371_, new_G335_,
    new_II374_, new_G456_, new_G87_, new_II386_, new_G414_, new_G486_,
    new_G231_, new_G160_, new_G265_, new_G64_, new_G180_, new_G107_,
    new_G207_, new_G167_, new_G124_, new_G203_, new_G489_, new_G495_,
    new_G177_, new_G212_, new_II493_, new_G404_, new_II502_, new_G468_,
    new_G173_, new_G487_, new_II529_, new_G149_, new_II536_, new_G446_,
    new_G494_, new_G500_, new_G214_, new_G492_, new_G483_, new_G282_,
    new_II573_, new_G403_, new_II576_, new_G447_, new_G479_, new_G491_,
    new_G554_, new_G170_, new_G172_, new_G525_, new_G493_, new_G545_,
    new_G488_, new_G499_, new_II624_, new_G303_, new_G480_, new_II631_,
    new_G336_, new_G496_, new_G174_, new_II662_, new_G405_, new_G478_,
    new_II692_, new_G432_, new_G359_, new_G469_, new_G461_, new_G431_,
    new_G362_, new_G81_, new_G348_, new_G352_, new_G379_, new_G385_,
    new_G376_, new_G387_, new_G462_, new_G436_, new_G363_, new_G410_,
    new_G399_, new_G437_, new_G307_, new_G306_, new_G283_, new_G339_,
    new_G472_, new_G351_, new_G440_, new_G382_, new_G386_, new_G321_,
    new_G378_, new_G471_, new_G377_, new_G358_, new_G400_, new_G308_,
    new_G411_, new_G413_, new_G434_, new_G373_, new_G357_, new_G444_,
    new_G361_, new_G346_, new_G457_, new_G364_, new_G445_, new_G412_,
    new_G371_, new_G353_, new_G388_, new_G473_, new_G331_, new_G429_,
    new_G380_, new_G360_, new_G338_, new_G337_, new_G340_, new_G322_,
    new_G330_, new_G430_, new_G344_, new_G428_, new_G349_, new_G460_,
    new_G463_, new_G393_, new_G470_, new_G341_, new_G342_, new_G324_,
    new_G323_, new_G354_, new_G312_, new_G315_, new_G474_, new_G343_,
    new_G304_, new_G398_, new_G365_, new_G417_, new_G290_, new_G327_,
    new_G367_, new_G397_, new_G451_, new_G406_, new_G418_, new_G453_,
    new_G289_, new_G311_, new_G402_, new_G433_, new_G449_, new_G452_,
    new_G329_, new_G291_, new_G328_, new_G366_, new_G372_, new_G383_,
    new_G392_, new_G396_, new_G401_, new_G422_, new_G415_, new_G425_,
    new_G438_, new_G424_, new_G439_, new_G317_, new_G426_, new_G443_,
    new_G416_, new_G427_, new_G442_, new_G423_, new_G448_, new_G419_,
    new_G193_, new_G394_, new_G407_, new_G314_, new_G395_, new_G288_,
    new_G302_, new_G224_, new_G355_, new_G316_, new_G350_, new_G368_,
    new_G381_, new_G384_, new_G389_, new_G374_, new_G286_, new_G293_,
    new_G375_, new_G356_, new_G313_, new_G420_, new_G421_, new_G320_,
    new_G310_, new_G408_, new_G305_, new_G409_, new_G296_, new_G325_,
    new_G464_, new_G391_, new_G292_, new_G345_, new_G465_, new_G454_,
    new_G269_, new_G287_, new_G318_, new_G326_, new_G390_, new_G298_,
    new_G300_, new_G261_, new_G301_, new_G92_, new_G47_, new_G114_,
    new_G297_, new_G93_, new_G106_, new_G110_, new_G455_, new_G152_,
    new_G60_, new_G133_, new_G105_, new_G108_, new_G115_, new_G126_,
    new_G79_, new_G319_, new_G131_, new_G118_, new_G73_, new_G91_,
    new_G137_, new_G242_, new_G147_, new_G284_, new_G294_, new_G553_,
    new_G141_, new_G142_, new_G88_, new_G544_, new_G285_, new_G295_,
    new_G450_, new_G150_, new_G146_, new_G244_, new_G61_, new_G95_,
    new_G121_, new_G279_, new_G128_, new_G145_, new_G139_, new_G57_,
    new_G58_, new_G76_, new_G101_, new_G117_, new_G271_, new_G97_,
    new_G134_, new_G54_, new_G116_, new_G71_, new_G274_, new_G74_,
    new_G112_, new_G245_, new_G122_, new_G238_, new_G129_, new_G240_,
    new_G252_, new_G77_, new_G103_, new_G200_, new_G248_, new_G89_,
    new_G222_, new_G239_, new_G235_, new_G220_, new_G49_, new_G251_,
    new_G276_, new_G263_, new_G226_, new_G210_, new_G66_, new_G233_,
    new_G104_, new_G86_, new_G219_, new_G68_, new_G232_, new_G136_,
    new_G161_, new_G100_, new_G85_, new_G243_, new_G63_, new_G237_,
    new_G56_, new_G83_, new_G96_, new_G278_, new_G255_, new_G69_,
    new_G181_, new_G277_, new_G151_, new_G48_, new_G264_, new_G208_,
    new_G168_, new_G84_, new_G258_, new_G166_, new_G259_, new_G217_,
    new_G257_, new_G260_, new_G266_, new_G262_, new_G138_, new_G256_,
    new_G82_, new_G109_, new_G206_, new_G204_, new_G53_, new_G273_,
    new_G267_, new_G113_, new_G143_, new_G213_, new_G51_, new_G102_,
    new_G52_, new_G80_, new_G270_, new_G94_, new_G249_, new_G268_,
    new_G111_, new_G534_, new_G253_, new_G148_, new_G254_, new_G127_,
    new_G215_, new_G62_, new_G523_, new_G144_, new_G250_, new_G281_,
    new_G171_, new_G526_, new_G280_, new_G246_, new_G119_, new_G120_,
    new_G185_, new_G159_, new_G163_, new_G216_, new_G169_, new_G225_,
    new_G190_, new_G241_, new_G198_, new_G178_, new_G229_, new_G209_,
    new_G195_, new_G189_, new_G201_, new_G164_, new_G211_, new_G156_,
    new_G205_, new_G227_, new_G230_, new_G191_, new_G196_, new_G197_,
    new_G202_, new_G218_, new_G183_, new_G182_, new_G176_, new_G175_,
    new_G187_, new_G158_, new_G194_, new_G157_, new_G186_, new_G247_,
    new_G179_, new_G188_, new_G154_, new_G184_, new_G155_, new_G162_;
  assign new_G520_ = ~G0;
  assign new_G521_ = ~G1;
  assign new_G522_ = ~G2;
  assign new_G524_ = ~G3;
  assign new_II156_ = ~G4;
  assign new_G334_ = ~new_II156_;
  assign new_G527_ = ~G4;
  assign new_G528_ = ~G5;
  assign new_G529_ = ~G6;
  assign new_G531_ = ~G7;
  assign new_G533_ = ~G8;
  assign new_G536_ = ~G9;
  assign new_G538_ = ~G10;
  assign new_G540_ = ~G11;
  assign new_G541_ = ~G12;
  assign new_G543_ = ~G13;
  assign new_G476_ = ~G30;
  assign new_G484_ = ~G30;
  assign new_G125_ = ~G40;
  assign new_G140_ = ~G33;
  assign G546 = ~G41;
  assign new_G132_ = ~G42;
  assign new_G70_ = ~G43;
  assign new_G67_ = ~G44;
  assign new_G99_ = ~G29;
  assign new_G475_ = ~new_G57_;
  assign new_G59_ = ~new_G58_;
  assign new_G228_ = ~new_G524_;
  assign new_G272_ = ~new_G271_;
  assign new_G98_ = ~new_G97_;
  assign new_G135_ = ~new_G134_;
  assign new_II218_ = ~new_G528_;
  assign new_G333_ = ~new_II218_;
  assign new_G55_ = ~new_G54_;
  assign new_G165_ = ~new_G529_;
  assign new_G72_ = ~new_G71_;
  assign new_G236_ = ~new_G274_;
  assign new_G275_ = ~new_G274_;
  assign new_II249_ = ~new_G538_;
  assign new_G370_ = ~new_II249_;
  assign new_G75_ = ~new_G74_;
  assign new_G490_ = ~new_G190_;
  assign new_G482_ = ~new_G241_;
  assign new_G153_ = ~new_G522_;
  assign new_G192_ = ~new_G193_;
  assign new_G123_ = ~new_G122_;
  assign new_II272_ = ~new_G209_;
  assign new_G458_ = ~new_II272_;
  assign new_II276_ = ~new_G238_;
  assign new_G332_ = ~new_II276_;
  assign new_II280_ = ~new_G272_;
  assign new_G309_ = ~new_II280_;
  assign new_II287_ = ~new_G135_;
  assign new_G347_ = ~new_II287_;
  assign new_G498_ = ~new_G195_;
  assign new_G78_ = ~new_G77_;
  assign new_II295_ = ~new_G198_;
  assign new_G459_ = ~new_II295_;
  assign new_G199_ = ~new_G200_;
  assign new_G90_ = ~new_G89_;
  assign new_G221_ = ~new_G222_;
  assign new_G223_ = ~new_G224_;
  assign new_II316_ = ~new_G239_;
  assign new_G369_ = ~new_II316_;
  assign new_G234_ = ~new_G235_;
  assign new_II327_ = ~new_G135_;
  assign new_G435_ = ~new_II327_;
  assign new_II330_ = ~new_G236_;
  assign new_G441_ = ~new_II330_;
  assign new_G50_ = ~new_G49_;
  assign new_G130_ = ~G9;
  assign new_G501_ = ~new_G156_;
  assign new_G477_ = ~new_G276_;
  assign new_G485_ = ~new_G276_;
  assign new_II352_ = ~new_G77_;
  assign new_G299_ = ~new_II352_;
  assign new_G497_ = ~new_G205_;
  assign new_II371_ = ~G1;
  assign new_G335_ = ~new_II371_;
  assign new_II374_ = ~new_G520_;
  assign new_G456_ = ~new_II374_;
  assign new_G87_ = ~new_G86_;
  assign new_II386_ = ~new_G199_;
  assign new_G414_ = ~new_II386_;
  assign new_G486_ = ~new_G68_;
  assign new_G231_ = ~new_G232_;
  assign new_G160_ = ~new_G161_;
  assign new_G265_ = ~new_G50_;
  assign new_G64_ = ~new_G63_;
  assign new_G180_ = ~new_G181_;
  assign new_G107_ = ~new_G456_;
  assign new_G207_ = ~new_G208_;
  assign new_G167_ = ~new_G168_;
  assign new_G124_ = ~new_G206_;
  assign new_G203_ = ~new_G204_;
  assign new_G489_ = ~new_G273_;
  assign new_G495_ = ~new_G273_;
  assign new_G177_ = ~new_G357_;
  assign new_G212_ = ~new_G213_;
  assign new_II493_ = ~new_G218_;
  assign new_G404_ = ~new_II493_;
  assign new_II502_ = ~new_G124_;
  assign new_G468_ = ~new_II502_;
  assign new_G173_ = ~new_G495_;
  assign new_G487_ = ~new_G534_;
  assign new_II529_ = ~new_G468_;
  assign new_G149_ = ~new_II529_;
  assign new_II536_ = ~new_G79_;
  assign new_G446_ = ~new_II536_;
  assign new_G494_ = ~new_G173_;
  assign new_G500_ = ~new_G173_;
  assign new_G214_ = ~new_G215_;
  assign new_G492_ = ~new_G62_;
  assign new_G483_ = ~new_G182_;
  assign new_G282_ = ~new_G281_;
  assign new_II573_ = ~new_G176_;
  assign new_G403_ = ~new_II573_;
  assign new_II576_ = ~new_G175_;
  assign new_G447_ = ~new_II576_;
  assign new_G479_ = ~new_G194_;
  assign new_G491_ = ~new_G194_;
  assign new_G554_ = ~new_G553_;
  assign new_G170_ = ~new_G171_;
  assign new_G172_ = ~new_G171_;
  assign new_G525_ = ~new_G526_;
  assign new_G493_ = ~new_G544_;
  assign new_G545_ = ~new_G544_;
  assign new_G488_ = ~new_G172_;
  assign new_G499_ = ~new_G280_;
  assign new_II624_ = ~new_G120_;
  assign new_G303_ = ~new_II624_;
  assign new_G480_ = ~new_G179_;
  assign new_II631_ = ~new_G188_;
  assign new_G336_ = ~new_II631_;
  assign new_G496_ = ~new_G188_;
  assign new_G174_ = ~new_G496_;
  assign new_II662_ = ~new_G174_;
  assign new_G405_ = ~new_II662_;
  assign new_G478_ = ~new_G279_;
  assign new_II692_ = ~new_G145_;
  assign new_G432_ = ~new_II692_;
  assign new_G359_ = G6 & G31;
  assign new_G469_ = new_G163_ & G3;
  assign new_G461_ = new_G529_ & new_G531_;
  assign new_G431_ = new_G524_ & new_G67_;
  assign new_G362_ = new_G129_ & new_G77_;
  assign new_G81_ = new_G288_ & new_G240_;
  assign new_G348_ = new_G97_ & new_G55_;
  assign new_G352_ = new_G164_ & G37 & G8 & new_G135_;
  assign G511 = new_G163_ & new_G164_;
  assign new_G379_ = G9 & new_G211_;
  assign new_G385_ = new_G49_ & new_G529_ & G7;
  assign new_G376_ = new_G533_ & new_G75_;
  assign new_G387_ = new_G75_ & G6 & new_G274_;
  assign new_G462_ = new_G192_ & new_G538_;
  assign new_G436_ = new_G123_ & new_G77_;
  assign new_G363_ = new_G77_ & new_G205_;
  assign new_G410_ = G1 & new_G205_;
  assign new_G399_ = new_G520_ & G1;
  assign new_G437_ = new_G66_ & new_G229_;
  assign new_G307_ = G6 & new_G104_;
  assign new_G306_ = new_G524_ & new_G78_;
  assign new_G283_ = new_G122_ & new_G219_;
  assign new_G339_ = new_G209_ & new_G533_ & new_G199_;
  assign new_G472_ = new_G190_ & new_G136_ & G9;
  assign new_G351_ = new_G234_ & new_G221_ & new_G524_ & new_G169_;
  assign new_G440_ = G38 & new_G234_;
  assign new_G382_ = G34 & G9 & new_G100_;
  assign new_G386_ = new_G536_ & new_G85_;
  assign new_G321_ = new_G90_ & new_G50_;
  assign new_G378_ = new_G89_ & new_G50_;
  assign new_G471_ = new_G112_ & new_G191_ & new_G103_;
  assign new_G377_ = new_G90_ & new_G56_;
  assign new_G358_ = G7 & new_G83_;
  assign new_G400_ = G0 & new_G277_;
  assign new_G308_ = G5 & new_G151_;
  assign new_G411_ = new_G48_ & new_G59_;
  assign new_G413_ = new_G197_ & new_G201_;
  assign new_G434_ = new_G165_ & new_G231_;
  assign new_G373_ = G34 & new_G160_;
  assign new_G357_ = new_G265_ & new_G232_;
  assign new_G444_ = new_G211_ & new_G64_ & new_G78_;
  assign new_G361_ = G6 & new_G202_;
  assign new_G346_ = G2 & new_G82_;
  assign new_G457_ = G4 & new_G107_;
  assign new_G364_ = G2 & new_G109_;
  assign new_G445_ = new_G53_ & new_G225_;
  assign new_G412_ = G3 & new_G207_;
  assign new_G371_ = new_G267_ & new_G161_ & new_G168_;
  assign new_G353_ = new_G163_ & G11 & new_G92_;
  assign new_G388_ = G11 & new_G114_;
  assign new_G473_ = G11 & new_G143_;
  assign new_G331_ = new_G213_ & new_G257_;
  assign new_G429_ = new_G51_ & new_G225_;
  assign new_G380_ = G6 & new_G93_;
  assign new_G360_ = G8 & new_G106_;
  assign new_G338_ = new_G202_ & new_G203_;
  assign new_G337_ = new_G270_ & new_G167_;
  assign new_G340_ = G8 & new_G270_;
  assign new_G322_ = new_G196_ & new_G522_ & new_G105_;
  assign new_G330_ = new_G248_ & new_G249_;
  assign new_G430_ = new_G177_ & new_G196_;
  assign new_G344_ = new_G195_ & new_G111_ & new_G189_;
  assign new_G428_ = new_G212_ & new_G227_;
  assign new_G349_ = G6 & new_G108_;
  assign new_G460_ = new_G115_ & G2 & new_G81_;
  assign new_G463_ = new_G521_ & new_G148_;
  assign new_G393_ = new_G127_ & G34;
  assign new_G470_ = new_G528_ & new_G149_;
  assign new_G341_ = new_G531_ & new_G118_;
  assign new_G342_ = new_G73_ & new_G197_;
  assign new_G324_ = new_G522_ & new_G183_;
  assign new_G323_ = G2 & new_G144_;
  assign new_G354_ = G0 & new_G214_;
  assign new_G312_ = new_G180_ & new_G182_;
  assign new_G315_ = new_G250_ & new_G251_;
  assign new_G474_ = new_G242_ & new_G77_;
  assign new_G343_ = new_G147_ & G2 & new_G528_;
  assign new_G304_ = new_G52_ & new_G158_;
  assign new_G398_ = new_G158_ & new_G94_ & new_G156_;
  assign new_G365_ = new_G156_ & new_G282_ & new_G137_;
  assign new_G417_ = new_G70_ & G13 & new_G282_;
  assign new_G290_ = new_G157_ & new_G117_ & new_G135_;
  assign new_G327_ = new_G157_ & G4 & G39;
  assign new_G367_ = new_G126_ & new_G157_;
  assign new_G397_ = new_G157_ & new_G101_ & new_G98_;
  assign new_G451_ = new_G187_ & new_G541_ & new_G554_;
  assign new_G406_ = new_G87_ & new_G172_;
  assign new_G418_ = new_G172_ & new_G524_ & new_G60_;
  assign new_G453_ = new_G545_ & new_G186_;
  assign new_G289_ = new_G156_ & G2 & new_G119_;
  assign new_G311_ = new_G179_ & G0 & new_G178_;
  assign new_G402_ = new_G154_ & new_G183_;
  assign new_G433_ = new_G91_ & new_G154_;
  assign new_G449_ = new_G88_ & new_G154_;
  assign new_G452_ = new_G526_ & new_G184_;
  assign new_G329_ = new_G150_ & new_G156_;
  assign new_G291_ = new_G138_ & new_G155_;
  assign new_G328_ = new_G155_ & G5 & new_G102_;
  assign new_G366_ = new_G125_ & new_G155_;
  assign new_G372_ = new_G155_ & new_G116_ & new_G275_;
  assign new_G383_ = new_G131_ & new_G155_;
  assign new_G392_ = new_G132_ & new_G155_;
  assign new_G396_ = new_G155_ & new_G76_ & new_G272_;
  assign new_G401_ = new_G155_ & G2 & new_G110_;
  assign new_G422_ = new_G155_ & G0 & new_G80_;
  assign new_G415_ = new_G165_ & new_G146_ & new_G142_;
  assign new_G425_ = new_G146_ & new_G176_;
  assign new_G438_ = new_G133_ & G8 & new_G146_;
  assign new_G424_ = new_G177_ & new_G78_ & new_G174_;
  assign new_G439_ = new_G174_ & new_G175_;
  assign new_G317_ = new_G159_ & new_G245_;
  assign new_G426_ = G38 & G37 & new_G162_;
  assign new_G443_ = new_G47_ & new_G162_;
  assign new_G416_ = new_G61_ & new_G167_;
  assign new_G427_ = new_G165_ & new_G541_ & new_G95_;
  assign new_G442_ = new_G541_ & new_G121_;
  assign new_G423_ = new_G541_ & new_G128_;
  assign new_G448_ = new_G139_ & new_G153_;
  assign new_G419_ = G3 | G5;
  assign new_G193_ = G6 | G30;
  assign new_G394_ = G5 | new_G58_;
  assign new_G407_ = G6 | new_G117_;
  assign new_G314_ = new_G527_ | new_G57_;
  assign new_G395_ = G4 | new_G134_;
  assign new_G288_ = G1 | new_G528_;
  assign new_G302_ = G4 | new_G529_;
  assign new_G224_ = new_G533_ | G31;
  assign new_G355_ = G11 | new_G116_;
  assign new_G316_ = new_G531_ | new_G536_;
  assign new_G350_ = G6 | new_G536_;
  assign new_G368_ = new_G533_ | new_G536_;
  assign new_G381_ = G7 | new_G71_;
  assign new_G384_ = new_G529_ | new_G71_;
  assign new_G389_ = G9 | new_G274_;
  assign new_G374_ = new_G536_ | new_G538_;
  assign new_G286_ = G9 | new_G540_;
  assign new_G293_ = G7 | new_G540_;
  assign new_G375_ = G10 | new_G540_;
  assign new_G356_ = G6 | new_G476_;
  assign new_G313_ = new_G521_ | new_G475_;
  assign new_G420_ = new_G522_ | new_G59_;
  assign new_G421_ = new_G228_ | new_G521_ | G2;
  assign new_G320_ = new_G76_ | new_G272_;
  assign new_G310_ = new_G522_ | new_G135_;
  assign new_G408_ = new_G529_ | new_G77_;
  assign new_G305_ = new_G524_ | new_G55_;
  assign new_G409_ = new_G528_ | new_G55_;
  assign new_G296_ = new_G89_ | new_G484_;
  assign new_G325_ = new_G222_ | G7 | new_G536_;
  assign new_G464_ = new_G72_ | new_G536_;
  assign new_G391_ = new_G74_ | new_G220_;
  assign new_G292_ = new_G538_ | new_G75_;
  assign new_G345_ = new_G529_ | new_G226_;
  assign new_G465_ = new_G524_ | new_G210_;
  assign new_G454_ = new_G122_ | new_G77_;
  assign new_G269_ = new_G362_ | new_G529_;
  assign new_G287_ = new_G522_ | new_G81_;
  assign new_G318_ = new_G232_ | G6 | G8;
  assign new_G326_ = new_G533_ | new_G232_;
  assign new_G390_ = new_G89_ | new_G50_;
  assign new_G298_ = G5 | new_G497_;
  assign new_G300_ = new_G87_ | new_G97_;
  assign new_G261_ = new_G283_ | new_G528_;
  assign new_G301_ = new_G122_ | new_G486_;
  assign new_G92_ = new_G351_ | new_G352_;
  assign new_G47_ = new_G440_ | new_G441_;
  assign new_G114_ = new_G385_ | new_G386_;
  assign new_G297_ = new_G64_ | new_G274_;
  assign new_G93_ = new_G378_ | new_G376_ | new_G377_;
  assign new_G106_ = new_G358_ | new_G359_;
  assign new_G110_ = new_G399_ | new_G400_;
  assign new_G455_ = new_G78_ | new_G206_;
  assign new_G152_ = new_G308_ | new_G306_ | new_G307_;
  assign new_G60_ = new_G413_ | new_G414_;
  assign new_G133_ = new_G434_ | new_G435_;
  assign new_G105_ = new_G321_ | new_G273_;
  assign new_G108_ = new_G346_ | new_G347_;
  assign new_G115_ = new_G459_ | new_G457_ | new_G458_;
  assign new_G126_ = new_G363_ | new_G364_;
  assign new_G79_ = new_G444_ | new_G445_;
  assign new_G319_ = new_G529_ | new_G489_;
  assign new_G131_ = new_G379_ | new_G380_;
  assign new_G118_ = new_G337_ | new_G338_;
  assign new_G73_ = new_G339_ | new_G340_;
  assign new_G91_ = new_G430_ | new_G431_;
  assign new_G137_ = new_G348_ | new_G349_;
  assign new_G242_ = new_G469_ | new_G470_;
  assign new_G147_ = new_G341_ | new_G342_;
  assign new_G284_ = new_G281_ | new_G528_ | new_G272_;
  assign new_G294_ = new_G281_ | G1 | new_G117_;
  assign new_G553_ = new_G324_ | new_G322_ | new_G323_;
  assign new_G141_ = new_G353_ | new_G354_;
  assign new_G142_ = new_G403_ | new_G404_;
  assign new_G88_ = new_G446_ | new_G447_;
  assign new_G544_ = new_G343_ | new_G344_;
  assign new_G285_ = G5 | new_G479_;
  assign new_G295_ = new_G122_ | new_G491_;
  assign new_G450_ = G12 | new_G171_;
  assign new_G150_ = new_G303_ | new_G304_;
  assign new_G146_ = new_G336_ | new_G170_;
  assign G539 = new_G453_ | new_G451_ | new_G452_;
  assign new_G244_ = new_G371_ | new_G159_;
  assign G550 = new_G485_ | new_G291_ | new_G289_ | new_G290_;
  assign G551 = new_G329_ | new_G327_ | new_G328_;
  assign G552 = new_G367_ | new_G365_ | new_G366_;
  assign G547 = new_G382_ | new_G383_;
  assign G548 = new_G392_ | new_G393_;
  assign G549 = new_G477_ | new_G398_ | new_G396_ | new_G397_;
  assign G530 = new_G401_ | new_G402_;
  assign new_G61_ = new_G405_ | new_G406_;
  assign new_G95_ = new_G424_ | new_G425_;
  assign new_G121_ = new_G438_ | new_G439_;
  assign new_G279_ = new_G317_ | new_G166_;
  assign new_G128_ = new_G418_ | new_G417_ | new_G415_ | new_G416_;
  assign new_G145_ = new_G426_ | new_G427_;
  assign new_G139_ = new_G442_ | new_G443_;
  assign G532 = new_G422_ | new_G423_;
  assign G535 = new_G432_ | new_G433_;
  assign G537 = new_G448_ | new_G449_;
  assign new_G57_ = ~G0 | ~G2;
  assign new_G58_ = ~G1 | ~G3;
  assign new_G76_ = ~G0 | ~G3;
  assign new_G101_ = ~G3 | ~G4;
  assign new_G117_ = ~G2 | ~G4;
  assign new_G271_ = ~G1 | ~G4;
  assign new_G97_ = ~G2 | ~G5;
  assign new_G134_ = ~G3 | ~G5;
  assign new_G54_ = ~G4 | ~G6;
  assign new_G116_ = ~G6 | ~G9;
  assign new_G71_ = ~G8 | ~G10;
  assign new_G274_ = ~G7 | ~G10;
  assign new_G74_ = ~G9 | ~G11;
  assign new_G112_ = ~G8 | ~G31;
  assign new_G245_ = ~G8 | ~G34;
  assign new_G122_ = ~new_G522_ | ~G3;
  assign new_G238_ = ~G2 | ~new_G524_;
  assign new_G129_ = ~new_G527_ | ~G5;
  assign new_G240_ = ~G4 | ~new_G134_;
  assign new_G252_ = ~new_G216_ | ~G35 | ~G3 | ~G11;
  assign new_G77_ = ~G4 | ~new_G528_;
  assign new_G103_ = ~G30 | ~new_G529_ | ~G7;
  assign new_G200_ = ~new_G527_ | ~new_G529_;
  assign new_G248_ = ~new_G529_ | ~G36;
  assign new_G89_ = ~new_G531_ | ~G8;
  assign new_G222_ = ~new_G533_ | ~G10;
  assign new_G239_ = ~G7 | ~new_G533_;
  assign new_G235_ = ~G6 | ~new_G536_;
  assign new_G220_ = ~G7 | ~new_G71_;
  assign new_G49_ = ~G9 | ~new_G538_;
  assign new_G251_ = ~new_G543_ | ~G32;
  assign new_G276_ = ~new_G140_ | ~G3 | ~new_G543_;
  assign new_G263_ = ~G0 | ~new_G99_;
  assign new_G226_ = ~new_G527_ | ~new_G59_;
  assign new_G210_ = ~new_G520_ | ~new_G272_;
  assign new_G66_ = ~new_G129_ | ~new_G101_;
  assign new_G233_ = ~new_G522_ | ~new_G135_;
  assign new_G104_ = ~new_G240_ | ~new_G122_ | ~new_G238_;
  assign new_G86_ = ~new_G55_ | ~G3;
  assign new_G219_ = ~new_G524_ | ~new_G55_;
  assign new_G68_ = ~new_G302_ | ~new_G528_;
  assign new_G232_ = ~new_G536_ | ~new_G164_;
  assign new_G136_ = ~new_G222_ | ~new_G224_;
  assign G510 = ~new_G350_ | ~new_G235_;
  assign new_G161_ = ~new_G316_ | ~new_G72_;
  assign new_G100_ = ~new_G381_ | ~new_G220_;
  assign new_G85_ = ~new_G384_ | ~new_G239_;
  assign new_G243_ = ~G34 | ~new_G368_ | ~new_G275_;
  assign new_G63_ = ~new_G75_ | ~G8;
  assign new_G237_ = ~new_G201_ | ~G10 | ~new_G75_;
  assign G503 = ~new_G286_ | ~new_G538_;
  assign new_G56_ = ~new_G374_ | ~new_G375_;
  assign new_G83_ = ~new_G355_ | ~new_G356_;
  assign new_G96_ = ~new_G313_ | ~new_G314_;
  assign new_G278_ = ~new_G332_ | ~new_G333_;
  assign new_G255_ = ~new_G529_ | ~new_G309_ | ~G2;
  assign new_G69_ = ~new_G233_ | ~new_G419_ | ~new_G420_;
  assign G512 = ~new_G310_ | ~new_G233_;
  assign new_G181_ = ~G2 | ~new_G78_;
  assign new_G277_ = ~new_G81_ | ~new_G394_ | ~new_G395_;
  assign new_G151_ = ~new_G305_ | ~new_G200_;
  assign new_G48_ = ~new_G409_ | ~new_G407_ | ~new_G408_;
  assign new_G264_ = ~new_G227_ | ~new_G241_;
  assign new_G208_ = ~new_G68_ | ~new_G229_;
  assign new_G168_ = ~new_G75_ | ~new_G221_;
  assign new_G84_ = ~new_G369_ | ~new_G370_;
  assign new_G258_ = ~new_G223_ | ~new_G464_ | ~new_G103_;
  assign new_G166_ = ~G7 | ~new_G50_;
  assign new_G259_ = ~new_G130_ | ~new_G225_;
  assign G504 = ~new_G292_ | ~new_G293_;
  assign new_G217_ = ~new_G50_ | ~new_G230_;
  assign new_G257_ = ~new_G538_ | ~new_G230_;
  assign new_G260_ = ~new_G191_ | ~new_G528_ | ~new_G529_;
  assign new_G266_ = ~new_G524_ | ~new_G96_;
  assign new_G262_ = ~new_G527_ | ~new_G278_;
  assign new_G138_ = ~new_G465_ | ~new_G263_;
  assign new_G256_ = ~G4 | ~new_G69_;
  assign new_G82_ = ~new_G334_ | ~new_G335_;
  assign new_G109_ = ~new_G269_ | ~new_G219_;
  assign new_G206_ = ~new_G287_ | ~new_G524_;
  assign new_G204_ = ~new_G521_ | ~new_G87_;
  assign new_G53_ = ~new_G264_ | ~new_G237_;
  assign new_G273_ = ~new_G325_ | ~new_G326_;
  assign new_G267_ = ~new_G536_ | ~new_G84_;
  assign new_G113_ = ~new_G389_ | ~new_G390_;
  assign new_G143_ = ~new_G259_ | ~new_G258_ | ~new_G193_;
  assign new_G213_ = ~new_G64_ | ~new_G275_;
  assign new_G51_ = ~new_G260_ | ~new_G237_;
  assign new_G102_ = ~new_G210_ | ~new_G320_ | ~new_G266_;
  assign new_G52_ = ~new_G219_ | ~new_G298_ | ~new_G299_;
  assign new_G80_ = ~new_G256_ | ~new_G421_ | ~new_G226_;
  assign new_G270_ = ~new_G345_ | ~new_G204_;
  assign new_G94_ = ~new_G262_ | ~new_G261_ | ~new_G181_;
  assign G505 = ~new_G181_ | ~new_G300_ | ~new_G301_;
  assign new_G249_ = ~new_G201_ | ~G11 | ~new_G273_;
  assign new_G268_ = ~G11 | ~new_G113_;
  assign new_G111_ = ~new_G213_ | ~new_G217_;
  assign new_G534_ = ~new_G166_ | ~new_G296_ | ~new_G297_;
  assign new_G253_ = ~new_G87_ | ~new_G218_;
  assign new_G148_ = ~G0 | ~new_G454_ | ~new_G455_;
  assign new_G254_ = ~G1 | ~new_G152_;
  assign new_G127_ = ~new_G391_ | ~new_G268_;
  assign new_G215_ = ~new_G212_ | ~new_G135_ | ~new_G55_;
  assign new_G62_ = ~new_G534_ | ~G32;
  assign new_G523_ = ~new_G208_ | ~new_G254_ | ~new_G255_;
  assign G508 = ~new_G318_ | ~new_G319_;
  assign new_G144_ = ~new_G253_ | ~new_G215_ | ~new_G252_;
  assign new_G250_ = ~G13 | ~new_G523_;
  assign new_G281_ = ~new_G523_ | ~new_G534_;
  assign new_G171_ = ~new_G553_ | ~new_G187_;
  assign new_G526_ = ~new_G141_ | ~G1 | ~G2;
  assign new_G280_ = ~G46 | ~new_G247_;
  assign new_G246_ = ~new_G544_ | ~new_G186_;
  assign new_G119_ = ~new_G284_ | ~new_G285_;
  assign new_G120_ = ~new_G294_ | ~new_G295_;
  assign new_G185_ = ~new_G525_ | ~new_G184_;
  assign new_G159_ = ~G6 | ~new_G155_;
  assign G518 = ~new_G246_ | ~new_G450_ | ~new_G185_;
  assign G542 = ~new_G279_ | ~new_G243_ | ~new_G244_;
  assign new_G163_ = ~G0 & ~G4;
  assign new_G216_ = ~G4 & ~G5;
  assign new_G169_ = ~G5 & ~G7;
  assign new_G225_ = ~G7 & ~G8;
  assign new_G190_ = ~G7 & ~G11;
  assign new_G241_ = ~G10 & ~G11;
  assign new_G198_ = ~new_G520_ & ~G3;
  assign new_G178_ = ~new_G521_ & ~G4;
  assign new_G229_ = ~G1 & ~new_G522_;
  assign new_G209_ = ~G1 & ~new_G524_;
  assign new_G195_ = ~new_G521_ & ~new_G134_;
  assign new_G189_ = ~new_G522_ & ~new_G54_;
  assign new_G201_ = ~new_G528_ & ~new_G54_;
  assign new_G164_ = ~new_G531_ & ~G10;
  assign new_G211_ = ~G6 & ~new_G274_;
  assign new_G156_ = ~G12 & ~new_G543_;
  assign new_G205_ = ~new_G529_ & ~new_G122_;
  assign new_G227_ = ~G5 & ~new_G200_;
  assign new_G230_ = ~G8 & ~new_G490_;
  assign new_G191_ = ~G9 & ~new_G482_;
  assign new_G196_ = ~new_G86_ & ~G5 & ~new_G540_;
  assign new_G197_ = ~new_G540_ & ~new_G232_;
  assign new_G202_ = ~G10 & ~new_G63_;
  assign G502 = ~new_G436_ & ~new_G437_;
  assign new_G218_ = ~new_G528_ & ~new_G217_;
  assign G516 = ~new_G412_ & ~new_G410_ & ~new_G411_;
  assign G515 = ~new_G387_ & ~new_G388_;
  assign G509 = ~new_G331_ & ~G5;
  assign G513 = ~new_G360_ & ~new_G361_;
  assign new_G183_ = ~new_G330_ & ~G3;
  assign G517 = ~new_G428_ & ~new_G429_;
  assign new_G182_ = ~G12 & ~new_G62_;
  assign G519 = ~new_G463_ & ~new_G462_ & ~new_G460_ & ~new_G461_;
  assign new_G176_ = ~G4 & ~new_G494_;
  assign new_G175_ = ~new_G86_ & ~new_G500_;
  assign new_G187_ = ~G13 & ~new_G492_;
  assign new_G158_ = ~new_G521_ & ~new_G281_;
  assign new_G194_ = ~new_G281_ & ~new_G271_;
  assign new_G157_ = ~G13 & ~new_G483_;
  assign G507 = ~new_G487_ & ~new_G315_ & ~G12;
  assign new_G186_ = ~new_G282_ & ~new_G501_;
  assign new_G247_ = ~new_G474_ & ~new_G473_ & ~new_G471_ & ~new_G472_;
  assign new_G179_ = ~new_G541_ & ~new_G280_;
  assign new_G188_ = ~new_G543_ & ~new_G493_;
  assign new_G154_ = ~G12 & ~new_G488_;
  assign new_G184_ = ~new_G499_ & ~new_G541_ & ~G13;
  assign G506 = ~new_G311_ & ~new_G312_;
  assign new_G155_ = ~G13 & ~new_G480_;
  assign new_G162_ = ~new_G185_ & ~new_G498_;
  assign G514 = ~new_G478_ & ~new_G372_ & ~new_G373_;
endmodule


