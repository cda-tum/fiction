// Benchmark "top" written by ABC on Mon Feb 19 11:52:45 2024

module top ( 
    pa1, pb2, pp, pa0, pc2, pq, pb0, pc1, pr, pa2, pb1, pc0, ps, pd0, pe1,
    pf2, pt, pd1, pe0, pg2, pu, pd2, pf0, pg1, pv, pe2, pf1, pg0, pw, ph0,
    pi1, pj2, px, ph1, pi0, pk2, py, ph2, pk1, pz, pi2, pj1, pk0, pl0, pm1,
    pn2, pl1, pm0, po2, pl2, pn0, po1, pm2, pn1, po0, pp0, pq1, pr2, pa,
    pp1, pq0, ps2, pb, pp2, pr0, ps1, pq2, pr1, ps0, pt0, pu1, pv2, pt1,
    pu0, pt2, pv0, pw1, pg, pu2, pv1, pw0, ph, px0, py1, pi, px1, py0, pz0,
    pk, pz1, pl, pm, pn, po,
    pc3, pd4, pe5, pb3, pd5, pe4, pa3, pf4, pg5, pf5, pg4, pa5, pg3, pa4,
    pf3, pb4, pc5, pe3, pb5, pc4, pd3, pk3, pl4, pm5, pj3, pl5, pm4, pi3,
    pn4, po5, ph3, pn5, po4, ph4, pi5, po3, ph5, pi4, pn3, pj4, pk5, pm3,
    pj5, pk4, pl3, ps3, pt4, pr3, pu4, pq3, pv4, pp3, pw4, pp4, pw3, pq4,
    pv3, pw2, pr4, pu3, ps4, pt3, pz2, pz3, px2, py3, px3, py2, px4, py4,
    pz4  );
  input  pa1, pb2, pp, pa0, pc2, pq, pb0, pc1, pr, pa2, pb1, pc0, ps,
    pd0, pe1, pf2, pt, pd1, pe0, pg2, pu, pd2, pf0, pg1, pv, pe2, pf1, pg0,
    pw, ph0, pi1, pj2, px, ph1, pi0, pk2, py, ph2, pk1, pz, pi2, pj1, pk0,
    pl0, pm1, pn2, pl1, pm0, po2, pl2, pn0, po1, pm2, pn1, po0, pp0, pq1,
    pr2, pa, pp1, pq0, ps2, pb, pp2, pr0, ps1, pq2, pr1, ps0, pt0, pu1,
    pv2, pt1, pu0, pt2, pv0, pw1, pg, pu2, pv1, pw0, ph, px0, py1, pi, px1,
    py0, pz0, pk, pz1, pl, pm, pn, po;
  output pc3, pd4, pe5, pb3, pd5, pe4, pa3, pf4, pg5, pf5, pg4, pa5, pg3, pa4,
    pf3, pb4, pc5, pe3, pb5, pc4, pd3, pk3, pl4, pm5, pj3, pl5, pm4, pi3,
    pn4, po5, ph3, pn5, po4, ph4, pi5, po3, ph5, pi4, pn3, pj4, pk5, pm3,
    pj5, pk4, pl3, ps3, pt4, pr3, pu4, pq3, pv4, pp3, pw4, pp4, pw3, pq4,
    pv3, pw2, pr4, pu3, ps4, pt3, pz2, pz3, px2, py3, px3, py2, px4, py4,
    pz4;
  wire new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n262,
    new_n263, new_n264, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n340, new_n341, new_n342,
    new_n343, new_n344, new_n345, new_n346, new_n347, new_n348, new_n349,
    new_n350, new_n351, new_n352, new_n354, new_n355, new_n356, new_n357,
    new_n358, new_n359, new_n360, new_n361, new_n363, new_n364, new_n365,
    new_n366, new_n367, new_n368, new_n369, new_n370, new_n371, new_n372,
    new_n373, new_n374, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n389, new_n390, new_n391, new_n392, new_n393, new_n394, new_n395,
    new_n396, new_n397, new_n398, new_n399, new_n400, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n408, new_n410, new_n411, new_n412,
    new_n413, new_n414, new_n415, new_n416, new_n417, new_n418, new_n419,
    new_n421, new_n422, new_n423, new_n424, new_n425, new_n426, new_n427,
    new_n428, new_n429, new_n430, new_n431, new_n432, new_n434, new_n435,
    new_n436, new_n437, new_n438, new_n439, new_n440, new_n442, new_n444,
    new_n445, new_n446, new_n447, new_n448, new_n449, new_n450, new_n451,
    new_n452, new_n453, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n464, new_n466, new_n467, new_n468,
    new_n469, new_n470, new_n471, new_n472, new_n473, new_n474, new_n475,
    new_n476, new_n478, new_n479, new_n480, new_n481, new_n482, new_n483,
    new_n484, new_n485, new_n486, new_n487, new_n489, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n502, new_n503, new_n504, new_n505, new_n506, new_n507,
    new_n508, new_n509, new_n510, new_n511, new_n513, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914;
  assign new_n166 = ~ph0 & pt2;
  assign new_n167 = ph0 & ~pt2;
  assign new_n168 = ~pq2 & ~pi;
  assign new_n169 = ~new_n166 & ~new_n167;
  assign new_n170 = ~new_n168 & new_n169;
  assign new_n171 = pn2 & ~pp2;
  assign new_n172 = ~po2 & pr2;
  assign new_n173 = new_n171 & new_n172;
  assign new_n174 = pe1 & new_n170;
  assign new_n175 = new_n173 & new_n174;
  assign new_n176 = ~pi0 & new_n175;
  assign new_n177 = pe1 & ~new_n168;
  assign new_n178 = pn2 & ~po2;
  assign new_n179 = new_n177 & new_n178;
  assign new_n180 = pr2 & new_n179;
  assign new_n181 = ~pp2 & new_n180;
  assign new_n182 = ps2 & ~new_n181;
  assign new_n183 = ~pi0 & new_n182;
  assign pc3 = new_n176 | new_n183;
  assign new_n185 = po2 & ~pq2;
  assign new_n186 = ~pp2 & new_n185;
  assign new_n187 = ~pr2 & new_n186;
  assign new_n188 = ~pc1 & pk1;
  assign new_n189 = ~new_n187 & new_n188;
  assign new_n190 = ~pp2 & ~pq2;
  assign new_n191 = ~pr2 & new_n190;
  assign new_n192 = ~pn2 & new_n191;
  assign new_n193 = pe1 & po2;
  assign new_n194 = new_n192 & new_n193;
  assign new_n195 = ~pc1 & new_n194;
  assign new_n196 = pn2 & new_n195;
  assign new_n197 = ~pe1 & new_n188;
  assign new_n198 = pt0 & new_n188;
  assign new_n199 = pn2 & new_n188;
  assign new_n200 = ~new_n187 & new_n195;
  assign new_n201 = ~pe1 & new_n195;
  assign new_n202 = pt0 & new_n195;
  assign new_n203 = ~new_n189 & ~new_n196;
  assign new_n204 = ~new_n197 & ~new_n198;
  assign new_n205 = new_n203 & new_n204;
  assign new_n206 = ~new_n201 & ~new_n202;
  assign new_n207 = ~new_n199 & ~new_n200;
  assign new_n208 = new_n206 & new_n207;
  assign pd4 = ~new_n205 | ~new_n208;
  assign new_n210 = pb & ~pu0;
  assign new_n211 = ~pk2 & ~pl2;
  assign new_n212 = ~pk2 & pm2;
  assign new_n213 = ~new_n211 & ~new_n212;
  assign new_n214 = ~pc1 & new_n213;
  assign new_n215 = new_n210 & new_n214;
  assign new_n216 = ~pk2 & new_n215;
  assign new_n217 = ~pl2 & new_n215;
  assign new_n218 = pu2 & new_n214;
  assign new_n219 = ~pk2 & new_n218;
  assign new_n220 = ~pl2 & new_n218;
  assign new_n221 = pl2 & new_n214;
  assign new_n222 = ~pk2 & new_n221;
  assign new_n223 = ~pu2 & ~new_n210;
  assign new_n224 = new_n214 & new_n223;
  assign new_n225 = new_n210 & new_n224;
  assign new_n226 = pl2 & new_n224;
  assign new_n227 = pu2 & new_n224;
  assign new_n228 = ~new_n216 & ~new_n217;
  assign new_n229 = ~new_n219 & ~new_n220;
  assign new_n230 = new_n228 & new_n229;
  assign new_n231 = ~new_n226 & ~new_n227;
  assign new_n232 = ~new_n222 & ~new_n225;
  assign new_n233 = new_n231 & new_n232;
  assign pe5 = ~new_n230 | ~new_n233;
  assign new_n235 = pk2 & pu2;
  assign new_n236 = pk2 & pb;
  assign new_n237 = ~pu0 & new_n236;
  assign new_n238 = ~new_n235 & ~new_n237;
  assign new_n239 = ~pc1 & new_n238;
  assign new_n240 = pk2 & new_n239;
  assign new_n241 = new_n210 & new_n239;
  assign new_n242 = pu2 & new_n239;
  assign new_n243 = ~new_n240 & ~new_n241;
  assign pd5 = new_n242 | ~new_n243;
  assign new_n245 = ~po2 & ~pq2;
  assign new_n246 = ~pr2 & ~pp2;
  assign new_n247 = new_n245 & new_n246;
  assign new_n248 = pe1 & new_n247;
  assign new_n249 = pn2 & new_n248;
  assign new_n250 = ~pc1 & new_n249;
  assign new_n251 = ~pc1 & pl1;
  assign pe4 = new_n250 | new_n251;
  assign new_n253 = pg0 & pv2;
  assign new_n254 = ~pi0 & ~new_n253;
  assign new_n255 = pl2 & pm2;
  assign new_n256 = ~ph & new_n255;
  assign new_n257 = ~pk2 & ~pg;
  assign new_n258 = new_n256 & new_n257;
  assign new_n259 = new_n254 & new_n258;
  assign new_n260 = pm1 & new_n254;
  assign pf4 = new_n259 | new_n260;
  assign new_n262 = pn2 & pm2;
  assign new_n263 = pl2 & new_n262;
  assign new_n264 = ~pk2 & new_n263;
  assign new_n265 = pe1 & pn2;
  assign new_n266 = pd1 & pn2;
  assign new_n267 = ~new_n264 & ~new_n265;
  assign new_n268 = ~pc1 & ~new_n266;
  assign new_n269 = new_n267 & new_n268;
  assign new_n270 = ~pk2 & pl2;
  assign new_n271 = pm2 & new_n270;
  assign new_n272 = new_n269 & new_n271;
  assign new_n273 = pe1 & new_n269;
  assign new_n274 = pd1 & new_n269;
  assign new_n275 = pn2 & new_n269;
  assign new_n276 = ~new_n272 & ~new_n273;
  assign new_n277 = ~new_n274 & ~new_n275;
  assign pg5 = ~new_n276 | ~new_n277;
  assign new_n279 = ~pl2 & ~pm2;
  assign new_n280 = ~pk2 & ~pm2;
  assign new_n281 = ~new_n270 & ~new_n279;
  assign new_n282 = ~pc1 & ~new_n280;
  assign new_n283 = new_n281 & new_n282;
  assign new_n284 = new_n210 & new_n283;
  assign new_n285 = ~pl2 & new_n284;
  assign new_n286 = ~pm2 & new_n284;
  assign new_n287 = pu2 & new_n283;
  assign new_n288 = ~pl2 & new_n287;
  assign new_n289 = ~pm2 & new_n287;
  assign new_n290 = pm2 & new_n283;
  assign new_n291 = ~pl2 & new_n290;
  assign new_n292 = new_n223 & new_n283;
  assign new_n293 = new_n210 & new_n292;
  assign new_n294 = pm2 & new_n292;
  assign new_n295 = pu2 & new_n292;
  assign new_n296 = ~new_n285 & ~new_n286;
  assign new_n297 = ~new_n288 & ~new_n289;
  assign new_n298 = new_n296 & new_n297;
  assign new_n299 = ~new_n294 & ~new_n295;
  assign new_n300 = ~new_n291 & ~new_n293;
  assign new_n301 = new_n299 & new_n300;
  assign pf5 = ~new_n298 | ~new_n301;
  assign new_n303 = pg0 & pm1;
  assign new_n304 = pv2 & new_n303;
  assign new_n305 = ph & new_n304;
  assign new_n306 = ~ph0 & new_n304;
  assign new_n307 = pg & new_n304;
  assign new_n308 = ~new_n305 & ~new_n306;
  assign new_n309 = ~new_n307 & new_n308;
  assign new_n310 = pe1 & ~po1;
  assign new_n311 = ~pm0 & new_n309;
  assign new_n312 = new_n310 & new_n311;
  assign new_n313 = ~pi0 & new_n312;
  assign new_n314 = pm1 & pv2;
  assign new_n315 = pg0 & new_n314;
  assign new_n316 = pi & new_n315;
  assign new_n317 = ~pi0 & new_n316;
  assign new_n318 = ph & new_n303;
  assign new_n319 = pv2 & new_n318;
  assign new_n320 = ~ph0 & new_n315;
  assign new_n321 = pg & new_n303;
  assign new_n322 = pv2 & new_n321;
  assign new_n323 = pe1 & ~pm0;
  assign new_n324 = ~new_n319 & ~new_n320;
  assign new_n325 = ~new_n322 & ~new_n323;
  assign new_n326 = new_n324 & new_n325;
  assign new_n327 = pn1 & new_n326;
  assign new_n328 = ~pi0 & new_n327;
  assign new_n329 = ~new_n313 & ~new_n317;
  assign pg4 = new_n328 | ~new_n329;
  assign new_n331 = ~pg & ~pi;
  assign new_n332 = ~ph & new_n331;
  assign new_n333 = ph0 & new_n332;
  assign new_n334 = ~pi0 & pm1;
  assign new_n335 = pv2 & new_n334;
  assign new_n336 = pc0 & ~new_n333;
  assign new_n337 = new_n335 & new_n336;
  assign new_n338 = pg0 & new_n337;
  assign new_n339 = pe1 & pi2;
  assign new_n340 = pi & new_n304;
  assign new_n341 = ~new_n307 & ~new_n340;
  assign new_n342 = new_n308 & new_n341;
  assign new_n343 = ~pm0 & new_n339;
  assign new_n344 = new_n342 & new_n343;
  assign new_n345 = ~pi0 & new_n344;
  assign new_n346 = pm1 & ~new_n333;
  assign new_n347 = pg0 & new_n346;
  assign new_n348 = pv2 & new_n347;
  assign new_n349 = ~new_n323 & ~new_n348;
  assign new_n350 = ph2 & new_n349;
  assign new_n351 = ~pi0 & new_n350;
  assign new_n352 = ~new_n338 & ~new_n345;
  assign pa5 = new_n351 | ~new_n352;
  assign new_n354 = ~pn0 & ~new_n191;
  assign new_n355 = ~pn2 & ~pn0;
  assign new_n356 = ~pe1 & ~pn0;
  assign new_n357 = po2 & ~pn0;
  assign new_n358 = ~new_n354 & ~new_n355;
  assign new_n359 = ~new_n356 & ~new_n357;
  assign new_n360 = new_n358 & new_n359;
  assign new_n361 = ~pi0 & new_n360;
  assign pg3 = ~pc1 & new_n361;
  assign new_n363 = ~pc1 & ph1;
  assign new_n364 = ~new_n187 & new_n363;
  assign new_n365 = ~pe1 & new_n363;
  assign new_n366 = pq0 & new_n363;
  assign new_n367 = pn2 & new_n363;
  assign new_n368 = pq0 & new_n195;
  assign new_n369 = ~new_n196 & ~new_n364;
  assign new_n370 = ~new_n365 & ~new_n366;
  assign new_n371 = new_n369 & new_n370;
  assign new_n372 = ~new_n201 & ~new_n368;
  assign new_n373 = ~new_n200 & ~new_n367;
  assign new_n374 = new_n372 & new_n373;
  assign pa4 = ~new_n371 | ~new_n374;
  assign new_n376 = ~ph0 & pm1;
  assign new_n377 = pm1 & ph;
  assign new_n378 = pm1 & pi;
  assign new_n379 = pm1 & pg;
  assign new_n380 = ~new_n376 & ~new_n377;
  assign new_n381 = ~new_n378 & ~new_n379;
  assign new_n382 = new_n380 & new_n381;
  assign new_n383 = pg0 & new_n382;
  assign new_n384 = pv2 & new_n383;
  assign new_n385 = ~pi0 & new_n253;
  assign new_n386 = ~pi0 & ~pm0;
  assign new_n387 = ~new_n385 & ~new_n386;
  assign pf3 = new_n384 | new_n387;
  assign new_n389 = ~pc1 & pi1;
  assign new_n390 = ~new_n187 & new_n389;
  assign new_n391 = ~pe1 & new_n389;
  assign new_n392 = pr0 & new_n389;
  assign new_n393 = pn2 & new_n389;
  assign new_n394 = pr0 & new_n195;
  assign new_n395 = ~new_n196 & ~new_n390;
  assign new_n396 = ~new_n391 & ~new_n392;
  assign new_n397 = new_n395 & new_n396;
  assign new_n398 = ~new_n201 & ~new_n394;
  assign new_n399 = ~new_n200 & ~new_n393;
  assign new_n400 = new_n398 & new_n399;
  assign pb4 = ~new_n397 | ~new_n400;
  assign new_n402 = pe0 & ~new_n333;
  assign new_n403 = new_n335 & new_n402;
  assign new_n404 = pg0 & new_n403;
  assign new_n405 = ~pi0 & new_n349;
  assign new_n406 = pj2 & new_n405;
  assign pc5 = new_n404 | new_n406;
  assign new_n408 = ~pc1 & pl0;
  assign pe3 = new_n250 | new_n408;
  assign new_n410 = pd0 & ~new_n333;
  assign new_n411 = new_n335 & new_n410;
  assign new_n412 = pg0 & new_n411;
  assign new_n413 = pe1 & pj2;
  assign new_n414 = ~pm0 & new_n413;
  assign new_n415 = new_n342 & new_n414;
  assign new_n416 = ~pi0 & new_n415;
  assign new_n417 = pi2 & new_n349;
  assign new_n418 = ~pi0 & new_n417;
  assign new_n419 = ~new_n412 & ~new_n416;
  assign pb5 = new_n418 | ~new_n419;
  assign new_n421 = ~pc1 & pj1;
  assign new_n422 = ~new_n187 & new_n421;
  assign new_n423 = ~pe1 & new_n421;
  assign new_n424 = ps0 & new_n421;
  assign new_n425 = pn2 & new_n421;
  assign new_n426 = ps0 & new_n195;
  assign new_n427 = ~new_n196 & ~new_n422;
  assign new_n428 = ~new_n423 & ~new_n424;
  assign new_n429 = new_n427 & new_n428;
  assign new_n430 = ~new_n201 & ~new_n426;
  assign new_n431 = ~new_n200 & ~new_n425;
  assign new_n432 = new_n430 & new_n431;
  assign pc4 = ~new_n429 | ~new_n432;
  assign new_n434 = ~pc1 & new_n382;
  assign new_n435 = pg0 & new_n434;
  assign new_n436 = pv2 & new_n435;
  assign new_n437 = ~pf0 & ~pk0;
  assign new_n438 = ~pk0 & ~pv2;
  assign new_n439 = ~new_n437 & ~new_n438;
  assign new_n440 = ~pc1 & new_n439;
  assign pd3 = new_n436 | new_n440;
  assign new_n442 = ~pi0 & pr0;
  assign pk3 = ~pc1 & new_n442;
  assign new_n444 = pn & ~new_n333;
  assign new_n445 = new_n335 & new_n444;
  assign new_n446 = pg0 & new_n445;
  assign new_n447 = pe1 & pt1;
  assign new_n448 = ~pm0 & new_n447;
  assign new_n449 = new_n342 & new_n448;
  assign new_n450 = ~pi0 & new_n449;
  assign new_n451 = ps1 & new_n349;
  assign new_n452 = ~pi0 & new_n451;
  assign new_n453 = ~new_n446 & ~new_n450;
  assign pl4 = new_n452 | ~new_n453;
  assign new_n455 = ~ps2 & pt2;
  assign new_n456 = ~pc1 & new_n455;
  assign new_n457 = pl1 & ~pt2;
  assign new_n458 = ps2 & new_n457;
  assign new_n459 = ~pc1 & new_n458;
  assign new_n460 = ~pl1 & pt2;
  assign new_n461 = ~pc1 & new_n460;
  assign new_n462 = ~new_n456 & ~new_n459;
  assign pm5 = new_n461 | ~new_n462;
  assign new_n464 = ~pi0 & pq0;
  assign pj3 = ~pc1 & new_n464;
  assign new_n466 = ~pm0 & pn1;
  assign new_n467 = pe1 & new_n466;
  assign new_n468 = ~pi0 & new_n467;
  assign new_n469 = pb1 & ~pe1;
  assign new_n470 = ~pi0 & new_n469;
  assign new_n471 = pb1 & pn1;
  assign new_n472 = ~pi0 & new_n471;
  assign new_n473 = pb1 & pm0;
  assign new_n474 = ~pi0 & new_n473;
  assign new_n475 = ~new_n468 & ~new_n470;
  assign new_n476 = ~new_n472 & ~new_n474;
  assign pl5 = ~new_n475 | ~new_n476;
  assign new_n478 = po & ~new_n333;
  assign new_n479 = new_n335 & new_n478;
  assign new_n480 = pg0 & new_n479;
  assign new_n481 = pe1 & pu1;
  assign new_n482 = ~pm0 & new_n481;
  assign new_n483 = new_n342 & new_n482;
  assign new_n484 = ~pi0 & new_n483;
  assign new_n485 = pt1 & new_n349;
  assign new_n486 = ~pi0 & new_n485;
  assign new_n487 = ~new_n480 & ~new_n484;
  assign pm4 = new_n486 | ~new_n487;
  assign new_n489 = ~pi0 & pp0;
  assign pi3 = ~pc1 & new_n489;
  assign new_n491 = pp & ~new_n333;
  assign new_n492 = new_n335 & new_n491;
  assign new_n493 = pg0 & new_n492;
  assign new_n494 = pe1 & pv1;
  assign new_n495 = ~pm0 & new_n494;
  assign new_n496 = new_n342 & new_n495;
  assign new_n497 = ~pi0 & new_n496;
  assign new_n498 = pu1 & new_n349;
  assign new_n499 = ~pi0 & new_n498;
  assign new_n500 = ~new_n493 & ~new_n497;
  assign pn4 = new_n499 | ~new_n500;
  assign new_n502 = pv2 & new_n254;
  assign new_n503 = ~pf0 & new_n502;
  assign new_n504 = pr2 & ~pp2;
  assign new_n505 = ~po2 & new_n504;
  assign new_n506 = pq2 & new_n505;
  assign new_n507 = pi & new_n505;
  assign new_n508 = ~new_n506 & ~new_n507;
  assign new_n509 = pn2 & ~new_n508;
  assign new_n510 = pe1 & new_n509;
  assign new_n511 = new_n254 & new_n510;
  assign po5 = new_n503 | new_n511;
  assign new_n513 = ~pi0 & po0;
  assign ph3 = ~pc1 & new_n513;
  assign new_n515 = ~pb & ~pu2;
  assign new_n516 = pu0 & ~pu2;
  assign new_n517 = ~new_n515 & ~new_n516;
  assign new_n518 = ~pi0 & new_n517;
  assign new_n519 = new_n210 & new_n518;
  assign new_n520 = ~pl2 & new_n518;
  assign new_n521 = pk2 & new_n518;
  assign new_n522 = ~pm2 & new_n518;
  assign new_n523 = ~new_n519 & ~new_n520;
  assign new_n524 = ~new_n521 & ~new_n522;
  assign pn5 = ~new_n523 | ~new_n524;
  assign new_n526 = pq & ~new_n333;
  assign new_n527 = new_n335 & new_n526;
  assign new_n528 = pg0 & new_n527;
  assign new_n529 = pe1 & pw1;
  assign new_n530 = ~pm0 & new_n529;
  assign new_n531 = new_n342 & new_n530;
  assign new_n532 = ~pi0 & new_n531;
  assign new_n533 = pv1 & new_n349;
  assign new_n534 = ~pi0 & new_n533;
  assign new_n535 = ~new_n528 & ~new_n532;
  assign po4 = new_n534 | ~new_n535;
  assign new_n537 = ~pm0 & pp1;
  assign new_n538 = pe1 & new_n537;
  assign new_n539 = ~pi0 & new_n538;
  assign new_n540 = ~pe1 & ~po1;
  assign new_n541 = ~pi0 & new_n540;
  assign new_n542 = ~po1 & pp1;
  assign new_n543 = ~pi0 & new_n542;
  assign new_n544 = pm0 & ~po1;
  assign new_n545 = ~pi0 & new_n544;
  assign new_n546 = ~new_n539 & ~new_n541;
  assign new_n547 = ~new_n543 & ~new_n545;
  assign new_n548 = new_n546 & new_n547;
  assign ph4 = new_n348 | new_n548;
  assign new_n550 = ~pn2 & ~pp2;
  assign new_n551 = ~po2 & ~pp2;
  assign new_n552 = ~new_n550 & ~new_n551;
  assign new_n553 = ~pc1 & new_n552;
  assign new_n554 = pe1 & new_n553;
  assign new_n555 = ~po2 & new_n554;
  assign new_n556 = ~pp2 & new_n554;
  assign new_n557 = pp2 & new_n553;
  assign new_n558 = ~po2 & new_n557;
  assign new_n559 = ~pn2 & new_n554;
  assign new_n560 = ~pn2 & new_n557;
  assign new_n561 = ~pk2 & new_n255;
  assign new_n562 = ~pd1 & ~new_n561;
  assign new_n563 = ~pe1 & new_n562;
  assign new_n564 = new_n553 & new_n563;
  assign new_n565 = pe1 & new_n564;
  assign new_n566 = pd1 & new_n564;
  assign new_n567 = new_n271 & new_n564;
  assign new_n568 = new_n271 & new_n553;
  assign new_n569 = ~pp2 & new_n568;
  assign new_n570 = pp2 & new_n564;
  assign new_n571 = ~po2 & new_n568;
  assign new_n572 = pd1 & new_n553;
  assign new_n573 = ~pp2 & new_n572;
  assign new_n574 = ~pn2 & new_n568;
  assign new_n575 = ~pn2 & new_n572;
  assign new_n576 = ~po2 & new_n572;
  assign new_n577 = ~new_n555 & ~new_n556;
  assign new_n578 = ~new_n558 & ~new_n559;
  assign new_n579 = new_n577 & new_n578;
  assign new_n580 = ~new_n566 & ~new_n567;
  assign new_n581 = ~new_n560 & ~new_n565;
  assign new_n582 = new_n580 & new_n581;
  assign new_n583 = new_n579 & new_n582;
  assign new_n584 = ~new_n574 & ~new_n575;
  assign new_n585 = ~new_n576 & new_n584;
  assign new_n586 = ~new_n571 & ~new_n573;
  assign new_n587 = ~new_n569 & ~new_n570;
  assign new_n588 = new_n586 & new_n587;
  assign new_n589 = new_n585 & new_n588;
  assign pi5 = ~new_n583 | ~new_n589;
  assign po3 = ~pi0 & pa;
  assign new_n592 = ~pn2 & ~po2;
  assign new_n593 = ~pc1 & ~new_n592;
  assign new_n594 = pd1 & new_n593;
  assign new_n595 = ~pn2 & new_n594;
  assign new_n596 = ~po2 & new_n594;
  assign new_n597 = pe1 & new_n593;
  assign new_n598 = ~pn2 & new_n597;
  assign new_n599 = ~po2 & new_n597;
  assign new_n600 = po2 & new_n593;
  assign new_n601 = ~pn2 & new_n600;
  assign new_n602 = new_n563 & new_n593;
  assign new_n603 = new_n271 & new_n602;
  assign new_n604 = pd1 & new_n602;
  assign new_n605 = po2 & new_n602;
  assign new_n606 = pe1 & new_n602;
  assign new_n607 = new_n271 & new_n593;
  assign new_n608 = ~pn2 & new_n607;
  assign new_n609 = ~po2 & new_n607;
  assign new_n610 = ~new_n608 & ~new_n609;
  assign new_n611 = ~new_n604 & ~new_n605;
  assign new_n612 = ~new_n606 & new_n611;
  assign new_n613 = new_n610 & new_n612;
  assign new_n614 = ~new_n595 & ~new_n596;
  assign new_n615 = ~new_n598 & new_n614;
  assign new_n616 = ~new_n599 & ~new_n601;
  assign new_n617 = ~new_n603 & new_n616;
  assign new_n618 = new_n615 & new_n617;
  assign ph5 = ~new_n613 | ~new_n618;
  assign new_n620 = ~new_n333 & new_n335;
  assign new_n621 = pk & new_n620;
  assign new_n622 = pg0 & new_n621;
  assign new_n623 = pe1 & pq1;
  assign new_n624 = ~pm0 & new_n342;
  assign new_n625 = new_n623 & new_n624;
  assign new_n626 = ~pi0 & new_n625;
  assign new_n627 = pp1 & new_n349;
  assign new_n628 = ~pi0 & new_n627;
  assign new_n629 = ~new_n622 & ~new_n626;
  assign pi4 = new_n628 | ~new_n629;
  assign pn3 = ~pi0 & pb;
  assign new_n632 = pl & ~new_n333;
  assign new_n633 = new_n335 & new_n632;
  assign new_n634 = pg0 & new_n633;
  assign new_n635 = pe1 & pr1;
  assign new_n636 = ~pm0 & new_n635;
  assign new_n637 = new_n342 & new_n636;
  assign new_n638 = ~pi0 & new_n637;
  assign new_n639 = pq1 & new_n349;
  assign new_n640 = ~pi0 & new_n639;
  assign new_n641 = ~new_n634 & ~new_n638;
  assign pj4 = new_n640 | ~new_n641;
  assign new_n643 = pp2 & pq2;
  assign new_n644 = pr2 & new_n643;
  assign new_n645 = ~pc1 & ~new_n644;
  assign new_n646 = pr2 & new_n645;
  assign new_n647 = pn2 & pp2;
  assign new_n648 = po2 & pq2;
  assign new_n649 = new_n647 & new_n648;
  assign new_n650 = ~pc1 & pe1;
  assign new_n651 = new_n649 & new_n650;
  assign new_n652 = ~pn2 & new_n651;
  assign new_n653 = ~pc1 & pr2;
  assign new_n654 = ~po2 & new_n653;
  assign new_n655 = ~pc1 & new_n563;
  assign new_n656 = pr2 & new_n655;
  assign new_n657 = ~pn2 & new_n653;
  assign new_n658 = new_n649 & new_n655;
  assign new_n659 = new_n271 & new_n658;
  assign new_n660 = new_n645 & new_n649;
  assign new_n661 = pe1 & new_n660;
  assign new_n662 = pd1 & new_n660;
  assign new_n663 = new_n271 & new_n660;
  assign new_n664 = pe1 & new_n658;
  assign new_n665 = pd1 & new_n658;
  assign new_n666 = ~pc1 & new_n271;
  assign new_n667 = new_n649 & new_n666;
  assign new_n668 = ~po2 & new_n667;
  assign new_n669 = ~pc1 & pd1;
  assign new_n670 = new_n649 & new_n669;
  assign new_n671 = ~po2 & new_n670;
  assign new_n672 = ~pn2 & new_n667;
  assign new_n673 = ~po2 & new_n651;
  assign new_n674 = ~pn2 & new_n670;
  assign new_n675 = ~new_n646 & ~new_n652;
  assign new_n676 = ~new_n654 & ~new_n656;
  assign new_n677 = new_n675 & new_n676;
  assign new_n678 = ~new_n661 & ~new_n662;
  assign new_n679 = ~new_n657 & ~new_n659;
  assign new_n680 = new_n678 & new_n679;
  assign new_n681 = new_n677 & new_n680;
  assign new_n682 = ~new_n665 & ~new_n668;
  assign new_n683 = ~new_n663 & ~new_n664;
  assign new_n684 = new_n682 & new_n683;
  assign new_n685 = ~new_n671 & ~new_n672;
  assign new_n686 = ~new_n673 & ~new_n674;
  assign new_n687 = new_n685 & new_n686;
  assign new_n688 = new_n684 & new_n687;
  assign pk5 = ~new_n681 | ~new_n688;
  assign new_n690 = ~pi0 & pt0;
  assign pm3 = ~pc1 & new_n690;
  assign new_n692 = ~pn2 & ~pq2;
  assign new_n693 = ~new_n190 & ~new_n692;
  assign new_n694 = ~pc1 & ~new_n245;
  assign new_n695 = new_n693 & new_n694;
  assign new_n696 = pq2 & new_n695;
  assign new_n697 = new_n563 & new_n696;
  assign new_n698 = pe1 & new_n695;
  assign new_n699 = ~po2 & new_n698;
  assign new_n700 = ~pn2 & new_n696;
  assign new_n701 = ~new_n643 & new_n696;
  assign new_n702 = ~po2 & new_n696;
  assign new_n703 = new_n271 & new_n695;
  assign new_n704 = ~po2 & new_n703;
  assign new_n705 = ~pn2 & new_n703;
  assign new_n706 = ~new_n643 & new_n703;
  assign new_n707 = new_n563 & new_n703;
  assign new_n708 = pd1 & new_n695;
  assign new_n709 = ~new_n643 & new_n708;
  assign new_n710 = new_n563 & new_n708;
  assign new_n711 = ~pn2 & new_n708;
  assign new_n712 = new_n563 & new_n698;
  assign new_n713 = ~po2 & new_n708;
  assign new_n714 = ~pn2 & new_n698;
  assign new_n715 = ~new_n643 & new_n698;
  assign new_n716 = ~new_n697 & ~new_n699;
  assign new_n717 = ~new_n700 & ~new_n701;
  assign new_n718 = new_n716 & new_n717;
  assign new_n719 = ~new_n705 & ~new_n706;
  assign new_n720 = ~new_n702 & ~new_n704;
  assign new_n721 = new_n719 & new_n720;
  assign new_n722 = new_n718 & new_n721;
  assign new_n723 = ~new_n710 & ~new_n711;
  assign new_n724 = ~new_n707 & ~new_n709;
  assign new_n725 = new_n723 & new_n724;
  assign new_n726 = ~new_n712 & ~new_n713;
  assign new_n727 = ~new_n714 & ~new_n715;
  assign new_n728 = new_n726 & new_n727;
  assign new_n729 = new_n725 & new_n728;
  assign pj5 = ~new_n722 | ~new_n729;
  assign new_n731 = pm & ~new_n333;
  assign new_n732 = new_n335 & new_n731;
  assign new_n733 = pg0 & new_n732;
  assign new_n734 = pe1 & ps1;
  assign new_n735 = ~pm0 & new_n734;
  assign new_n736 = new_n342 & new_n735;
  assign new_n737 = ~pi0 & new_n736;
  assign new_n738 = pr1 & new_n349;
  assign new_n739 = ~pi0 & new_n738;
  assign new_n740 = ~new_n733 & ~new_n737;
  assign pk4 = new_n739 | ~new_n740;
  assign new_n742 = ~pi0 & ps0;
  assign pl3 = ~pc1 & new_n742;
  assign ps3 = ~pi0 & py0;
  assign new_n745 = pv & ~new_n333;
  assign new_n746 = new_n335 & new_n745;
  assign new_n747 = pg0 & new_n746;
  assign new_n748 = pb2 & pe1;
  assign new_n749 = ~pm0 & new_n748;
  assign new_n750 = new_n342 & new_n749;
  assign new_n751 = ~pi0 & new_n750;
  assign new_n752 = pa2 & new_n349;
  assign new_n753 = ~pi0 & new_n752;
  assign new_n754 = ~new_n747 & ~new_n751;
  assign pt4 = new_n753 | ~new_n754;
  assign pr3 = ~pi0 & px0;
  assign new_n757 = pw & ~new_n333;
  assign new_n758 = new_n335 & new_n757;
  assign new_n759 = pg0 & new_n758;
  assign new_n760 = pc2 & pe1;
  assign new_n761 = ~pm0 & new_n760;
  assign new_n762 = new_n342 & new_n761;
  assign new_n763 = ~pi0 & new_n762;
  assign new_n764 = pb2 & new_n349;
  assign new_n765 = ~pi0 & new_n764;
  assign new_n766 = ~new_n759 & ~new_n763;
  assign pu4 = new_n765 | ~new_n766;
  assign pq3 = ~pi0 & pw0;
  assign new_n769 = px & ~new_n333;
  assign new_n770 = new_n335 & new_n769;
  assign new_n771 = pg0 & new_n770;
  assign new_n772 = pe1 & pd2;
  assign new_n773 = ~pm0 & new_n772;
  assign new_n774 = new_n342 & new_n773;
  assign new_n775 = ~pi0 & new_n774;
  assign new_n776 = pc2 & new_n349;
  assign new_n777 = ~pi0 & new_n776;
  assign new_n778 = ~new_n771 & ~new_n775;
  assign pv4 = new_n777 | ~new_n778;
  assign pp3 = ~pi0 & pv0;
  assign new_n781 = py & ~new_n333;
  assign new_n782 = new_n335 & new_n781;
  assign new_n783 = pg0 & new_n782;
  assign new_n784 = pe1 & pe2;
  assign new_n785 = ~pm0 & new_n784;
  assign new_n786 = new_n342 & new_n785;
  assign new_n787 = ~pi0 & new_n786;
  assign new_n788 = pd2 & new_n349;
  assign new_n789 = ~pi0 & new_n788;
  assign new_n790 = ~new_n783 & ~new_n787;
  assign pw4 = new_n789 | ~new_n790;
  assign new_n792 = pr & ~new_n333;
  assign new_n793 = new_n335 & new_n792;
  assign new_n794 = pg0 & new_n793;
  assign new_n795 = pe1 & px1;
  assign new_n796 = ~pm0 & new_n795;
  assign new_n797 = new_n342 & new_n796;
  assign new_n798 = ~pi0 & new_n797;
  assign new_n799 = pw1 & new_n349;
  assign new_n800 = ~pi0 & new_n799;
  assign new_n801 = ~new_n794 & ~new_n798;
  assign pp4 = new_n800 | ~new_n801;
  assign new_n803 = ph0 & ~ph;
  assign new_n804 = ~pi & new_n803;
  assign new_n805 = ~pg & new_n804;
  assign new_n806 = ~pg0 & ~new_n805;
  assign new_n807 = pi0 & ~pm1;
  assign new_n808 = new_n806 & new_n807;
  assign pw3 = pv2 & new_n808;
  assign new_n810 = ps & ~new_n333;
  assign new_n811 = new_n335 & new_n810;
  assign new_n812 = pg0 & new_n811;
  assign new_n813 = pe1 & py1;
  assign new_n814 = ~pm0 & new_n813;
  assign new_n815 = new_n342 & new_n814;
  assign new_n816 = ~pi0 & new_n815;
  assign new_n817 = px1 & new_n349;
  assign new_n818 = ~pi0 & new_n817;
  assign new_n819 = ~new_n812 & ~new_n816;
  assign pq4 = new_n818 | ~new_n819;
  assign new_n821 = pr2 & new_n551;
  assign new_n822 = new_n177 & new_n821;
  assign new_n823 = pn2 & new_n822;
  assign new_n824 = ~pi0 & ~pv2;
  assign new_n825 = ~pf0 & ~pi0;
  assign new_n826 = ~new_n824 & ~new_n825;
  assign new_n827 = ~new_n384 & ~new_n823;
  assign pv3 = new_n826 | ~new_n827;
  assign new_n829 = pt & ~new_n333;
  assign new_n830 = new_n335 & new_n829;
  assign new_n831 = pg0 & new_n830;
  assign new_n832 = pe1 & pz1;
  assign new_n833 = ~pm0 & new_n832;
  assign new_n834 = new_n342 & new_n833;
  assign new_n835 = ~pi0 & new_n834;
  assign new_n836 = py1 & new_n349;
  assign new_n837 = ~pi0 & new_n836;
  assign new_n838 = ~new_n831 & ~new_n835;
  assign pr4 = new_n837 | ~new_n838;
  assign pu3 = pa1 & ~pi0;
  assign new_n841 = pu & ~new_n333;
  assign new_n842 = new_n335 & new_n841;
  assign new_n843 = pg0 & new_n842;
  assign new_n844 = pa2 & pe1;
  assign new_n845 = ~pm0 & new_n844;
  assign new_n846 = new_n342 & new_n845;
  assign new_n847 = ~pi0 & new_n846;
  assign new_n848 = pz1 & new_n349;
  assign new_n849 = ~pi0 & new_n848;
  assign new_n850 = ~new_n843 & ~new_n847;
  assign ps4 = new_n849 | ~new_n850;
  assign pt3 = ~pi0 & pz0;
  assign new_n853 = ~pc1 & pg1;
  assign new_n854 = ~new_n187 & new_n853;
  assign new_n855 = ~pe1 & new_n853;
  assign new_n856 = pp0 & new_n853;
  assign new_n857 = pn2 & new_n853;
  assign new_n858 = pp0 & new_n195;
  assign new_n859 = ~new_n196 & ~new_n854;
  assign new_n860 = ~new_n855 & ~new_n856;
  assign new_n861 = new_n859 & new_n860;
  assign new_n862 = ~new_n201 & ~new_n858;
  assign new_n863 = ~new_n200 & ~new_n857;
  assign new_n864 = new_n862 & new_n863;
  assign pz3 = ~new_n861 | ~new_n864;
  assign new_n866 = ~pc1 & pf1;
  assign new_n867 = ~new_n187 & new_n866;
  assign new_n868 = ~pe1 & new_n866;
  assign new_n869 = po0 & new_n866;
  assign new_n870 = pn2 & new_n866;
  assign new_n871 = po0 & new_n195;
  assign new_n872 = ~new_n196 & ~new_n867;
  assign new_n873 = ~new_n868 & ~new_n869;
  assign new_n874 = new_n872 & new_n873;
  assign new_n875 = ~new_n201 & ~new_n871;
  assign new_n876 = ~new_n200 & ~new_n870;
  assign new_n877 = new_n875 & new_n876;
  assign py3 = ~new_n874 | ~new_n877;
  assign new_n879 = pl2 & new_n212;
  assign new_n880 = ~pc1 & new_n879;
  assign new_n881 = ~new_n669 & ~new_n880;
  assign px3 = new_n650 | ~new_n881;
  assign new_n883 = pz & ~new_n333;
  assign new_n884 = new_n335 & new_n883;
  assign new_n885 = pg0 & new_n884;
  assign new_n886 = pe1 & pf2;
  assign new_n887 = ~pm0 & new_n886;
  assign new_n888 = new_n342 & new_n887;
  assign new_n889 = ~pi0 & new_n888;
  assign new_n890 = pe2 & new_n349;
  assign new_n891 = ~pi0 & new_n890;
  assign new_n892 = ~new_n885 & ~new_n889;
  assign px4 = new_n891 | ~new_n892;
  assign new_n894 = pa0 & ~new_n333;
  assign new_n895 = new_n335 & new_n894;
  assign new_n896 = pg0 & new_n895;
  assign new_n897 = pe1 & pg2;
  assign new_n898 = ~pm0 & new_n897;
  assign new_n899 = new_n342 & new_n898;
  assign new_n900 = ~pi0 & new_n899;
  assign new_n901 = pf2 & new_n349;
  assign new_n902 = ~pi0 & new_n901;
  assign new_n903 = ~new_n896 & ~new_n900;
  assign py4 = new_n902 | ~new_n903;
  assign new_n905 = pb0 & ~new_n333;
  assign new_n906 = new_n335 & new_n905;
  assign new_n907 = pg0 & new_n906;
  assign new_n908 = pe1 & ph2;
  assign new_n909 = ~pm0 & new_n908;
  assign new_n910 = new_n342 & new_n909;
  assign new_n911 = ~pi0 & new_n910;
  assign new_n912 = pg2 & new_n349;
  assign new_n913 = ~pi0 & new_n912;
  assign new_n914 = ~new_n907 & ~new_n911;
  assign pz4 = new_n913 | ~new_n914;
  assign pb3 = ~pk1;
  assign pa3 = ~pj1;
  assign pw2 = ~pf1;
  assign pz2 = ~pi1;
  assign px2 = ~pg1;
  assign py2 = ~ph1;
endmodule


