// Benchmark "top" written by ABC on Mon Feb 19 11:52:42 2024

module top ( 
    ic3_35_, ic7_39_, id4_4_, id22_22_, id26_26_, id21_21_, id27_27_,
    id29_29_, ic4_36_, id5_5_, id20_20_, id28_28_, ic6_38_, id6_6_,
    id17_17_, id31_31_, id18_18_, id23_23_, id25_25_, id30_30_, ic0_32_,
    id7_7_, id19_19_, id24_24_, ic1_33_, ic5_37_, r_40_, id0_0_, id8_8_,
    id14_14_, id16_16_, id1_1_, id9_9_, id15_15_, ic2_34_, id2_2_,
    id13_13_, id10_10_, id12_12_, id3_3_, id11_11_,
    od10_232_, od11_231_, od12_230_, od4_238_, od8_234_, od1_241_,
    od20_222_, od21_221_, od22_220_, od5_237_, od9_233_, od2_240_,
    od23_219_, od24_218_, od25_217_, od26_216_, od27_215_, od28_214_,
    od29_213_, od30_212_, od31_211_, od6_236_, od13_229_, od14_228_,
    od15_227_, od16_226_, od17_225_, od18_224_, od19_223_, od3_239_,
    od7_235_, od0_242_  );
  input  ic3_35_, ic7_39_, id4_4_, id22_22_, id26_26_, id21_21_,
    id27_27_, id29_29_, ic4_36_, id5_5_, id20_20_, id28_28_, ic6_38_,
    id6_6_, id17_17_, id31_31_, id18_18_, id23_23_, id25_25_, id30_30_,
    ic0_32_, id7_7_, id19_19_, id24_24_, ic1_33_, ic5_37_, r_40_, id0_0_,
    id8_8_, id14_14_, id16_16_, id1_1_, id9_9_, id15_15_, ic2_34_, id2_2_,
    id13_13_, id10_10_, id12_12_, id3_3_, id11_11_;
  output od10_232_, od11_231_, od12_230_, od4_238_, od8_234_, od1_241_,
    od20_222_, od21_221_, od22_220_, od5_237_, od9_233_, od2_240_,
    od23_219_, od24_218_, od25_217_, od26_216_, od27_215_, od28_214_,
    od29_213_, od30_212_, od31_211_, od6_236_, od13_229_, od14_228_,
    od15_227_, od16_226_, od17_225_, od18_224_, od19_223_, od3_239_,
    od7_235_, od0_242_;
  wire new_n74, new_n75, new_n76, new_n77, new_n78, new_n79, new_n80,
    new_n81, new_n82, new_n83, new_n84, new_n85, new_n86, new_n87, new_n88,
    new_n89, new_n90, new_n91, new_n92, new_n93, new_n94, new_n95, new_n96,
    new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n140, new_n141, new_n142, new_n143, new_n144, new_n145,
    new_n146, new_n147, new_n148, new_n149, new_n150, new_n151, new_n152,
    new_n153, new_n154, new_n155, new_n156, new_n157, new_n158, new_n159,
    new_n160, new_n161, new_n162, new_n163, new_n164, new_n165, new_n166,
    new_n167, new_n168, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n320, new_n321,
    new_n322, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n332, new_n333, new_n334, new_n335, new_n336, new_n337,
    new_n339, new_n340, new_n341, new_n343, new_n344, new_n345, new_n346,
    new_n347, new_n348, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n372, new_n373, new_n374, new_n376, new_n377,
    new_n378, new_n380, new_n381, new_n382, new_n384, new_n385, new_n386,
    new_n388, new_n389, new_n390, new_n392, new_n393, new_n394, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n404,
    new_n405, new_n406, new_n408, new_n409, new_n410, new_n412, new_n413,
    new_n414, new_n416, new_n417, new_n418, new_n419, new_n420, new_n421,
    new_n423, new_n424, new_n425, new_n427, new_n428, new_n429, new_n431,
    new_n432, new_n433, new_n435, new_n436, new_n437, new_n439, new_n440,
    new_n441, new_n443, new_n444, new_n445, new_n447, new_n448, new_n449,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n458,
    new_n459, new_n460, new_n462, new_n463, new_n464, new_n466, new_n467,
    new_n468, new_n470, new_n471, new_n472, new_n474, new_n475, new_n476,
    new_n478, new_n479, new_n480;
  assign new_n74 = id14_14_ & ~id15_15_;
  assign new_n75 = ~id14_14_ & id15_15_;
  assign new_n76 = ~new_n74 & ~new_n75;
  assign new_n77 = ~id13_13_ & id12_12_;
  assign new_n78 = id13_13_ & ~id12_12_;
  assign new_n79 = ~new_n77 & ~new_n78;
  assign new_n80 = new_n76 & ~new_n79;
  assign new_n81 = ~new_n76 & new_n79;
  assign new_n82 = ~new_n80 & ~new_n81;
  assign new_n83 = id6_6_ & ~id7_7_;
  assign new_n84 = ~id6_6_ & id7_7_;
  assign new_n85 = ~new_n83 & ~new_n84;
  assign new_n86 = id4_4_ & ~id5_5_;
  assign new_n87 = ~id4_4_ & id5_5_;
  assign new_n88 = ~new_n86 & ~new_n87;
  assign new_n89 = new_n85 & ~new_n88;
  assign new_n90 = ~new_n85 & new_n88;
  assign new_n91 = ~new_n89 & ~new_n90;
  assign new_n92 = new_n82 & ~new_n91;
  assign new_n93 = ~new_n82 & new_n91;
  assign new_n94 = ~new_n92 & ~new_n93;
  assign new_n95 = ic7_39_ & r_40_;
  assign new_n96 = new_n94 & new_n95;
  assign new_n97 = ~new_n94 & ~new_n95;
  assign new_n98 = ~new_n96 & ~new_n97;
  assign new_n99 = id27_27_ & ~id31_31_;
  assign new_n100 = ~id27_27_ & id31_31_;
  assign new_n101 = ~new_n99 & ~new_n100;
  assign new_n102 = ~id23_23_ & id19_19_;
  assign new_n103 = id23_23_ & ~id19_19_;
  assign new_n104 = ~new_n102 & ~new_n103;
  assign new_n105 = new_n101 & ~new_n104;
  assign new_n106 = ~new_n101 & new_n104;
  assign new_n107 = ~new_n105 & ~new_n106;
  assign new_n108 = new_n98 & ~new_n107;
  assign new_n109 = ~new_n98 & new_n107;
  assign new_n110 = ~new_n108 & ~new_n109;
  assign new_n111 = ~id31_31_ & id30_30_;
  assign new_n112 = id31_31_ & ~id30_30_;
  assign new_n113 = ~new_n111 & ~new_n112;
  assign new_n114 = ~id29_29_ & id28_28_;
  assign new_n115 = id29_29_ & ~id28_28_;
  assign new_n116 = ~new_n114 & ~new_n115;
  assign new_n117 = new_n113 & ~new_n116;
  assign new_n118 = ~new_n113 & new_n116;
  assign new_n119 = ~new_n117 & ~new_n118;
  assign new_n120 = id22_22_ & ~id23_23_;
  assign new_n121 = ~id22_22_ & id23_23_;
  assign new_n122 = ~new_n120 & ~new_n121;
  assign new_n123 = ~id21_21_ & id20_20_;
  assign new_n124 = id21_21_ & ~id20_20_;
  assign new_n125 = ~new_n123 & ~new_n124;
  assign new_n126 = new_n122 & ~new_n125;
  assign new_n127 = ~new_n122 & new_n125;
  assign new_n128 = ~new_n126 & ~new_n127;
  assign new_n129 = new_n119 & ~new_n128;
  assign new_n130 = ~new_n119 & new_n128;
  assign new_n131 = ~new_n129 & ~new_n130;
  assign new_n132 = ic3_35_ & r_40_;
  assign new_n133 = new_n131 & new_n132;
  assign new_n134 = ~new_n131 & ~new_n132;
  assign new_n135 = ~new_n133 & ~new_n134;
  assign new_n136 = ~id15_15_ & id11_11_;
  assign new_n137 = id15_15_ & ~id11_11_;
  assign new_n138 = ~new_n136 & ~new_n137;
  assign new_n139 = ~id7_7_ & id3_3_;
  assign new_n140 = id7_7_ & ~id3_3_;
  assign new_n141 = ~new_n139 & ~new_n140;
  assign new_n142 = new_n138 & ~new_n141;
  assign new_n143 = ~new_n138 & new_n141;
  assign new_n144 = ~new_n142 & ~new_n143;
  assign new_n145 = new_n135 & ~new_n144;
  assign new_n146 = ~new_n135 & new_n144;
  assign new_n147 = ~new_n145 & ~new_n146;
  assign new_n148 = id26_26_ & ~id27_27_;
  assign new_n149 = ~id26_26_ & id27_27_;
  assign new_n150 = ~new_n148 & ~new_n149;
  assign new_n151 = ~id25_25_ & id24_24_;
  assign new_n152 = id25_25_ & ~id24_24_;
  assign new_n153 = ~new_n151 & ~new_n152;
  assign new_n154 = new_n150 & ~new_n153;
  assign new_n155 = ~new_n150 & new_n153;
  assign new_n156 = ~new_n154 & ~new_n155;
  assign new_n157 = new_n119 & ~new_n156;
  assign new_n158 = ~new_n119 & new_n156;
  assign new_n159 = ~new_n157 & ~new_n158;
  assign new_n160 = ic1_33_ & r_40_;
  assign new_n161 = new_n159 & new_n160;
  assign new_n162 = ~new_n159 & ~new_n160;
  assign new_n163 = ~new_n161 & ~new_n162;
  assign new_n164 = id9_9_ & ~id13_13_;
  assign new_n165 = ~id9_9_ & id13_13_;
  assign new_n166 = ~new_n164 & ~new_n165;
  assign new_n167 = ~id5_5_ & id1_1_;
  assign new_n168 = id5_5_ & ~id1_1_;
  assign new_n169 = ~new_n167 & ~new_n168;
  assign new_n170 = new_n166 & ~new_n169;
  assign new_n171 = ~new_n166 & new_n169;
  assign new_n172 = ~new_n170 & ~new_n171;
  assign new_n173 = new_n163 & ~new_n172;
  assign new_n174 = ~new_n163 & new_n172;
  assign new_n175 = ~new_n173 & ~new_n174;
  assign new_n176 = id18_18_ & ~id19_19_;
  assign new_n177 = ~id18_18_ & id19_19_;
  assign new_n178 = ~new_n176 & ~new_n177;
  assign new_n179 = ~id17_17_ & id16_16_;
  assign new_n180 = id17_17_ & ~id16_16_;
  assign new_n181 = ~new_n179 & ~new_n180;
  assign new_n182 = new_n178 & ~new_n181;
  assign new_n183 = ~new_n178 & new_n181;
  assign new_n184 = ~new_n182 & ~new_n183;
  assign new_n185 = new_n156 & ~new_n184;
  assign new_n186 = ~new_n156 & new_n184;
  assign new_n187 = ~new_n185 & ~new_n186;
  assign new_n188 = r_40_ & ic2_34_;
  assign new_n189 = new_n187 & new_n188;
  assign new_n190 = ~new_n187 & ~new_n188;
  assign new_n191 = ~new_n189 & ~new_n190;
  assign new_n192 = ~id14_14_ & id10_10_;
  assign new_n193 = id14_14_ & ~id10_10_;
  assign new_n194 = ~new_n192 & ~new_n193;
  assign new_n195 = ~id6_6_ & id2_2_;
  assign new_n196 = id6_6_ & ~id2_2_;
  assign new_n197 = ~new_n195 & ~new_n196;
  assign new_n198 = new_n194 & ~new_n197;
  assign new_n199 = ~new_n194 & new_n197;
  assign new_n200 = ~new_n198 & ~new_n199;
  assign new_n201 = new_n191 & ~new_n200;
  assign new_n202 = ~new_n191 & new_n200;
  assign new_n203 = ~new_n201 & ~new_n202;
  assign new_n204 = new_n128 & ~new_n184;
  assign new_n205 = ~new_n128 & new_n184;
  assign new_n206 = ~new_n204 & ~new_n205;
  assign new_n207 = ic0_32_ & r_40_;
  assign new_n208 = new_n206 & new_n207;
  assign new_n209 = ~new_n206 & ~new_n207;
  assign new_n210 = ~new_n208 & ~new_n209;
  assign new_n211 = id8_8_ & ~id12_12_;
  assign new_n212 = ~id8_8_ & id12_12_;
  assign new_n213 = ~new_n211 & ~new_n212;
  assign new_n214 = ~id4_4_ & id0_0_;
  assign new_n215 = id4_4_ & ~id0_0_;
  assign new_n216 = ~new_n214 & ~new_n215;
  assign new_n217 = new_n213 & ~new_n216;
  assign new_n218 = ~new_n213 & new_n216;
  assign new_n219 = ~new_n217 & ~new_n218;
  assign new_n220 = new_n210 & ~new_n219;
  assign new_n221 = ~new_n210 & new_n219;
  assign new_n222 = ~new_n220 & ~new_n221;
  assign new_n223 = new_n147 & new_n175;
  assign new_n224 = new_n203 & new_n223;
  assign new_n225 = ~new_n222 & new_n224;
  assign new_n226 = ~new_n203 & new_n223;
  assign new_n227 = new_n222 & new_n226;
  assign new_n228 = new_n147 & ~new_n175;
  assign new_n229 = new_n203 & new_n228;
  assign new_n230 = new_n222 & new_n229;
  assign new_n231 = ~new_n147 & new_n175;
  assign new_n232 = new_n203 & new_n231;
  assign new_n233 = new_n222 & new_n232;
  assign new_n234 = ~new_n225 & ~new_n227;
  assign new_n235 = ~new_n230 & new_n234;
  assign new_n236 = ~new_n233 & new_n235;
  assign new_n237 = id10_10_ & ~id11_11_;
  assign new_n238 = ~id10_10_ & id11_11_;
  assign new_n239 = ~new_n237 & ~new_n238;
  assign new_n240 = id8_8_ & ~id9_9_;
  assign new_n241 = ~id8_8_ & id9_9_;
  assign new_n242 = ~new_n240 & ~new_n241;
  assign new_n243 = new_n239 & ~new_n242;
  assign new_n244 = ~new_n239 & new_n242;
  assign new_n245 = ~new_n243 & ~new_n244;
  assign new_n246 = new_n82 & ~new_n245;
  assign new_n247 = ~new_n82 & new_n245;
  assign new_n248 = ~new_n246 & ~new_n247;
  assign new_n249 = ic5_37_ & r_40_;
  assign new_n250 = new_n248 & new_n249;
  assign new_n251 = ~new_n248 & ~new_n249;
  assign new_n252 = ~new_n250 & ~new_n251;
  assign new_n253 = ~id29_29_ & id25_25_;
  assign new_n254 = id29_29_ & ~id25_25_;
  assign new_n255 = ~new_n253 & ~new_n254;
  assign new_n256 = ~id21_21_ & id17_17_;
  assign new_n257 = id21_21_ & ~id17_17_;
  assign new_n258 = ~new_n256 & ~new_n257;
  assign new_n259 = new_n255 & ~new_n258;
  assign new_n260 = ~new_n255 & new_n258;
  assign new_n261 = ~new_n259 & ~new_n260;
  assign new_n262 = new_n252 & ~new_n261;
  assign new_n263 = ~new_n252 & new_n261;
  assign new_n264 = ~new_n262 & ~new_n263;
  assign new_n265 = id2_2_ & ~id3_3_;
  assign new_n266 = ~id2_2_ & id3_3_;
  assign new_n267 = ~new_n265 & ~new_n266;
  assign new_n268 = id0_0_ & ~id1_1_;
  assign new_n269 = ~id0_0_ & id1_1_;
  assign new_n270 = ~new_n268 & ~new_n269;
  assign new_n271 = new_n267 & ~new_n270;
  assign new_n272 = ~new_n267 & new_n270;
  assign new_n273 = ~new_n271 & ~new_n272;
  assign new_n274 = new_n245 & ~new_n273;
  assign new_n275 = ~new_n245 & new_n273;
  assign new_n276 = ~new_n274 & ~new_n275;
  assign new_n277 = ic6_38_ & r_40_;
  assign new_n278 = new_n276 & new_n277;
  assign new_n279 = ~new_n276 & ~new_n277;
  assign new_n280 = ~new_n278 & ~new_n279;
  assign new_n281 = id26_26_ & ~id30_30_;
  assign new_n282 = ~id26_26_ & id30_30_;
  assign new_n283 = ~new_n281 & ~new_n282;
  assign new_n284 = ~id22_22_ & id18_18_;
  assign new_n285 = id22_22_ & ~id18_18_;
  assign new_n286 = ~new_n284 & ~new_n285;
  assign new_n287 = new_n283 & ~new_n286;
  assign new_n288 = ~new_n283 & new_n286;
  assign new_n289 = ~new_n287 & ~new_n288;
  assign new_n290 = new_n280 & ~new_n289;
  assign new_n291 = ~new_n280 & new_n289;
  assign new_n292 = ~new_n290 & ~new_n291;
  assign new_n293 = new_n91 & ~new_n273;
  assign new_n294 = ~new_n91 & new_n273;
  assign new_n295 = ~new_n293 & ~new_n294;
  assign new_n296 = ic4_36_ & r_40_;
  assign new_n297 = new_n295 & new_n296;
  assign new_n298 = ~new_n295 & ~new_n296;
  assign new_n299 = ~new_n297 & ~new_n298;
  assign new_n300 = ~id28_28_ & id24_24_;
  assign new_n301 = id28_28_ & ~id24_24_;
  assign new_n302 = ~new_n300 & ~new_n301;
  assign new_n303 = ~id20_20_ & id16_16_;
  assign new_n304 = id20_20_ & ~id16_16_;
  assign new_n305 = ~new_n303 & ~new_n304;
  assign new_n306 = new_n302 & ~new_n305;
  assign new_n307 = ~new_n302 & new_n305;
  assign new_n308 = ~new_n306 & ~new_n307;
  assign new_n309 = new_n299 & ~new_n308;
  assign new_n310 = ~new_n299 & new_n308;
  assign new_n311 = ~new_n309 & ~new_n310;
  assign new_n312 = new_n110 & ~new_n236;
  assign new_n313 = ~new_n264 & new_n312;
  assign new_n314 = ~new_n292 & new_n313;
  assign new_n315 = new_n311 & new_n314;
  assign new_n316 = ~new_n203 & new_n315;
  assign new_n317 = id10_10_ & ~new_n316;
  assign new_n318 = ~id10_10_ & new_n316;
  assign od10_232_ = new_n317 | new_n318;
  assign new_n320 = ~new_n147 & new_n315;
  assign new_n321 = id11_11_ & ~new_n320;
  assign new_n322 = ~id11_11_ & new_n320;
  assign od11_231_ = new_n321 | new_n322;
  assign new_n324 = ~new_n110 & ~new_n236;
  assign new_n325 = ~new_n264 & new_n324;
  assign new_n326 = new_n292 & new_n325;
  assign new_n327 = new_n311 & new_n326;
  assign new_n328 = ~new_n222 & new_n327;
  assign new_n329 = id12_12_ & ~new_n328;
  assign new_n330 = ~id12_12_ & new_n328;
  assign od12_230_ = new_n329 | new_n330;
  assign new_n332 = new_n264 & new_n324;
  assign new_n333 = new_n292 & new_n332;
  assign new_n334 = ~new_n311 & new_n333;
  assign new_n335 = ~new_n222 & new_n334;
  assign new_n336 = id4_4_ & ~new_n335;
  assign new_n337 = ~id4_4_ & new_n335;
  assign od4_238_ = new_n336 | new_n337;
  assign new_n339 = ~new_n222 & new_n315;
  assign new_n340 = id8_8_ & ~new_n339;
  assign new_n341 = ~id8_8_ & new_n339;
  assign od8_234_ = new_n340 | new_n341;
  assign new_n343 = new_n264 & new_n312;
  assign new_n344 = ~new_n292 & new_n343;
  assign new_n345 = ~new_n311 & new_n344;
  assign new_n346 = ~new_n175 & new_n345;
  assign new_n347 = id1_1_ & ~new_n346;
  assign new_n348 = ~id1_1_ & new_n346;
  assign od1_241_ = new_n347 | new_n348;
  assign new_n350 = new_n110 & new_n264;
  assign new_n351 = new_n292 & new_n350;
  assign new_n352 = ~new_n311 & new_n351;
  assign new_n353 = ~new_n292 & new_n350;
  assign new_n354 = new_n311 & new_n353;
  assign new_n355 = new_n110 & ~new_n264;
  assign new_n356 = new_n292 & new_n355;
  assign new_n357 = new_n311 & new_n356;
  assign new_n358 = ~new_n110 & new_n264;
  assign new_n359 = new_n292 & new_n358;
  assign new_n360 = new_n311 & new_n359;
  assign new_n361 = ~new_n352 & ~new_n354;
  assign new_n362 = ~new_n357 & new_n361;
  assign new_n363 = ~new_n360 & new_n362;
  assign new_n364 = ~new_n147 & ~new_n363;
  assign new_n365 = new_n175 & new_n364;
  assign new_n366 = new_n203 & new_n365;
  assign new_n367 = ~new_n222 & new_n366;
  assign new_n368 = ~new_n311 & new_n367;
  assign new_n369 = id20_20_ & ~new_n368;
  assign new_n370 = ~id20_20_ & new_n368;
  assign od20_222_ = new_n369 | new_n370;
  assign new_n372 = ~new_n264 & new_n367;
  assign new_n373 = id21_21_ & ~new_n372;
  assign new_n374 = ~id21_21_ & new_n372;
  assign od21_221_ = new_n373 | new_n374;
  assign new_n376 = ~new_n292 & new_n367;
  assign new_n377 = id22_22_ & ~new_n376;
  assign new_n378 = ~id22_22_ & new_n376;
  assign od22_220_ = new_n377 | new_n378;
  assign new_n380 = ~new_n175 & new_n334;
  assign new_n381 = id5_5_ & ~new_n380;
  assign new_n382 = ~id5_5_ & new_n380;
  assign od5_237_ = new_n381 | new_n382;
  assign new_n384 = ~new_n175 & new_n315;
  assign new_n385 = id9_9_ & ~new_n384;
  assign new_n386 = ~id9_9_ & new_n384;
  assign od9_233_ = new_n385 | new_n386;
  assign new_n388 = ~new_n203 & new_n345;
  assign new_n389 = id2_2_ & ~new_n388;
  assign new_n390 = ~id2_2_ & new_n388;
  assign od2_240_ = new_n389 | new_n390;
  assign new_n392 = ~new_n110 & new_n367;
  assign new_n393 = id23_23_ & ~new_n392;
  assign new_n394 = ~id23_23_ & new_n392;
  assign od23_219_ = new_n393 | new_n394;
  assign new_n396 = new_n147 & ~new_n363;
  assign new_n397 = ~new_n175 & new_n396;
  assign new_n398 = ~new_n203 & new_n397;
  assign new_n399 = new_n222 & new_n398;
  assign new_n400 = ~new_n311 & new_n399;
  assign new_n401 = id24_24_ & ~new_n400;
  assign new_n402 = ~id24_24_ & new_n400;
  assign od24_218_ = new_n401 | new_n402;
  assign new_n404 = ~new_n264 & new_n399;
  assign new_n405 = id25_25_ & ~new_n404;
  assign new_n406 = ~id25_25_ & new_n404;
  assign od25_217_ = new_n405 | new_n406;
  assign new_n408 = ~new_n292 & new_n399;
  assign new_n409 = id26_26_ & ~new_n408;
  assign new_n410 = ~id26_26_ & new_n408;
  assign od26_216_ = new_n409 | new_n410;
  assign new_n412 = ~new_n110 & new_n399;
  assign new_n413 = id27_27_ & ~new_n412;
  assign new_n414 = ~id27_27_ & new_n412;
  assign od27_215_ = new_n413 | new_n414;
  assign new_n416 = ~new_n175 & new_n364;
  assign new_n417 = new_n203 & new_n416;
  assign new_n418 = new_n222 & new_n417;
  assign new_n419 = ~new_n311 & new_n418;
  assign new_n420 = id28_28_ & ~new_n419;
  assign new_n421 = ~id28_28_ & new_n419;
  assign od28_214_ = new_n420 | new_n421;
  assign new_n423 = ~new_n264 & new_n418;
  assign new_n424 = id29_29_ & ~new_n423;
  assign new_n425 = ~id29_29_ & new_n423;
  assign od29_213_ = new_n424 | new_n425;
  assign new_n427 = ~new_n292 & new_n418;
  assign new_n428 = id30_30_ & ~new_n427;
  assign new_n429 = ~id30_30_ & new_n427;
  assign od30_212_ = new_n428 | new_n429;
  assign new_n431 = ~new_n110 & new_n418;
  assign new_n432 = id31_31_ & ~new_n431;
  assign new_n433 = ~id31_31_ & new_n431;
  assign od31_211_ = new_n432 | new_n433;
  assign new_n435 = ~new_n203 & new_n334;
  assign new_n436 = id6_6_ & ~new_n435;
  assign new_n437 = ~id6_6_ & new_n435;
  assign od6_236_ = new_n436 | new_n437;
  assign new_n439 = ~new_n175 & new_n327;
  assign new_n440 = id13_13_ & ~new_n439;
  assign new_n441 = ~id13_13_ & new_n439;
  assign od13_229_ = new_n440 | new_n441;
  assign new_n443 = ~new_n203 & new_n327;
  assign new_n444 = id14_14_ & ~new_n443;
  assign new_n445 = ~id14_14_ & new_n443;
  assign od14_228_ = new_n444 | new_n445;
  assign new_n447 = ~new_n147 & new_n327;
  assign new_n448 = id15_15_ & ~new_n447;
  assign new_n449 = ~id15_15_ & new_n447;
  assign od15_227_ = new_n448 | new_n449;
  assign new_n451 = new_n175 & new_n396;
  assign new_n452 = ~new_n203 & new_n451;
  assign new_n453 = ~new_n222 & new_n452;
  assign new_n454 = ~new_n311 & new_n453;
  assign new_n455 = id16_16_ & ~new_n454;
  assign new_n456 = ~id16_16_ & new_n454;
  assign od16_226_ = new_n455 | new_n456;
  assign new_n458 = ~new_n264 & new_n453;
  assign new_n459 = id17_17_ & ~new_n458;
  assign new_n460 = ~id17_17_ & new_n458;
  assign od17_225_ = new_n459 | new_n460;
  assign new_n462 = ~new_n292 & new_n453;
  assign new_n463 = id18_18_ & ~new_n462;
  assign new_n464 = ~id18_18_ & new_n462;
  assign od18_224_ = new_n463 | new_n464;
  assign new_n466 = ~new_n110 & new_n453;
  assign new_n467 = id19_19_ & ~new_n466;
  assign new_n468 = ~id19_19_ & new_n466;
  assign od19_223_ = new_n467 | new_n468;
  assign new_n470 = ~new_n147 & new_n345;
  assign new_n471 = id3_3_ & ~new_n470;
  assign new_n472 = ~id3_3_ & new_n470;
  assign od3_239_ = new_n471 | new_n472;
  assign new_n474 = ~new_n147 & new_n334;
  assign new_n475 = id7_7_ & ~new_n474;
  assign new_n476 = ~id7_7_ & new_n474;
  assign od7_235_ = new_n475 | new_n476;
  assign new_n478 = ~new_n222 & new_n345;
  assign new_n479 = id0_0_ & ~new_n478;
  assign new_n480 = ~id0_0_ & new_n478;
  assign od0_242_ = new_n479 | new_n480;
endmodule


