// Benchmark "b14" written by ABC on Wed Sep  5 10:17:20 2018

module b14 ( clock, 
    DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
    DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
    DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
    DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
    DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
    DATAI_0_,
    ADDR_REG_19_, ADDR_REG_18_, ADDR_REG_17_, ADDR_REG_16_, ADDR_REG_15_,
    ADDR_REG_14_, ADDR_REG_13_, ADDR_REG_12_, ADDR_REG_11_, ADDR_REG_10_,
    ADDR_REG_9_, ADDR_REG_8_, ADDR_REG_7_, ADDR_REG_6_, ADDR_REG_5_,
    ADDR_REG_4_, ADDR_REG_3_, ADDR_REG_2_, ADDR_REG_1_, ADDR_REG_0_,
    DATAO_REG_31_, DATAO_REG_30_, DATAO_REG_29_, DATAO_REG_28_,
    DATAO_REG_27_, DATAO_REG_26_, DATAO_REG_25_, DATAO_REG_24_,
    DATAO_REG_23_, DATAO_REG_22_, DATAO_REG_21_, DATAO_REG_20_,
    DATAO_REG_19_, DATAO_REG_18_, DATAO_REG_17_, DATAO_REG_16_,
    DATAO_REG_15_, DATAO_REG_14_, DATAO_REG_13_, DATAO_REG_12_,
    DATAO_REG_11_, DATAO_REG_10_, DATAO_REG_9_, DATAO_REG_8_, DATAO_REG_7_,
    DATAO_REG_6_, DATAO_REG_5_, DATAO_REG_4_, DATAO_REG_3_, DATAO_REG_2_,
    DATAO_REG_1_, DATAO_REG_0_, RD_REG, WR_REG  );
  input  clock;
  input  DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_,
    DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_,
    DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_,
    DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_,
    DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_,
    DATAI_1_, DATAI_0_;
  output ADDR_REG_19_, ADDR_REG_18_, ADDR_REG_17_, ADDR_REG_16_, ADDR_REG_15_,
    ADDR_REG_14_, ADDR_REG_13_, ADDR_REG_12_, ADDR_REG_11_, ADDR_REG_10_,
    ADDR_REG_9_, ADDR_REG_8_, ADDR_REG_7_, ADDR_REG_6_, ADDR_REG_5_,
    ADDR_REG_4_, ADDR_REG_3_, ADDR_REG_2_, ADDR_REG_1_, ADDR_REG_0_,
    DATAO_REG_31_, DATAO_REG_30_, DATAO_REG_29_, DATAO_REG_28_,
    DATAO_REG_27_, DATAO_REG_26_, DATAO_REG_25_, DATAO_REG_24_,
    DATAO_REG_23_, DATAO_REG_22_, DATAO_REG_21_, DATAO_REG_20_,
    DATAO_REG_19_, DATAO_REG_18_, DATAO_REG_17_, DATAO_REG_16_,
    DATAO_REG_15_, DATAO_REG_14_, DATAO_REG_13_, DATAO_REG_12_,
    DATAO_REG_11_, DATAO_REG_10_, DATAO_REG_9_, DATAO_REG_8_, DATAO_REG_7_,
    DATAO_REG_6_, DATAO_REG_5_, DATAO_REG_4_, DATAO_REG_3_, DATAO_REG_2_,
    DATAO_REG_1_, DATAO_REG_0_, RD_REG, WR_REG;
  reg IR_REG_0_, IR_REG_1_, IR_REG_2_, IR_REG_3_, IR_REG_4_, IR_REG_5_,
    IR_REG_6_, IR_REG_7_, IR_REG_8_, IR_REG_9_, IR_REG_10_, IR_REG_11_,
    IR_REG_12_, IR_REG_13_, IR_REG_14_, IR_REG_15_, IR_REG_16_, IR_REG_17_,
    IR_REG_18_, IR_REG_19_, IR_REG_20_, IR_REG_21_, IR_REG_22_, IR_REG_23_,
    IR_REG_24_, IR_REG_25_, IR_REG_26_, IR_REG_27_, IR_REG_28_, IR_REG_29_,
    IR_REG_30_, IR_REG_31_, D_REG_0_, D_REG_1_, D_REG_2_, D_REG_3_,
    D_REG_4_, D_REG_5_, D_REG_6_, D_REG_7_, D_REG_8_, D_REG_9_, D_REG_10_,
    D_REG_11_, D_REG_12_, D_REG_13_, D_REG_14_, D_REG_15_, D_REG_16_,
    D_REG_17_, D_REG_18_, D_REG_19_, D_REG_20_, D_REG_21_, D_REG_22_,
    D_REG_23_, D_REG_24_, D_REG_25_, D_REG_26_, D_REG_27_, D_REG_28_,
    D_REG_29_, D_REG_30_, D_REG_31_, REG0_REG_0_, REG0_REG_1_, REG0_REG_2_,
    REG0_REG_3_, REG0_REG_4_, REG0_REG_5_, REG0_REG_6_, REG0_REG_7_,
    REG0_REG_8_, REG0_REG_9_, REG0_REG_10_, REG0_REG_11_, REG0_REG_12_,
    REG0_REG_13_, REG0_REG_14_, REG0_REG_15_, REG0_REG_16_, REG0_REG_17_,
    REG0_REG_18_, REG0_REG_19_, REG0_REG_20_, REG0_REG_21_, REG0_REG_22_,
    REG0_REG_23_, REG0_REG_24_, REG0_REG_25_, REG0_REG_26_, REG0_REG_27_,
    REG0_REG_28_, REG0_REG_29_, REG0_REG_30_, REG0_REG_31_, REG1_REG_0_,
    REG1_REG_1_, REG1_REG_2_, REG1_REG_3_, REG1_REG_4_, REG1_REG_5_,
    REG1_REG_6_, REG1_REG_7_, REG1_REG_8_, REG1_REG_9_, REG1_REG_10_,
    REG1_REG_11_, REG1_REG_12_, REG1_REG_13_, REG1_REG_14_, REG1_REG_15_,
    REG1_REG_16_, REG1_REG_17_, REG1_REG_18_, REG1_REG_19_, REG1_REG_20_,
    REG1_REG_21_, REG1_REG_22_, REG1_REG_23_, REG1_REG_24_, REG1_REG_25_,
    REG1_REG_26_, REG1_REG_27_, REG1_REG_28_, REG1_REG_29_, REG1_REG_30_,
    REG1_REG_31_, REG2_REG_0_, REG2_REG_1_, REG2_REG_2_, REG2_REG_3_,
    REG2_REG_4_, REG2_REG_5_, REG2_REG_6_, REG2_REG_7_, REG2_REG_8_,
    REG2_REG_9_, REG2_REG_10_, REG2_REG_11_, REG2_REG_12_, REG2_REG_13_,
    REG2_REG_14_, REG2_REG_15_, REG2_REG_16_, REG2_REG_17_, REG2_REG_18_,
    REG2_REG_19_, REG2_REG_20_, REG2_REG_21_, REG2_REG_22_, REG2_REG_23_,
    REG2_REG_24_, REG2_REG_25_, REG2_REG_26_, REG2_REG_27_, REG2_REG_28_,
    REG2_REG_29_, REG2_REG_30_, REG2_REG_31_, ADDR_REG_19_, ADDR_REG_18_,
    ADDR_REG_17_, ADDR_REG_16_, ADDR_REG_15_, ADDR_REG_14_, ADDR_REG_13_,
    ADDR_REG_12_, ADDR_REG_11_, ADDR_REG_10_, ADDR_REG_9_, ADDR_REG_8_,
    ADDR_REG_7_, ADDR_REG_6_, ADDR_REG_5_, ADDR_REG_4_, ADDR_REG_3_,
    ADDR_REG_2_, ADDR_REG_1_, ADDR_REG_0_, DATAO_REG_0_, DATAO_REG_1_,
    DATAO_REG_2_, DATAO_REG_3_, DATAO_REG_4_, DATAO_REG_5_, DATAO_REG_6_,
    DATAO_REG_7_, DATAO_REG_8_, DATAO_REG_9_, DATAO_REG_10_, DATAO_REG_11_,
    DATAO_REG_12_, DATAO_REG_13_, DATAO_REG_14_, DATAO_REG_15_,
    DATAO_REG_16_, DATAO_REG_17_, DATAO_REG_18_, DATAO_REG_19_,
    DATAO_REG_20_, DATAO_REG_21_, DATAO_REG_22_, DATAO_REG_23_,
    DATAO_REG_24_, DATAO_REG_25_, DATAO_REG_26_, DATAO_REG_27_,
    DATAO_REG_28_, DATAO_REG_29_, DATAO_REG_30_, DATAO_REG_31_, B_REG,
    REG3_REG_15_, REG3_REG_26_, REG3_REG_6_, REG3_REG_18_, REG3_REG_2_,
    REG3_REG_11_, REG3_REG_22_, REG3_REG_13_, REG3_REG_20_, REG3_REG_0_,
    REG3_REG_9_, REG3_REG_4_, REG3_REG_24_, REG3_REG_17_, REG3_REG_5_,
    REG3_REG_16_, REG3_REG_25_, REG3_REG_12_, REG3_REG_21_, REG3_REG_1_,
    REG3_REG_8_, REG3_REG_28_, REG3_REG_19_, REG3_REG_3_, REG3_REG_10_,
    REG3_REG_23_, REG3_REG_14_, REG3_REG_27_, REG3_REG_7_, STATE_REG,
    RD_REG, WR_REG;
  wire n822, n823, n824_1, n825, n826, n827, n829_1, n830, n831, n832, n833,
    n834_1, n835, n837, n838, n839_1, n840, n841, n842, n843, n844_1, n846,
    n847, n848, n849_1, n850, n851, n852, n854_1, n855, n856, n857, n858,
    n859_1, n860, n862, n863, n864_1, n865, n866, n867, n868, n869_1, n870,
    n871, n872, n874_1, n875, n876, n877, n878, n879_1, n880, n882, n883,
    n884_1, n885, n886, n887, n888, n889_1, n891, n892, n893, n894_1, n895,
    n896, n897, n899_1, n900, n901, n902, n903, n904_1, n905, n906, n907,
    n909_1, n910, n911, n912, n913, n914_1, n915, n917, n918, n919_1, n920,
    n921, n922, n923, n924_1, n926, n927, n928, n929_1, n930, n931, n932,
    n934_1, n935, n936, n937, n938, n939_1, n940, n941, n942, n943, n944_1,
    n945, n946, n947, n948, n949_1, n951, n952, n953, n954_1, n955, n956,
    n957, n959_1, n960, n961, n962, n963, n964_1, n965, n966, n968, n969_1,
    n970, n971, n972, n973, n974_1, n976, n977, n978_1, n979, n980, n981,
    n982_1, n983, n984, n986_1, n987, n988, n989, n990_1, n991, n992,
    n994_1, n995, n996, n997, n998_1, n999, n1000, n1001, n1003, n1004,
    n1005, n1006_1, n1007, n1008, n1009, n1011, n1012, n1013, n1014_1,
    n1015, n1016, n1017, n1018_1, n1020, n1021, n1022_1, n1023, n1024,
    n1025, n1026_1, n1028, n1029, n1030_1, n1031, n1032, n1033, n1034_1,
    n1036, n1037, n1038_1, n1039, n1040, n1041, n1042_1, n1043, n1044,
    n1045, n1046_1, n1047, n1048, n1049, n1050_1, n1051, n1052, n1054_1,
    n1055, n1056, n1057, n1058_1, n1059, n1060, n1061, n1063, n1064, n1065,
    n1066_1, n1067, n1068, n1069, n1071, n1072, n1073, n1074_1, n1075,
    n1076, n1077, n1079, n1080, n1081, n1082_1, n1083, n1084, n1085,
    n1086_1, n1087, n1088, n1089, n1090_1, n1091, n1093, n1094_1, n1095,
    n1096, n1097, n1098_1, n1099, n1100, n1101, n1103, n1104, n1105,
    n1106_1, n1107, n1108, n1109, n1111, n1112, n1113, n1114_1, n1115,
    n1116, n1117, n1119, n1120, n1121, n1122_1, n1123, n1124, n1125,
    n1126_1, n1127, n1128, n1129, n1130_1, n1131, n1132, n1133, n1134_1,
    n1135, n1136, n1137, n1138_1, n1139, n1140, n1141, n1142_1, n1143,
    n1144, n1146_1, n1147, n1148, n1180, n1181, n1182_1, n1183, n1184,
    n1185, n1186, n1187_1, n1188, n1189, n1190, n1191, n1192_1, n1193,
    n1194, n1195, n1196, n1197_1, n1198, n1199, n1200, n1201, n1202_1,
    n1203, n1204, n1205, n1206, n1207_1, n1208, n1209, n1210, n1211,
    n1212_1, n1213, n1214, n1215, n1216, n1217_1, n1218, n1219, n1220,
    n1221, n1222_1, n1223, n1224, n1225, n1226, n1227_1, n1228, n1229,
    n1230, n1231, n1232_1, n1233, n1234, n1235, n1236, n1237_1, n1238,
    n1239, n1240, n1241, n1242_1, n1243, n1244, n1245, n1246, n1247_1,
    n1248, n1249, n1250, n1251, n1252_1, n1253, n1254, n1255, n1256,
    n1257_1, n1258, n1259, n1260, n1261, n1262_1, n1263, n1264, n1265,
    n1266, n1267_1, n1268, n1269, n1270, n1271, n1272_1, n1273, n1274,
    n1275, n1276, n1277_1, n1278, n1279, n1280, n1281, n1282_1, n1283,
    n1284, n1285, n1286, n1287_1, n1288, n1289, n1290, n1291, n1292_1,
    n1293, n1294, n1295, n1296, n1297_1, n1298, n1299, n1300, n1301,
    n1302_1, n1303, n1304, n1305, n1306, n1307_1, n1308, n1309, n1310,
    n1311, n1312_1, n1313, n1314, n1315, n1316, n1317_1, n1318, n1319,
    n1320, n1321, n1322_1, n1323, n1324, n1325, n1326, n1327_1, n1328,
    n1329, n1330, n1331, n1332_1, n1333, n1334, n1335, n1336, n1337_1,
    n1338, n1339, n1340, n1341_1, n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
    n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1409,
    n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
    n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1536, n1537, n1538, n1539, n1540, n1541,
    n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
    n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
    n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
    n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
    n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
    n1602, n1603, n1604, n1605, n1607, n1608, n1609, n1610, n1611, n1612,
    n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
    n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
    n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
    n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
    n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
    n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1672, n1673,
    n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1753, n1754,
    n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
    n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
    n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
    n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1825,
    n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
    n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
    n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
    n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
    n1886, n1887, n1888, n1889, n1890, n1891, n1893, n1894, n1895, n1896,
    n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
    n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
    n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
    n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
    n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
    n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
    n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1966, n1967,
    n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
    n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
    n2028, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
    n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
    n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
    n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
    n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
    n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
    n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
    n2099, n2100, n2101, n2102, n2103, n2104, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
    n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
    n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
    n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
    n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
    n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
    n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
    n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
    n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
    n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
    n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
    n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
    n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
    n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
    n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
    n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
    n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
    n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
    n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
    n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
    n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
    n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
    n2444, n2445, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
    n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
    n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
    n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
    n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
    n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
    n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
    n2515, n2516, n2517, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
    n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
    n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
    n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
    n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
    n2586, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
    n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
    n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
    n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
    n2647, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
    n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
    n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
    n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2708,
    n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
    n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
    n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
    n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
    n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
    n2769, n2770, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
    n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
    n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
    n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
    n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
    n2840, n2841, n2842, n2843, n2845, n2846, n2847, n2848, n2849, n2850,
    n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
    n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
    n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
    n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
    n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
    n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
    n2931, n2932, n2933, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
    n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
    n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
    n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
    n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
    n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
    n3002, n3003, n3004, n3005, n3007, n3008, n3009, n3010, n3011, n3012,
    n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
    n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
    n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
    n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
    n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
    n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
    n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
    n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
    n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
    n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
    n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
    n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
    n3144, n3145, n3146, n3147, n3148, n3150, n3151, n3152, n3153, n3154,
    n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
    n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
    n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
    n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
    n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
    n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
    n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
    n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
    n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
    n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
    n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
    n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
    n3306, n3307, n3308, n3309, n3310, n3311, n3313, n3314, n3315, n3316,
    n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
    n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
    n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
    n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
    n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
    n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
    n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
    n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
    n3408, n3409, n3410, n3411, n3413, n3414, n3415, n3416, n3417, n3418,
    n3419, n3420, n3421, n3422, n3423, n3424, n3426, n3427, n3428, n3429,
    n3431, n3432, n3434, n3435, n3437, n3438, n3440, n3441, n3443, n3444,
    n3446, n3447, n3449, n3450, n3452, n3453, n3455, n3456, n3458, n3459,
    n3461, n3462, n3464, n3465, n3467, n3468, n3470, n3471, n3473, n3474,
    n3476, n3477, n3479, n3480, n3482, n3483, n3485, n3486, n3488, n3489,
    n3491, n3492, n3494, n3495, n3497, n3498, n3500, n3501, n3503, n3504,
    n3506, n3507, n3509, n3510, n3512, n3513, n3515, n3516, n3518, n3519,
    n3521, n3522, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
    n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
    n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3552,
    n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
    n3563, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
    n3574, n3575, n3576, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3591, n3592, n3593, n3594, n3595,
    n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3604, n3605, n3606,
    n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3617,
    n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
    n3628, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
    n3650, n3651, n3652, n3653, n3654, n3656, n3657, n3658, n3659, n3660,
    n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3669, n3670, n3671,
    n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3682,
    n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
    n3693, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
    n3704, n3705, n3706, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
    n3715, n3716, n3717, n3718, n3719, n3721, n3722, n3723, n3724, n3725,
    n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3734, n3735, n3736,
    n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3747,
    n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
    n3758, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
    n3769, n3770, n3771, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
    n3780, n3781, n3782, n3783, n3784, n3786, n3787, n3788, n3789, n3790,
    n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3812,
    n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
    n3823, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
    n3834, n3835, n3836, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
    n3845, n3846, n3847, n3848, n3849, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3864, n3865, n3866,
    n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3877,
    n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
    n3888, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
    n3899, n3900, n3901, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3916, n3917, n3918, n3919, n3920,
    n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3930, n3931,
    n3932, n3933, n3934, n3935, n3937, n3938, n3939, n3940, n3941, n3943,
    n3944, n3945, n3946, n3947, n3949, n3950, n3951, n3952, n3953, n3954,
    n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
    n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
    n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
    n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
    n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
    n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
    n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
    n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
    n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
    n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
    n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
    n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
    n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
    n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
    n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
    n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
    n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
    n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
    n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
    n4145, n4146, n4147, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
    n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
    n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
    n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
    n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
    n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4205, n4206, n4207,
    n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
    n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
    n4228, n4229, n4230, n4231, n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
    n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4259,
    n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
    n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
    n4280, n4281, n4282, n4283, n4285, n4286, n4287, n4288, n4289, n4290,
    n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
    n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4311,
    n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
    n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
    n4332, n4333, n4334, n4335, n4336, n4337, n4339, n4340, n4341, n4342,
    n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
    n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
    n4363, n4364, n4365, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
    n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
    n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4393, n4394,
    n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
    n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
    n4415, n4416, n4417, n4418, n4419, n4421, n4422, n4423, n4424, n4425,
    n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
    n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
    n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
    n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
    n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4475, n4476, n4477,
    n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
    n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
    n4498, n4499, n4500, n4501, n4503, n4504, n4505, n4506, n4507, n4508,
    n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
    n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4529,
    n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
    n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
    n4550, n4551, n4552, n4553, n4555, n4556, n4557, n4558, n4559, n4560,
    n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
    n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
    n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
    n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
    n4601, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
    n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
    n4622, n4623, n4624, n4625, n4626, n4627, n4629, n4630, n4631, n4632,
    n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
    n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
    n4653, n4654, n4655, n4656, n4658, n4659, n4660, n4661, n4662, n4663,
    n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
    n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
    n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4692, n4693, n4694,
    n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
    n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4714, n4715,
    n4717, n4718, n4720, n4721, n4723, n4724, n4726, n4727, n4729, n4730,
    n4732, n4733, n4735, n4736, n4738, n4739, n4741, n4742, n4744, n4745,
    n4747, n4748, n4750, n4751, n4753, n4754, n4756, n4757, n4759, n4760,
    n4762, n4763, n4765, n4766, n4768, n4769, n4771, n4772, n4774, n4775,
    n4777, n4778, n4780, n4781, n4783, n4784, n4786, n4787, n4789, n4790,
    n4792, n4793, n4795, n4796, n4798, n4799, n4801, n4802, n4804, n4805,
    n4807, n4808, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
    n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
    n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
    n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
    n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
    n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
    n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
    n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
    n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
    n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
    n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
    n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
    n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
    n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
    n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
    n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
    n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
    n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
    n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
    n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
    n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
    n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
    n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
    n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
    n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
    n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
    n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
    n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
    n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
    n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
    n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
    n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
    n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
    n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
    n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
    n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
    n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
    n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
    n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
    n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
    n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
    n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
    n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
    n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
    n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
    n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
    n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
    n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
    n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
    n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
    n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
    n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
    n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
    n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
    n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
    n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
    n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
    n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
    n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
    n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
    n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
    n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
    n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
    n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
    n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
    n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
    n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
    n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
    n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
    n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
    n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
    n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
    n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
    n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
    n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
    n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
    n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
    n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
    n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
    n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
    n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
    n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
    n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
    n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
    n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
    n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
    n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
    n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
    n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
    n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
    n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
    n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
    n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
    n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
    n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
    n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
    n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
    n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
    n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
    n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
    n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
    n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
    n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
    n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
    n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
    n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
    n5868, n5869, n5870, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
    n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
    n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
    n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
    n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
    n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
    n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
    n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
    n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
    n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
    n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
    n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
    n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
    n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
    n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
    n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
    n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
    n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
    n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
    n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
    n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
    n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
    n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
    n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
    n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
    n6119, n6120, n6121, n6122, n6124, n6125, n6126, n6127, n6128, n6129,
    n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
    n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
    n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
    n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
    n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
    n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
    n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
    n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
    n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
    n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
    n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
    n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
    n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
    n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
    n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
    n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
    n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
    n6300, n6301, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
    n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
    n6321, n6322, n6323, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
    n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
    n6342, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
    n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
    n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
    n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
    n6384, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
    n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
    n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
    n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
    n6426, n6427, n6428, n6429, n6431, n6432, n6433, n6434, n6435, n6436,
    n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
    n6447, n6448, n6449, n6450, n6451, n6452, n6454, n6455, n6456, n6457,
    n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6466, n6467, n6468,
    n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
    n6479, n6480, n6481, n6482, n6483, n6485, n6486, n6487, n6488, n6489,
    n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
    n6500, n6501, n6502, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
    n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
    n6521, n6522, n6523, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
    n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
    n6542, n6543, n6544, n6545, n6546, n6547, n6549, n6550, n6551, n6552,
    n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
    n6563, n6564, n6565, n6566, n6568, n6569, n6570, n6571, n6572, n6573,
    n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
    n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
    n6605, n6606, n6607, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
    n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
    n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
    n6647, n6648, n6649, n6650, n6651, n6653, n6654, n6655, n6656, n6657,
    n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
    n6668, n6669, n6670, n6671, n6673, n6674, n6675, n6676, n6677, n6678,
    n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
    n6689, n6690, n6691, n6692, n6694, n6695, n6696, n6697, n6698, n6699,
    n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
    n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
    n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
    n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
    n6740, n6741, n6742, n6743, n6744, n6746, n6747, n6748, n6749, n6750,
    n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
    n6761, n6762, n6763, n6764, n6766, n6767, n6768, n6769, n6770, n6771,
    n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
    n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6790, n6791, n6792,
    n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
    n6803, n6804, n6805, n6806, n6807, n6809, n6810, n6811, n6812, n6813,
    n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
    n6824, n6825, n6826, n6827, n6829, n6830, n6831, n6832, n6833, n6834,
    n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
    n6845, n6846, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
    n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
    n6866, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
    n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
    n6887, n6888, n6889, n6890, n174, n179, n184, n189, n194, n199, n204,
    n209, n214, n219, n224, n229, n234, n239, n244, n249, n254, n259, n264,
    n269, n274, n279, n284, n289, n294, n299, n304, n309, n314, n319, n324,
    n329, n334, n339, n344, n349, n354, n359, n364, n369, n374, n379, n384,
    n389, n394, n399, n404, n409, n414, n419, n424, n429, n434, n439, n444,
    n449, n454, n459, n464, n469, n474, n479, n484, n489, n494, n499, n504,
    n509, n514, n519, n524, n529, n534, n539, n544, n549, n554, n559, n564,
    n569, n574, n579, n584, n589, n594, n599, n604, n609, n614, n619, n624,
    n629, n634, n639, n644, n649, n654, n659, n664, n669, n674, n679, n684,
    n689, n694, n699, n704, n709, n714, n719, n724, n729, n734, n739, n744,
    n749, n754, n759, n764, n769, n774, n779, n784, n789, n794, n799, n804,
    n809, n814, n819, n824, n829, n834, n839, n844, n849, n854, n859, n864,
    n869, n874, n879, n884, n889, n894, n899, n904, n909, n914, n919, n924,
    n929, n934, n939, n944, n949, n954, n959, n964, n969, n974, n978, n982,
    n986, n990, n994, n998, n1002, n1006, n1010, n1014, n1018, n1022,
    n1026, n1030, n1034, n1038, n1042, n1046, n1050, n1054, n1058, n1062,
    n1066, n1070, n1074, n1078, n1082, n1086, n1090, n1094, n1098, n1102,
    n1106, n1110, n1114, n1118, n1122, n1126, n1130, n1134, n1138, n1142,
    n1146, n1150, n1154, n1158, n1162, n1166, n1170, n1174, n1178, n1182,
    n1187, n1192, n1197, n1202, n1207, n1212, n1217, n1222, n1227, n1232,
    n1237, n1242, n1247, n1252, n1257, n1262, n1267, n1272, n1277, n1282,
    n1287, n1292, n1297, n1302, n1307, n1312, n1317, n1322, n1327, n1332,
    n1337, n1341;
  assign n822 = ~IR_REG_31_ & STATE_REG;
  assign n823 = IR_REG_0_ & n822;
  assign n824_1 = DATAI_0_ & ~STATE_REG;
  assign n825 = ~n823 & ~n824_1;
  assign n826 = STATE_REG & ~n822;
  assign n827 = IR_REG_0_ & n826;
  assign n174 = ~n825 | n827;
  assign n829_1 = IR_REG_1_ & n822;
  assign n830 = DATAI_1_ & ~STATE_REG;
  assign n831 = ~n829_1 & ~n830;
  assign n832 = IR_REG_0_ & ~IR_REG_1_;
  assign n833 = ~IR_REG_0_ & IR_REG_1_;
  assign n834_1 = ~n832 & ~n833;
  assign n835 = n826 & ~n834_1;
  assign n179 = ~n831 | n835;
  assign n837 = IR_REG_2_ & n822;
  assign n838 = DATAI_2_ & ~STATE_REG;
  assign n839_1 = ~n837 & ~n838;
  assign n840 = ~IR_REG_0_ & ~IR_REG_1_;
  assign n841 = IR_REG_2_ & ~n840;
  assign n842 = ~IR_REG_2_ & n840;
  assign n843 = ~n841 & ~n842;
  assign n844_1 = n826 & n843;
  assign n184 = ~n839_1 | n844_1;
  assign n846 = IR_REG_3_ & n822;
  assign n847 = DATAI_3_ & ~STATE_REG;
  assign n848 = ~n846 & ~n847;
  assign n849_1 = IR_REG_3_ & ~n842;
  assign n850 = ~IR_REG_3_ & n842;
  assign n851 = ~n849_1 & ~n850;
  assign n852 = n826 & n851;
  assign n189 = ~n848 | n852;
  assign n854_1 = IR_REG_4_ & n822;
  assign n855 = DATAI_4_ & ~STATE_REG;
  assign n856 = ~n854_1 & ~n855;
  assign n857 = ~IR_REG_4_ & n850;
  assign n858 = IR_REG_4_ & ~n850;
  assign n859_1 = ~n857 & ~n858;
  assign n860 = n826 & n859_1;
  assign n194 = ~n856 | n860;
  assign n862 = IR_REG_5_ & n822;
  assign n863 = DATAI_5_ & ~STATE_REG;
  assign n864_1 = ~n862 & ~n863;
  assign n865 = IR_REG_5_ & ~n857;
  assign n866 = ~IR_REG_3_ & ~IR_REG_5_;
  assign n867 = ~IR_REG_4_ & n866;
  assign n868 = ~IR_REG_1_ & ~IR_REG_2_;
  assign n869_1 = ~IR_REG_0_ & n868;
  assign n870 = n867 & n869_1;
  assign n871 = ~n865 & ~n870;
  assign n872 = n826 & n871;
  assign n199 = ~n864_1 | n872;
  assign n874_1 = IR_REG_6_ & n822;
  assign n875 = DATAI_6_ & ~STATE_REG;
  assign n876 = ~n874_1 & ~n875;
  assign n877 = IR_REG_6_ & ~n870;
  assign n878 = ~IR_REG_6_ & n870;
  assign n879_1 = ~n877 & ~n878;
  assign n880 = n826 & n879_1;
  assign n204 = ~n876 | n880;
  assign n882 = IR_REG_7_ & n822;
  assign n883 = DATAI_7_ & ~STATE_REG;
  assign n884_1 = ~n882 & ~n883;
  assign n885 = IR_REG_7_ & ~n878;
  assign n886 = ~IR_REG_6_ & ~IR_REG_7_;
  assign n887 = n870 & n886;
  assign n888 = ~n885 & ~n887;
  assign n889_1 = n826 & n888;
  assign n209 = ~n884_1 | n889_1;
  assign n891 = IR_REG_8_ & n822;
  assign n892 = DATAI_8_ & ~STATE_REG;
  assign n893 = ~n891 & ~n892;
  assign n894_1 = ~IR_REG_8_ & n887;
  assign n895 = IR_REG_8_ & ~n887;
  assign n896 = ~n894_1 & ~n895;
  assign n897 = n826 & n896;
  assign n214 = ~n893 | n897;
  assign n899_1 = IR_REG_9_ & n822;
  assign n900 = DATAI_9_ & ~STATE_REG;
  assign n901 = ~n899_1 & ~n900;
  assign n902 = IR_REG_9_ & ~n894_1;
  assign n903 = ~IR_REG_8_ & n886;
  assign n904_1 = ~IR_REG_9_ & n903;
  assign n905 = n870 & n904_1;
  assign n906 = ~n902 & ~n905;
  assign n907 = n826 & n906;
  assign n219 = ~n901 | n907;
  assign n909_1 = IR_REG_10_ & n822;
  assign n910 = DATAI_10_ & ~STATE_REG;
  assign n911 = ~n909_1 & ~n910;
  assign n912 = IR_REG_10_ & ~n905;
  assign n913 = ~IR_REG_10_ & n905;
  assign n914_1 = ~n912 & ~n913;
  assign n915 = n826 & n914_1;
  assign n224 = ~n911 | n915;
  assign n917 = IR_REG_11_ & n822;
  assign n918 = DATAI_11_ & ~STATE_REG;
  assign n919_1 = ~n917 & ~n918;
  assign n920 = IR_REG_11_ & ~n913;
  assign n921 = ~IR_REG_10_ & ~IR_REG_11_;
  assign n922 = n905 & n921;
  assign n923 = ~n920 & ~n922;
  assign n924_1 = n826 & n923;
  assign n229 = ~n919_1 | n924_1;
  assign n926 = IR_REG_12_ & n822;
  assign n927 = DATAI_12_ & ~STATE_REG;
  assign n928 = ~n926 & ~n927;
  assign n929_1 = ~IR_REG_12_ & n922;
  assign n930 = IR_REG_12_ & ~n922;
  assign n931 = ~n929_1 & ~n930;
  assign n932 = n826 & n931;
  assign n234 = ~n928 | n932;
  assign n934_1 = IR_REG_13_ & n822;
  assign n935 = DATAI_13_ & ~STATE_REG;
  assign n936 = ~n934_1 & ~n935;
  assign n937 = IR_REG_13_ & ~n929_1;
  assign n938 = ~IR_REG_7_ & ~IR_REG_9_;
  assign n939_1 = ~IR_REG_8_ & n938;
  assign n940 = ~IR_REG_3_ & ~IR_REG_4_;
  assign n941 = ~IR_REG_5_ & n940;
  assign n942 = ~IR_REG_6_ & n941;
  assign n943 = ~IR_REG_12_ & n921;
  assign n944_1 = ~IR_REG_13_ & n943;
  assign n945 = n939_1 & n942;
  assign n946 = n869_1 & n945;
  assign n947 = n944_1 & n946;
  assign n948 = ~n937 & ~n947;
  assign n949_1 = n826 & n948;
  assign n239 = ~n936 | n949_1;
  assign n951 = IR_REG_14_ & n822;
  assign n952 = DATAI_14_ & ~STATE_REG;
  assign n953 = ~n951 & ~n952;
  assign n954_1 = IR_REG_14_ & ~n947;
  assign n955 = ~IR_REG_14_ & n947;
  assign n956 = ~n954_1 & ~n955;
  assign n957 = n826 & n956;
  assign n244 = ~n953 | n957;
  assign n959_1 = IR_REG_15_ & n822;
  assign n960 = DATAI_15_ & ~STATE_REG;
  assign n961 = ~n959_1 & ~n960;
  assign n962 = IR_REG_15_ & ~n955;
  assign n963 = ~IR_REG_14_ & ~IR_REG_15_;
  assign n964_1 = n947 & n963;
  assign n965 = ~n962 & ~n964_1;
  assign n966 = n826 & n965;
  assign n249 = ~n961 | n966;
  assign n968 = IR_REG_16_ & n822;
  assign n969_1 = DATAI_16_ & ~STATE_REG;
  assign n970 = ~n968 & ~n969_1;
  assign n971 = ~IR_REG_16_ & n964_1;
  assign n972 = IR_REG_16_ & ~n964_1;
  assign n973 = ~n971 & ~n972;
  assign n974_1 = n826 & n973;
  assign n254 = ~n970 | n974_1;
  assign n976 = IR_REG_17_ & n822;
  assign n977 = DATAI_17_ & ~STATE_REG;
  assign n978_1 = ~n976 & ~n977;
  assign n979 = IR_REG_17_ & ~n971;
  assign n980 = ~IR_REG_16_ & n963;
  assign n981 = ~IR_REG_17_ & n980;
  assign n982_1 = n947 & n981;
  assign n983 = ~n979 & ~n982_1;
  assign n984 = n826 & n983;
  assign n259 = ~n978_1 | n984;
  assign n986_1 = IR_REG_18_ & n822;
  assign n987 = DATAI_18_ & ~STATE_REG;
  assign n988 = ~n986_1 & ~n987;
  assign n989 = IR_REG_18_ & ~n982_1;
  assign n990_1 = ~IR_REG_18_ & n982_1;
  assign n991 = ~n989 & ~n990_1;
  assign n992 = n826 & n991;
  assign n264 = ~n988 | n992;
  assign n994_1 = IR_REG_19_ & n822;
  assign n995 = DATAI_19_ & ~STATE_REG;
  assign n996 = ~n994_1 & ~n995;
  assign n997 = IR_REG_19_ & ~n990_1;
  assign n998_1 = ~IR_REG_18_ & ~IR_REG_19_;
  assign n999 = n982_1 & n998_1;
  assign n1000 = ~n997 & ~n999;
  assign n1001 = n826 & n1000;
  assign n269 = ~n996 | n1001;
  assign n1003 = IR_REG_20_ & n822;
  assign n1004 = DATAI_20_ & ~STATE_REG;
  assign n1005 = ~n1003 & ~n1004;
  assign n1006_1 = ~IR_REG_20_ & n999;
  assign n1007 = IR_REG_20_ & ~n999;
  assign n1008 = ~n1006_1 & ~n1007;
  assign n1009 = n826 & n1008;
  assign n274 = ~n1005 | n1009;
  assign n1011 = IR_REG_21_ & n822;
  assign n1012 = DATAI_21_ & ~STATE_REG;
  assign n1013 = ~n1011 & ~n1012;
  assign n1014_1 = IR_REG_21_ & ~n1006_1;
  assign n1015 = ~IR_REG_20_ & ~IR_REG_21_;
  assign n1016 = n999 & n1015;
  assign n1017 = ~n1014_1 & ~n1016;
  assign n1018_1 = n826 & n1017;
  assign n279 = ~n1013 | n1018_1;
  assign n1020 = IR_REG_22_ & n822;
  assign n1021 = DATAI_22_ & ~STATE_REG;
  assign n1022_1 = ~n1020 & ~n1021;
  assign n1023 = IR_REG_22_ & ~n1016;
  assign n1024 = ~IR_REG_22_ & n1016;
  assign n1025 = ~n1023 & ~n1024;
  assign n1026_1 = n826 & n1025;
  assign n284 = ~n1022_1 | n1026_1;
  assign n1028 = IR_REG_23_ & n822;
  assign n1029 = DATAI_23_ & ~STATE_REG;
  assign n1030_1 = ~n1028 & ~n1029;
  assign n1031 = ~IR_REG_23_ & n1024;
  assign n1032 = IR_REG_23_ & ~n1024;
  assign n1033 = ~n1031 & ~n1032;
  assign n1034_1 = n826 & n1033;
  assign n289 = ~n1030_1 | n1034_1;
  assign n1036 = IR_REG_24_ & n822;
  assign n1037 = DATAI_24_ & ~STATE_REG;
  assign n1038_1 = ~n1036 & ~n1037;
  assign n1039 = ~IR_REG_22_ & ~IR_REG_23_;
  assign n1040 = ~IR_REG_21_ & n1039;
  assign n1041 = ~IR_REG_19_ & n1040;
  assign n1042_1 = ~IR_REG_20_ & n1041;
  assign n1043 = ~IR_REG_17_ & ~IR_REG_18_;
  assign n1044 = ~IR_REG_16_ & n1043;
  assign n1045 = ~IR_REG_14_ & n1044;
  assign n1046_1 = ~IR_REG_15_ & n1045;
  assign n1047 = n1042_1 & n1046_1;
  assign n1048 = n947 & n1047;
  assign n1049 = ~IR_REG_24_ & n1048;
  assign n1050_1 = IR_REG_24_ & ~n1048;
  assign n1051 = ~n1049 & ~n1050_1;
  assign n1052 = n826 & n1051;
  assign n294 = ~n1038_1 | n1052;
  assign n1054_1 = IR_REG_25_ & n822;
  assign n1055 = DATAI_25_ & ~STATE_REG;
  assign n1056 = ~n1054_1 & ~n1055;
  assign n1057 = IR_REG_25_ & ~n1049;
  assign n1058_1 = ~IR_REG_24_ & ~IR_REG_25_;
  assign n1059 = n1048 & n1058_1;
  assign n1060 = ~n1057 & ~n1059;
  assign n1061 = n826 & n1060;
  assign n299 = ~n1056 | n1061;
  assign n1063 = IR_REG_26_ & n822;
  assign n1064 = DATAI_26_ & ~STATE_REG;
  assign n1065 = ~n1063 & ~n1064;
  assign n1066_1 = IR_REG_26_ & ~n1059;
  assign n1067 = ~IR_REG_26_ & n1059;
  assign n1068 = ~n1066_1 & ~n1067;
  assign n1069 = n826 & n1068;
  assign n304 = ~n1065 | n1069;
  assign n1071 = IR_REG_27_ & n822;
  assign n1072 = DATAI_27_ & ~STATE_REG;
  assign n1073 = ~n1071 & ~n1072;
  assign n1074_1 = ~IR_REG_27_ & n1067;
  assign n1075 = IR_REG_27_ & ~n1067;
  assign n1076 = ~n1074_1 & ~n1075;
  assign n1077 = n826 & n1076;
  assign n309 = ~n1073 | n1077;
  assign n1079 = IR_REG_28_ & n822;
  assign n1080 = DATAI_28_ & ~STATE_REG;
  assign n1081 = ~n1079 & ~n1080;
  assign n1082_1 = ~IR_REG_26_ & ~IR_REG_27_;
  assign n1083 = ~IR_REG_24_ & n1082_1;
  assign n1084 = ~IR_REG_25_ & n1083;
  assign n1085 = n1048 & n1084;
  assign n1086_1 = IR_REG_28_ & ~n1085;
  assign n1087 = n947 & n1084;
  assign n1088 = n1047 & n1087;
  assign n1089 = ~IR_REG_28_ & n1088;
  assign n1090_1 = ~n1086_1 & ~n1089;
  assign n1091 = n826 & n1090_1;
  assign n314 = ~n1081 | n1091;
  assign n1093 = IR_REG_29_ & n822;
  assign n1094_1 = DATAI_29_ & ~STATE_REG;
  assign n1095 = ~n1093 & ~n1094_1;
  assign n1096 = IR_REG_29_ & ~n1089;
  assign n1097 = ~IR_REG_28_ & ~IR_REG_29_;
  assign n1098_1 = n1087 & n1097;
  assign n1099 = n1047 & n1098_1;
  assign n1100 = ~n1096 & ~n1099;
  assign n1101 = n826 & n1100;
  assign n319 = ~n1095 | n1101;
  assign n1103 = IR_REG_30_ & n822;
  assign n1104 = DATAI_30_ & ~STATE_REG;
  assign n1105 = ~n1103 & ~n1104;
  assign n1106_1 = ~IR_REG_30_ & n1099;
  assign n1107 = IR_REG_30_ & ~n1099;
  assign n1108 = ~n1106_1 & ~n1107;
  assign n1109 = n826 & n1108;
  assign n324 = ~n1105 | n1109;
  assign n1111 = IR_REG_31_ & n822;
  assign n1112 = DATAI_31_ & ~STATE_REG;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114_1 = IR_REG_31_ & n1106_1;
  assign n1115 = ~IR_REG_31_ & ~n1106_1;
  assign n1116 = ~n1114_1 & ~n1115;
  assign n1117 = n826 & ~n1116;
  assign n329 = ~n1113 | n1117;
  assign n1119 = IR_REG_31_ & n1033;
  assign n1120 = IR_REG_23_ & ~IR_REG_31_;
  assign n1121 = ~n1119 & ~n1120;
  assign n1122_1 = IR_REG_31_ & n1060;
  assign n1123 = IR_REG_25_ & ~IR_REG_31_;
  assign n1124 = ~n1122_1 & ~n1123;
  assign n1125 = IR_REG_31_ & n1068;
  assign n1126_1 = IR_REG_26_ & ~IR_REG_31_;
  assign n1127 = ~n1125 & ~n1126_1;
  assign n1128 = IR_REG_31_ & n1051;
  assign n1129 = IR_REG_24_ & ~IR_REG_31_;
  assign n1130_1 = ~n1128 & ~n1129;
  assign n1131 = ~n1124 & ~n1127;
  assign n1132 = ~n1130_1 & n1131;
  assign n1133 = n1121 & ~n1132;
  assign n1134_1 = STATE_REG & n1133;
  assign n1135 = n1124 & ~n1127;
  assign n1136 = n1130_1 & n1135;
  assign n1137 = B_REG & n1136;
  assign n1138_1 = ~B_REG & ~n1130_1;
  assign n1139 = ~n1137 & ~n1138_1;
  assign n1140 = ~n1127 & n1139;
  assign n1141 = n1134_1 & ~n1140;
  assign n1142_1 = n1130_1 & ~n1135;
  assign n1143 = n1141 & ~n1142_1;
  assign n1144 = D_REG_0_ & ~n1141;
  assign n334 = n1143 | n1144;
  assign n1146_1 = n1124 & ~n1135;
  assign n1147 = n1141 & ~n1146_1;
  assign n1148 = D_REG_1_ & ~n1141;
  assign n339 = n1147 | n1148;
  assign n344 = D_REG_2_ & ~n1141;
  assign n349 = D_REG_3_ & ~n1141;
  assign n354 = D_REG_4_ & ~n1141;
  assign n359 = D_REG_5_ & ~n1141;
  assign n364 = D_REG_6_ & ~n1141;
  assign n369 = D_REG_7_ & ~n1141;
  assign n374 = D_REG_8_ & ~n1141;
  assign n379 = D_REG_9_ & ~n1141;
  assign n384 = D_REG_10_ & ~n1141;
  assign n389 = D_REG_11_ & ~n1141;
  assign n394 = D_REG_12_ & ~n1141;
  assign n399 = D_REG_13_ & ~n1141;
  assign n404 = D_REG_14_ & ~n1141;
  assign n409 = D_REG_15_ & ~n1141;
  assign n414 = D_REG_16_ & ~n1141;
  assign n419 = D_REG_17_ & ~n1141;
  assign n424 = D_REG_18_ & ~n1141;
  assign n429 = D_REG_19_ & ~n1141;
  assign n434 = D_REG_20_ & ~n1141;
  assign n439 = D_REG_21_ & ~n1141;
  assign n444 = D_REG_22_ & ~n1141;
  assign n449 = D_REG_23_ & ~n1141;
  assign n454 = D_REG_24_ & ~n1141;
  assign n459 = D_REG_25_ & ~n1141;
  assign n464 = D_REG_26_ & ~n1141;
  assign n469 = D_REG_27_ & ~n1141;
  assign n474 = D_REG_28_ & ~n1141;
  assign n479 = D_REG_29_ & ~n1141;
  assign n484 = D_REG_30_ & ~n1141;
  assign n489 = D_REG_31_ & ~n1141;
  assign n1180 = D_REG_0_ & n1140;
  assign n1181 = n1127 & n1130_1;
  assign n1182_1 = ~n1140 & ~n1181;
  assign n1183 = ~n1180 & ~n1182_1;
  assign n1184 = n1134_1 & n1183;
  assign n1185 = ~n1140 & ~n1146_1;
  assign n1186 = D_REG_1_ & n1140;
  assign n1187_1 = ~n1185 & ~n1186;
  assign n1188 = IR_REG_31_ & n1008;
  assign n1189 = IR_REG_20_ & ~IR_REG_31_;
  assign n1190 = ~n1188 & ~n1189;
  assign n1191 = IR_REG_31_ & n1000;
  assign n1192_1 = IR_REG_19_ & ~IR_REG_31_;
  assign n1193 = ~n1191 & ~n1192_1;
  assign n1194 = n1190 & n1193;
  assign n1195 = IR_REG_31_ & n1017;
  assign n1196 = IR_REG_21_ & ~IR_REG_31_;
  assign n1197_1 = ~n1195 & ~n1196;
  assign n1198 = ~n1190 & n1197_1;
  assign n1199 = IR_REG_31_ & n1025;
  assign n1200 = IR_REG_22_ & ~IR_REG_31_;
  assign n1201 = ~n1199 & ~n1200;
  assign n1202_1 = ~n1197_1 & n1201;
  assign n1203 = n1197_1 & ~n1201;
  assign n1204 = ~n1194 & ~n1198;
  assign n1205 = ~n1202_1 & n1204;
  assign n1206 = ~n1203 & n1205;
  assign n1207_1 = n1187_1 & ~n1206;
  assign n1208 = D_REG_8_ & n1140;
  assign n1209 = D_REG_7_ & n1140;
  assign n1210 = D_REG_9_ & n1140;
  assign n1211 = ~n1208 & ~n1209;
  assign n1212_1 = ~n1210 & n1211;
  assign n1213 = D_REG_6_ & n1140;
  assign n1214 = D_REG_5_ & n1140;
  assign n1215 = D_REG_4_ & n1140;
  assign n1216 = D_REG_3_ & n1140;
  assign n1217_1 = ~n1213 & ~n1214;
  assign n1218 = ~n1215 & n1217_1;
  assign n1219 = ~n1216 & n1218;
  assign n1220 = D_REG_31_ & n1140;
  assign n1221 = D_REG_30_ & n1140;
  assign n1222_1 = D_REG_2_ & n1140;
  assign n1223 = D_REG_29_ & n1140;
  assign n1224 = ~n1220 & ~n1221;
  assign n1225 = ~n1222_1 & n1224;
  assign n1226 = ~n1223 & n1225;
  assign n1227_1 = D_REG_28_ & n1140;
  assign n1228 = D_REG_27_ & n1140;
  assign n1229 = D_REG_26_ & n1140;
  assign n1230 = D_REG_25_ & n1140;
  assign n1231 = ~n1227_1 & ~n1228;
  assign n1232_1 = ~n1229 & n1231;
  assign n1233 = ~n1230 & n1232_1;
  assign n1234 = n1212_1 & n1219;
  assign n1235 = n1226 & n1234;
  assign n1236 = n1233 & n1235;
  assign n1237_1 = D_REG_23_ & n1140;
  assign n1238 = D_REG_22_ & n1140;
  assign n1239 = D_REG_24_ & n1140;
  assign n1240 = ~n1237_1 & ~n1238;
  assign n1241 = ~n1239 & n1240;
  assign n1242_1 = D_REG_21_ & n1140;
  assign n1243 = D_REG_20_ & n1140;
  assign n1244 = D_REG_19_ & n1140;
  assign n1245 = D_REG_18_ & n1140;
  assign n1246 = ~n1242_1 & ~n1243;
  assign n1247_1 = ~n1244 & n1246;
  assign n1248 = ~n1245 & n1247_1;
  assign n1249 = D_REG_17_ & n1140;
  assign n1250 = D_REG_16_ & n1140;
  assign n1251 = D_REG_15_ & n1140;
  assign n1252_1 = D_REG_14_ & n1140;
  assign n1253 = ~n1249 & ~n1250;
  assign n1254 = ~n1251 & n1253;
  assign n1255 = ~n1252_1 & n1254;
  assign n1256 = D_REG_13_ & n1140;
  assign n1257_1 = D_REG_12_ & n1140;
  assign n1258 = D_REG_11_ & n1140;
  assign n1259 = D_REG_10_ & n1140;
  assign n1260 = ~n1256 & ~n1257_1;
  assign n1261 = ~n1258 & n1260;
  assign n1262_1 = ~n1259 & n1261;
  assign n1263 = n1241 & n1248;
  assign n1264 = n1255 & n1263;
  assign n1265 = n1262_1 & n1264;
  assign n1266 = n1236 & n1265;
  assign n1267_1 = n1207_1 & n1266;
  assign n1268 = n1184 & n1267_1;
  assign n1269 = IR_REG_31_ & n1076;
  assign n1270 = IR_REG_27_ & ~IR_REG_31_;
  assign n1271 = ~n1269 & ~n1270;
  assign n1272_1 = IR_REG_31_ & n1090_1;
  assign n1273 = IR_REG_28_ & ~IR_REG_31_;
  assign n1274 = ~n1272_1 & ~n1273;
  assign n1275 = n1271 & n1274;
  assign n1276 = IR_REG_0_ & IR_REG_31_;
  assign n1277_1 = IR_REG_0_ & ~IR_REG_31_;
  assign n1278 = ~n1276 & ~n1277_1;
  assign n1279 = n1275 & ~n1278;
  assign n1280 = DATAI_0_ & ~n1275;
  assign n1281 = ~n1279 & ~n1280;
  assign n1282_1 = n1198 & n1201;
  assign n1283 = ~n1281 & n1282_1;
  assign n1284 = ~n1197_1 & ~n1201;
  assign n1285 = n1274 & n1284;
  assign n1286 = IR_REG_31_ & n1108;
  assign n1287_1 = IR_REG_30_ & ~IR_REG_31_;
  assign n1288 = ~n1286 & ~n1287_1;
  assign n1289 = IR_REG_31_ & n1100;
  assign n1290 = IR_REG_29_ & ~IR_REG_31_;
  assign n1291 = ~n1289 & ~n1290;
  assign n1292_1 = ~n1288 & ~n1291;
  assign n1293 = REG3_REG_1_ & n1292_1;
  assign n1294 = n1288 & n1291;
  assign n1295 = REG0_REG_1_ & n1294;
  assign n1296 = n1288 & ~n1291;
  assign n1297_1 = REG1_REG_1_ & n1296;
  assign n1298 = ~n1288 & n1291;
  assign n1299 = REG2_REG_1_ & n1298;
  assign n1300 = ~n1293 & ~n1295;
  assign n1301 = ~n1297_1 & n1300;
  assign n1302_1 = ~n1299 & n1301;
  assign n1303 = n1285 & ~n1302_1;
  assign n1304 = n1190 & n1201;
  assign n1305 = n1197_1 & n1304;
  assign n1306 = ~n1281 & n1305;
  assign n1307_1 = REG3_REG_0_ & n1292_1;
  assign n1308 = REG2_REG_0_ & n1298;
  assign n1309 = REG1_REG_0_ & n1296;
  assign n1310 = REG0_REG_0_ & n1294;
  assign n1311 = ~n1307_1 & ~n1308;
  assign n1312_1 = ~n1309 & n1311;
  assign n1313 = ~n1310 & n1312_1;
  assign n1314 = ~n1281 & n1313;
  assign n1315 = n1281 & ~n1313;
  assign n1316 = ~n1314 & ~n1315;
  assign n1317_1 = ~n1193 & n1201;
  assign n1318 = n1190 & n1317_1;
  assign n1319 = ~n1316 & n1318;
  assign n1320 = ~n1306 & ~n1319;
  assign n1321 = ~n1283 & ~n1303;
  assign n1322_1 = n1320 & n1321;
  assign n1323 = n1190 & ~n1201;
  assign n1324 = n1193 & n1323;
  assign n1325 = n1197_1 & n1324;
  assign n1326 = ~n1316 & n1325;
  assign n1327_1 = ~n1190 & ~n1197_1;
  assign n1328 = n1193 & n1327_1;
  assign n1329 = ~n1316 & n1328;
  assign n1330 = n1194 & ~n1197_1;
  assign n1331 = n1201 & n1330;
  assign n1332_1 = ~n1316 & n1331;
  assign n1333 = ~n1193 & n1327_1;
  assign n1334 = ~n1316 & n1333;
  assign n1335 = n1193 & ~n1201;
  assign n1336 = ~n1190 & n1335;
  assign n1337_1 = ~n1316 & n1336;
  assign n1338 = ~n1334 & ~n1337_1;
  assign n1339 = ~n1193 & ~n1201;
  assign n1340 = ~n1190 & n1339;
  assign n1341_1 = ~n1316 & n1340;
  assign n1342 = ~n1193 & n1323;
  assign n1343 = ~n1316 & n1342;
  assign n1344 = ~n1341_1 & ~n1343;
  assign n1345 = ~n1326 & ~n1329;
  assign n1346 = ~n1332_1 & n1345;
  assign n1347 = n1338 & n1346;
  assign n1348 = n1344 & n1347;
  assign n1349 = n1322_1 & n1348;
  assign n1350 = n1268 & ~n1349;
  assign n1351 = REG0_REG_0_ & ~n1268;
  assign n494 = n1350 | n1351;
  assign n1353 = REG3_REG_2_ & n1292_1;
  assign n1354 = REG0_REG_2_ & n1294;
  assign n1355 = REG1_REG_2_ & n1296;
  assign n1356 = REG2_REG_2_ & n1298;
  assign n1357 = ~n1353 & ~n1354;
  assign n1358 = ~n1355 & n1357;
  assign n1359 = ~n1356 & n1358;
  assign n1360 = n1285 & ~n1359;
  assign n1361 = IR_REG_31_ & ~n834_1;
  assign n1362 = IR_REG_1_ & ~IR_REG_31_;
  assign n1363 = ~n1361 & ~n1362;
  assign n1364 = n1275 & ~n1363;
  assign n1365 = DATAI_1_ & ~n1275;
  assign n1366 = ~n1364 & ~n1365;
  assign n1367 = ~n1281 & n1366;
  assign n1368 = n1281 & ~n1366;
  assign n1369 = ~n1367 & ~n1368;
  assign n1370 = n1305 & ~n1369;
  assign n1371 = n1282_1 & ~n1366;
  assign n1372 = ~n1302_1 & ~n1366;
  assign n1373 = n1302_1 & n1366;
  assign n1374 = ~n1372 & ~n1373;
  assign n1375 = ~n1281 & ~n1313;
  assign n1376 = n1374 & ~n1375;
  assign n1377 = ~n1374 & n1375;
  assign n1378 = ~n1376 & ~n1377;
  assign n1379 = n1318 & ~n1378;
  assign n1380 = ~n1360 & ~n1370;
  assign n1381 = ~n1371 & n1380;
  assign n1382 = ~n1379 & n1381;
  assign n1383 = ~n1302_1 & n1366;
  assign n1384 = n1302_1 & ~n1366;
  assign n1385 = ~n1383 & ~n1384;
  assign n1386 = ~n1314 & ~n1385;
  assign n1387 = n1314 & n1385;
  assign n1388 = ~n1386 & ~n1387;
  assign n1389 = n1342 & ~n1388;
  assign n1390 = ~n1274 & n1284;
  assign n1391 = ~n1313 & n1390;
  assign n1392 = n1336 & ~n1378;
  assign n1393 = n1340 & ~n1388;
  assign n1394 = ~n1392 & ~n1393;
  assign n1395 = n1331 & ~n1378;
  assign n1396 = n1325 & ~n1378;
  assign n1397 = n1328 & ~n1388;
  assign n1398 = n1333 & ~n1388;
  assign n1399 = ~n1397 & ~n1398;
  assign n1400 = ~n1395 & ~n1396;
  assign n1401 = n1399 & n1400;
  assign n1402 = ~n1389 & ~n1391;
  assign n1403 = n1394 & n1402;
  assign n1404 = n1401 & n1403;
  assign n1405 = n1382 & n1404;
  assign n1406 = n1268 & ~n1405;
  assign n1407 = REG0_REG_1_ & ~n1268;
  assign n499 = n1406 | n1407;
  assign n1409 = ~REG3_REG_3_ & n1292_1;
  assign n1410 = REG0_REG_3_ & n1294;
  assign n1411 = REG1_REG_3_ & n1296;
  assign n1412 = REG2_REG_3_ & n1298;
  assign n1413 = ~n1409 & ~n1410;
  assign n1414 = ~n1411 & n1413;
  assign n1415 = ~n1412 & n1414;
  assign n1416 = n1285 & ~n1415;
  assign n1417 = IR_REG_31_ & n843;
  assign n1418 = IR_REG_2_ & ~IR_REG_31_;
  assign n1419 = ~n1417 & ~n1418;
  assign n1420 = n1275 & ~n1419;
  assign n1421 = DATAI_2_ & ~n1275;
  assign n1422 = ~n1420 & ~n1421;
  assign n1423 = n1281 & n1366;
  assign n1424 = ~n1422 & ~n1423;
  assign n1425 = n1422 & n1423;
  assign n1426 = ~n1424 & ~n1425;
  assign n1427 = n1305 & n1426;
  assign n1428 = n1282_1 & ~n1422;
  assign n1429 = ~n1359 & ~n1422;
  assign n1430 = n1359 & n1422;
  assign n1431 = ~n1429 & ~n1430;
  assign n1432 = ~n1373 & n1375;
  assign n1433 = ~n1372 & ~n1432;
  assign n1434 = n1431 & ~n1433;
  assign n1435 = n1359 & ~n1422;
  assign n1436 = ~n1359 & n1422;
  assign n1437 = ~n1435 & ~n1436;
  assign n1438 = ~n1372 & n1437;
  assign n1439 = ~n1432 & n1438;
  assign n1440 = ~n1434 & ~n1439;
  assign n1441 = n1318 & n1440;
  assign n1442 = ~n1416 & ~n1427;
  assign n1443 = ~n1428 & n1442;
  assign n1444 = ~n1441 & n1443;
  assign n1445 = ~n1302_1 & ~n1314;
  assign n1446 = ~n1314 & n1366;
  assign n1447 = ~n1445 & ~n1446;
  assign n1448 = ~n1383 & n1447;
  assign n1449 = n1437 & n1448;
  assign n1450 = ~n1437 & ~n1448;
  assign n1451 = ~n1449 & ~n1450;
  assign n1452 = n1342 & ~n1451;
  assign n1453 = ~n1302_1 & n1390;
  assign n1454 = n1336 & n1440;
  assign n1455 = n1340 & ~n1451;
  assign n1456 = ~n1454 & ~n1455;
  assign n1457 = n1331 & n1440;
  assign n1458 = n1325 & n1440;
  assign n1459 = n1328 & ~n1451;
  assign n1460 = n1333 & ~n1451;
  assign n1461 = ~n1459 & ~n1460;
  assign n1462 = ~n1457 & ~n1458;
  assign n1463 = n1461 & n1462;
  assign n1464 = ~n1452 & ~n1453;
  assign n1465 = n1456 & n1464;
  assign n1466 = n1463 & n1465;
  assign n1467 = n1444 & n1466;
  assign n1468 = n1268 & ~n1467;
  assign n1469 = REG0_REG_2_ & ~n1268;
  assign n504 = n1468 | n1469;
  assign n1471 = ~REG3_REG_4_ & REG3_REG_3_;
  assign n1472 = REG3_REG_4_ & ~REG3_REG_3_;
  assign n1473 = ~n1471 & ~n1472;
  assign n1474 = n1292_1 & ~n1473;
  assign n1475 = REG0_REG_4_ & n1294;
  assign n1476 = REG1_REG_4_ & n1296;
  assign n1477 = REG2_REG_4_ & n1298;
  assign n1478 = ~n1474 & ~n1475;
  assign n1479 = ~n1476 & n1478;
  assign n1480 = ~n1477 & n1479;
  assign n1481 = n1285 & ~n1480;
  assign n1482 = IR_REG_31_ & n851;
  assign n1483 = IR_REG_3_ & ~IR_REG_31_;
  assign n1484 = ~n1482 & ~n1483;
  assign n1485 = n1275 & ~n1484;
  assign n1486 = DATAI_3_ & ~n1275;
  assign n1487 = ~n1485 & ~n1486;
  assign n1488 = ~n1425 & ~n1487;
  assign n1489 = n1425 & n1487;
  assign n1490 = ~n1488 & ~n1489;
  assign n1491 = n1305 & n1490;
  assign n1492 = n1282_1 & ~n1487;
  assign n1493 = n1372 & ~n1430;
  assign n1494 = ~n1429 & ~n1493;
  assign n1495 = ~n1430 & n1432;
  assign n1496 = n1494 & ~n1495;
  assign n1497 = n1415 & ~n1487;
  assign n1498 = ~n1415 & n1487;
  assign n1499 = ~n1497 & ~n1498;
  assign n1500 = n1496 & ~n1499;
  assign n1501 = ~n1415 & ~n1487;
  assign n1502 = n1415 & n1487;
  assign n1503 = ~n1501 & ~n1502;
  assign n1504 = ~n1496 & ~n1503;
  assign n1505 = ~n1500 & ~n1504;
  assign n1506 = n1318 & ~n1505;
  assign n1507 = ~n1481 & ~n1491;
  assign n1508 = ~n1492 & n1507;
  assign n1509 = ~n1506 & n1508;
  assign n1510 = ~n1435 & ~n1499;
  assign n1511 = ~n1436 & n1448;
  assign n1512 = n1510 & ~n1511;
  assign n1513 = ~n1436 & n1499;
  assign n1514 = ~n1435 & ~n1448;
  assign n1515 = n1513 & ~n1514;
  assign n1516 = ~n1512 & ~n1515;
  assign n1517 = n1342 & ~n1516;
  assign n1518 = ~n1359 & n1390;
  assign n1519 = n1336 & ~n1505;
  assign n1520 = n1340 & ~n1516;
  assign n1521 = ~n1519 & ~n1520;
  assign n1522 = n1331 & ~n1505;
  assign n1523 = n1325 & ~n1505;
  assign n1524 = n1328 & ~n1516;
  assign n1525 = n1333 & ~n1516;
  assign n1526 = ~n1524 & ~n1525;
  assign n1527 = ~n1522 & ~n1523;
  assign n1528 = n1526 & n1527;
  assign n1529 = ~n1517 & ~n1518;
  assign n1530 = n1521 & n1529;
  assign n1531 = n1528 & n1530;
  assign n1532 = n1509 & n1531;
  assign n1533 = n1268 & ~n1532;
  assign n1534 = REG0_REG_3_ & ~n1268;
  assign n509 = n1533 | n1534;
  assign n1536 = REG3_REG_4_ & REG3_REG_3_;
  assign n1537 = ~REG3_REG_5_ & n1536;
  assign n1538 = REG3_REG_5_ & ~n1536;
  assign n1539 = ~n1537 & ~n1538;
  assign n1540 = n1292_1 & ~n1539;
  assign n1541 = REG0_REG_5_ & n1294;
  assign n1542 = REG1_REG_5_ & n1296;
  assign n1543 = REG2_REG_5_ & n1298;
  assign n1544 = ~n1540 & ~n1541;
  assign n1545 = ~n1542 & n1544;
  assign n1546 = ~n1543 & n1545;
  assign n1547 = n1285 & ~n1546;
  assign n1548 = IR_REG_31_ & n859_1;
  assign n1549 = IR_REG_4_ & ~IR_REG_31_;
  assign n1550 = ~n1548 & ~n1549;
  assign n1551 = n1275 & ~n1550;
  assign n1552 = DATAI_4_ & ~n1275;
  assign n1553 = ~n1551 & ~n1552;
  assign n1554 = ~n1489 & ~n1553;
  assign n1555 = n1487 & n1553;
  assign n1556 = n1425 & n1555;
  assign n1557 = ~n1554 & ~n1556;
  assign n1558 = n1305 & n1557;
  assign n1559 = n1282_1 & ~n1553;
  assign n1560 = n1480 & ~n1553;
  assign n1561 = ~n1480 & n1553;
  assign n1562 = ~n1560 & ~n1561;
  assign n1563 = ~n1430 & ~n1502;
  assign n1564 = n1432 & n1563;
  assign n1565 = ~n1501 & ~n1564;
  assign n1566 = ~n1494 & ~n1502;
  assign n1567 = n1565 & ~n1566;
  assign n1568 = ~n1562 & n1567;
  assign n1569 = n1480 & n1553;
  assign n1570 = ~n1480 & ~n1553;
  assign n1571 = ~n1569 & ~n1570;
  assign n1572 = ~n1567 & ~n1571;
  assign n1573 = ~n1568 & ~n1572;
  assign n1574 = n1318 & ~n1573;
  assign n1575 = ~n1547 & ~n1558;
  assign n1576 = ~n1559 & n1575;
  assign n1577 = ~n1574 & n1576;
  assign n1578 = ~n1415 & n1436;
  assign n1579 = n1415 & ~n1436;
  assign n1580 = n1487 & ~n1579;
  assign n1581 = ~n1578 & ~n1580;
  assign n1582 = ~n1435 & ~n1497;
  assign n1583 = ~n1448 & n1582;
  assign n1584 = n1581 & ~n1583;
  assign n1585 = n1562 & n1584;
  assign n1586 = ~n1562 & ~n1584;
  assign n1587 = ~n1585 & ~n1586;
  assign n1588 = n1342 & ~n1587;
  assign n1589 = n1390 & ~n1415;
  assign n1590 = n1336 & ~n1573;
  assign n1591 = n1340 & ~n1587;
  assign n1592 = ~n1590 & ~n1591;
  assign n1593 = n1331 & ~n1573;
  assign n1594 = n1325 & ~n1573;
  assign n1595 = n1328 & ~n1587;
  assign n1596 = n1333 & ~n1587;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = ~n1593 & ~n1594;
  assign n1599 = n1597 & n1598;
  assign n1600 = ~n1588 & ~n1589;
  assign n1601 = n1592 & n1600;
  assign n1602 = n1599 & n1601;
  assign n1603 = n1577 & n1602;
  assign n1604 = n1268 & ~n1603;
  assign n1605 = REG0_REG_4_ & ~n1268;
  assign n514 = n1604 | n1605;
  assign n1607 = REG3_REG_5_ & REG3_REG_3_;
  assign n1608 = REG3_REG_4_ & n1607;
  assign n1609 = ~REG3_REG_6_ & n1608;
  assign n1610 = REG3_REG_6_ & ~n1608;
  assign n1611 = ~n1609 & ~n1610;
  assign n1612 = n1292_1 & ~n1611;
  assign n1613 = REG0_REG_6_ & n1294;
  assign n1614 = REG1_REG_6_ & n1296;
  assign n1615 = REG2_REG_6_ & n1298;
  assign n1616 = ~n1612 & ~n1613;
  assign n1617 = ~n1614 & n1616;
  assign n1618 = ~n1615 & n1617;
  assign n1619 = n1285 & ~n1618;
  assign n1620 = IR_REG_31_ & n871;
  assign n1621 = IR_REG_5_ & ~IR_REG_31_;
  assign n1622 = ~n1620 & ~n1621;
  assign n1623 = n1275 & ~n1622;
  assign n1624 = DATAI_5_ & ~n1275;
  assign n1625 = ~n1623 & ~n1624;
  assign n1626 = ~n1556 & ~n1625;
  assign n1627 = n1556 & n1625;
  assign n1628 = ~n1626 & ~n1627;
  assign n1629 = n1305 & n1628;
  assign n1630 = n1282_1 & ~n1625;
  assign n1631 = ~n1546 & ~n1625;
  assign n1632 = n1546 & n1625;
  assign n1633 = ~n1569 & ~n1632;
  assign n1634 = ~n1631 & n1633;
  assign n1635 = n1567 & ~n1570;
  assign n1636 = n1634 & ~n1635;
  assign n1637 = n1546 & ~n1625;
  assign n1638 = ~n1546 & n1625;
  assign n1639 = ~n1637 & ~n1638;
  assign n1640 = ~n1570 & n1639;
  assign n1641 = ~n1567 & ~n1569;
  assign n1642 = n1640 & ~n1641;
  assign n1643 = ~n1636 & ~n1642;
  assign n1644 = n1318 & n1643;
  assign n1645 = ~n1619 & ~n1629;
  assign n1646 = ~n1630 & n1645;
  assign n1647 = ~n1644 & n1646;
  assign n1648 = ~n1560 & ~n1584;
  assign n1649 = ~n1561 & ~n1648;
  assign n1650 = n1639 & n1649;
  assign n1651 = ~n1639 & ~n1649;
  assign n1652 = ~n1650 & ~n1651;
  assign n1653 = n1342 & ~n1652;
  assign n1654 = n1390 & ~n1480;
  assign n1655 = n1336 & n1643;
  assign n1656 = n1340 & ~n1652;
  assign n1657 = ~n1655 & ~n1656;
  assign n1658 = n1331 & n1643;
  assign n1659 = n1325 & n1643;
  assign n1660 = n1328 & ~n1652;
  assign n1661 = n1333 & ~n1652;
  assign n1662 = ~n1660 & ~n1661;
  assign n1663 = ~n1658 & ~n1659;
  assign n1664 = n1662 & n1663;
  assign n1665 = ~n1653 & ~n1654;
  assign n1666 = n1657 & n1665;
  assign n1667 = n1664 & n1666;
  assign n1668 = n1647 & n1667;
  assign n1669 = n1268 & ~n1668;
  assign n1670 = REG0_REG_5_ & ~n1268;
  assign n519 = n1669 | n1670;
  assign n1672 = REG3_REG_4_ & REG3_REG_5_;
  assign n1673 = REG3_REG_6_ & n1672;
  assign n1674 = REG3_REG_3_ & n1673;
  assign n1675 = ~REG3_REG_7_ & n1674;
  assign n1676 = REG3_REG_7_ & ~n1674;
  assign n1677 = ~n1675 & ~n1676;
  assign n1678 = n1292_1 & ~n1677;
  assign n1679 = REG0_REG_7_ & n1294;
  assign n1680 = REG1_REG_7_ & n1296;
  assign n1681 = REG2_REG_7_ & n1298;
  assign n1682 = ~n1678 & ~n1679;
  assign n1683 = ~n1680 & n1682;
  assign n1684 = ~n1681 & n1683;
  assign n1685 = n1285 & ~n1684;
  assign n1686 = IR_REG_31_ & n879_1;
  assign n1687 = IR_REG_6_ & ~IR_REG_31_;
  assign n1688 = ~n1686 & ~n1687;
  assign n1689 = n1275 & ~n1688;
  assign n1690 = DATAI_6_ & ~n1275;
  assign n1691 = ~n1689 & ~n1690;
  assign n1692 = ~n1627 & ~n1691;
  assign n1693 = n1625 & n1691;
  assign n1694 = n1556 & n1693;
  assign n1695 = ~n1692 & ~n1694;
  assign n1696 = n1305 & n1695;
  assign n1697 = n1282_1 & ~n1691;
  assign n1698 = n1618 & ~n1691;
  assign n1699 = ~n1618 & n1691;
  assign n1700 = ~n1698 & ~n1699;
  assign n1701 = n1372 & n1633;
  assign n1702 = n1563 & n1701;
  assign n1703 = n1570 & ~n1625;
  assign n1704 = n1563 & n1633;
  assign n1705 = n1432 & n1704;
  assign n1706 = ~n1702 & ~n1703;
  assign n1707 = ~n1705 & n1706;
  assign n1708 = n1501 & n1633;
  assign n1709 = ~n1570 & n1625;
  assign n1710 = ~n1546 & ~n1709;
  assign n1711 = n1429 & ~n1502;
  assign n1712 = n1633 & n1711;
  assign n1713 = ~n1708 & ~n1710;
  assign n1714 = ~n1712 & n1713;
  assign n1715 = n1707 & n1714;
  assign n1716 = ~n1700 & n1715;
  assign n1717 = n1618 & n1691;
  assign n1718 = ~n1618 & ~n1691;
  assign n1719 = ~n1717 & ~n1718;
  assign n1720 = ~n1715 & ~n1719;
  assign n1721 = ~n1716 & ~n1720;
  assign n1722 = n1318 & ~n1721;
  assign n1723 = ~n1685 & ~n1696;
  assign n1724 = ~n1697 & n1723;
  assign n1725 = ~n1722 & n1724;
  assign n1726 = ~n1637 & ~n1700;
  assign n1727 = ~n1638 & n1649;
  assign n1728 = n1726 & ~n1727;
  assign n1729 = ~n1638 & ~n1699;
  assign n1730 = ~n1698 & n1729;
  assign n1731 = ~n1637 & ~n1649;
  assign n1732 = n1730 & ~n1731;
  assign n1733 = ~n1728 & ~n1732;
  assign n1734 = n1342 & ~n1733;
  assign n1735 = n1390 & ~n1546;
  assign n1736 = n1336 & ~n1721;
  assign n1737 = n1340 & ~n1733;
  assign n1738 = ~n1736 & ~n1737;
  assign n1739 = n1331 & ~n1721;
  assign n1740 = n1325 & ~n1721;
  assign n1741 = n1328 & ~n1733;
  assign n1742 = n1333 & ~n1733;
  assign n1743 = ~n1741 & ~n1742;
  assign n1744 = ~n1739 & ~n1740;
  assign n1745 = n1743 & n1744;
  assign n1746 = ~n1734 & ~n1735;
  assign n1747 = n1738 & n1746;
  assign n1748 = n1745 & n1747;
  assign n1749 = n1725 & n1748;
  assign n1750 = n1268 & ~n1749;
  assign n1751 = REG0_REG_6_ & ~n1268;
  assign n524 = n1750 | n1751;
  assign n1753 = REG3_REG_3_ & REG3_REG_7_;
  assign n1754 = REG3_REG_6_ & n1753;
  assign n1755 = REG3_REG_4_ & n1754;
  assign n1756 = REG3_REG_5_ & n1755;
  assign n1757 = ~REG3_REG_8_ & n1756;
  assign n1758 = REG3_REG_8_ & ~n1756;
  assign n1759 = ~n1757 & ~n1758;
  assign n1760 = n1292_1 & ~n1759;
  assign n1761 = REG0_REG_8_ & n1294;
  assign n1762 = REG1_REG_8_ & n1296;
  assign n1763 = REG2_REG_8_ & n1298;
  assign n1764 = ~n1760 & ~n1761;
  assign n1765 = ~n1762 & n1764;
  assign n1766 = ~n1763 & n1765;
  assign n1767 = n1285 & ~n1766;
  assign n1768 = IR_REG_31_ & n888;
  assign n1769 = IR_REG_7_ & ~IR_REG_31_;
  assign n1770 = ~n1768 & ~n1769;
  assign n1771 = n1275 & ~n1770;
  assign n1772 = DATAI_7_ & ~n1275;
  assign n1773 = ~n1771 & ~n1772;
  assign n1774 = ~n1694 & ~n1773;
  assign n1775 = n1694 & n1773;
  assign n1776 = ~n1774 & ~n1775;
  assign n1777 = n1305 & n1776;
  assign n1778 = n1282_1 & ~n1773;
  assign n1779 = n1684 & n1773;
  assign n1780 = ~n1717 & ~n1779;
  assign n1781 = ~n1684 & ~n1773;
  assign n1782 = n1780 & ~n1781;
  assign n1783 = n1715 & ~n1718;
  assign n1784 = n1782 & ~n1783;
  assign n1785 = n1684 & ~n1773;
  assign n1786 = ~n1684 & n1773;
  assign n1787 = ~n1785 & ~n1786;
  assign n1788 = ~n1718 & n1787;
  assign n1789 = ~n1715 & ~n1717;
  assign n1790 = n1788 & ~n1789;
  assign n1791 = ~n1784 & ~n1790;
  assign n1792 = n1318 & n1791;
  assign n1793 = ~n1767 & ~n1777;
  assign n1794 = ~n1778 & n1793;
  assign n1795 = ~n1792 & n1794;
  assign n1796 = n1561 & ~n1637;
  assign n1797 = n1729 & ~n1796;
  assign n1798 = ~n1698 & ~n1797;
  assign n1799 = ~n1637 & ~n1698;
  assign n1800 = ~n1560 & n1799;
  assign n1801 = ~n1584 & n1800;
  assign n1802 = ~n1798 & ~n1801;
  assign n1803 = n1787 & n1802;
  assign n1804 = ~n1787 & ~n1802;
  assign n1805 = ~n1803 & ~n1804;
  assign n1806 = n1342 & ~n1805;
  assign n1807 = n1390 & ~n1618;
  assign n1808 = n1336 & n1791;
  assign n1809 = n1340 & ~n1805;
  assign n1810 = ~n1808 & ~n1809;
  assign n1811 = n1331 & n1791;
  assign n1812 = n1325 & n1791;
  assign n1813 = n1328 & ~n1805;
  assign n1814 = n1333 & ~n1805;
  assign n1815 = ~n1813 & ~n1814;
  assign n1816 = ~n1811 & ~n1812;
  assign n1817 = n1815 & n1816;
  assign n1818 = ~n1806 & ~n1807;
  assign n1819 = n1810 & n1818;
  assign n1820 = n1817 & n1819;
  assign n1821 = n1795 & n1820;
  assign n1822 = n1268 & ~n1821;
  assign n1823 = REG0_REG_7_ & ~n1268;
  assign n529 = n1822 | n1823;
  assign n1825 = REG3_REG_8_ & n1756;
  assign n1826 = ~REG3_REG_9_ & n1825;
  assign n1827 = REG3_REG_9_ & ~n1825;
  assign n1828 = ~n1826 & ~n1827;
  assign n1829 = n1292_1 & ~n1828;
  assign n1830 = REG0_REG_9_ & n1294;
  assign n1831 = REG1_REG_9_ & n1296;
  assign n1832 = REG2_REG_9_ & n1298;
  assign n1833 = ~n1829 & ~n1830;
  assign n1834 = ~n1831 & n1833;
  assign n1835 = ~n1832 & n1834;
  assign n1836 = n1285 & ~n1835;
  assign n1837 = IR_REG_31_ & n896;
  assign n1838 = IR_REG_8_ & ~IR_REG_31_;
  assign n1839 = ~n1837 & ~n1838;
  assign n1840 = n1275 & ~n1839;
  assign n1841 = DATAI_8_ & ~n1275;
  assign n1842 = ~n1840 & ~n1841;
  assign n1843 = n1775 & n1842;
  assign n1844 = ~n1775 & ~n1842;
  assign n1845 = ~n1843 & ~n1844;
  assign n1846 = n1305 & n1845;
  assign n1847 = n1282_1 & ~n1842;
  assign n1848 = n1718 & ~n1773;
  assign n1849 = ~n1718 & n1773;
  assign n1850 = ~n1684 & ~n1849;
  assign n1851 = ~n1848 & ~n1850;
  assign n1852 = ~n1715 & n1780;
  assign n1853 = n1851 & ~n1852;
  assign n1854 = n1766 & ~n1842;
  assign n1855 = ~n1766 & n1842;
  assign n1856 = ~n1854 & ~n1855;
  assign n1857 = n1853 & ~n1856;
  assign n1858 = n1766 & n1842;
  assign n1859 = ~n1766 & ~n1842;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = ~n1853 & ~n1860;
  assign n1862 = ~n1857 & ~n1861;
  assign n1863 = n1318 & ~n1862;
  assign n1864 = ~n1836 & ~n1846;
  assign n1865 = ~n1847 & n1864;
  assign n1866 = ~n1863 & n1865;
  assign n1867 = ~n1785 & ~n1856;
  assign n1868 = ~n1786 & n1802;
  assign n1869 = n1867 & ~n1868;
  assign n1870 = ~n1786 & n1856;
  assign n1871 = ~n1785 & ~n1802;
  assign n1872 = n1870 & ~n1871;
  assign n1873 = ~n1869 & ~n1872;
  assign n1874 = n1342 & ~n1873;
  assign n1875 = n1390 & ~n1684;
  assign n1876 = n1336 & ~n1862;
  assign n1877 = n1340 & ~n1873;
  assign n1878 = ~n1876 & ~n1877;
  assign n1879 = n1331 & ~n1862;
  assign n1880 = n1325 & ~n1862;
  assign n1881 = n1328 & ~n1873;
  assign n1882 = n1333 & ~n1873;
  assign n1883 = ~n1881 & ~n1882;
  assign n1884 = ~n1879 & ~n1880;
  assign n1885 = n1883 & n1884;
  assign n1886 = ~n1874 & ~n1875;
  assign n1887 = n1878 & n1886;
  assign n1888 = n1885 & n1887;
  assign n1889 = n1866 & n1888;
  assign n1890 = n1268 & ~n1889;
  assign n1891 = REG0_REG_8_ & ~n1268;
  assign n534 = n1890 | n1891;
  assign n1893 = REG3_REG_9_ & REG3_REG_8_;
  assign n1894 = n1756 & n1893;
  assign n1895 = ~REG3_REG_10_ & n1894;
  assign n1896 = REG3_REG_10_ & ~n1894;
  assign n1897 = ~n1895 & ~n1896;
  assign n1898 = n1292_1 & ~n1897;
  assign n1899 = REG0_REG_10_ & n1294;
  assign n1900 = REG1_REG_10_ & n1296;
  assign n1901 = REG2_REG_10_ & n1298;
  assign n1902 = ~n1898 & ~n1899;
  assign n1903 = ~n1900 & n1902;
  assign n1904 = ~n1901 & n1903;
  assign n1905 = n1285 & ~n1904;
  assign n1906 = n1773 & n1842;
  assign n1907 = n1694 & n1906;
  assign n1908 = IR_REG_31_ & n906;
  assign n1909 = IR_REG_9_ & ~IR_REG_31_;
  assign n1910 = ~n1908 & ~n1909;
  assign n1911 = n1275 & ~n1910;
  assign n1912 = DATAI_9_ & ~n1275;
  assign n1913 = ~n1911 & ~n1912;
  assign n1914 = n1907 & n1913;
  assign n1915 = ~n1907 & ~n1913;
  assign n1916 = ~n1914 & ~n1915;
  assign n1917 = n1305 & n1916;
  assign n1918 = n1282_1 & ~n1913;
  assign n1919 = n1835 & ~n1913;
  assign n1920 = ~n1835 & n1913;
  assign n1921 = ~n1919 & ~n1920;
  assign n1922 = ~n1853 & ~n1858;
  assign n1923 = ~n1859 & ~n1922;
  assign n1924 = ~n1921 & n1923;
  assign n1925 = n1835 & n1913;
  assign n1926 = ~n1835 & ~n1913;
  assign n1927 = ~n1925 & ~n1926;
  assign n1928 = ~n1923 & ~n1927;
  assign n1929 = ~n1924 & ~n1928;
  assign n1930 = n1318 & ~n1929;
  assign n1931 = ~n1905 & ~n1917;
  assign n1932 = ~n1918 & n1931;
  assign n1933 = ~n1930 & n1932;
  assign n1934 = ~n1785 & ~n1854;
  assign n1935 = n1798 & n1934;
  assign n1936 = ~n1766 & n1786;
  assign n1937 = n1766 & ~n1786;
  assign n1938 = n1842 & ~n1937;
  assign n1939 = ~n1936 & ~n1938;
  assign n1940 = ~n1935 & n1939;
  assign n1941 = n1800 & n1934;
  assign n1942 = ~n1584 & n1941;
  assign n1943 = n1940 & ~n1942;
  assign n1944 = n1921 & n1943;
  assign n1945 = ~n1921 & ~n1943;
  assign n1946 = ~n1944 & ~n1945;
  assign n1947 = n1342 & ~n1946;
  assign n1948 = n1390 & ~n1766;
  assign n1949 = n1336 & ~n1929;
  assign n1950 = n1340 & ~n1946;
  assign n1951 = ~n1949 & ~n1950;
  assign n1952 = n1331 & ~n1929;
  assign n1953 = n1325 & ~n1929;
  assign n1954 = n1328 & ~n1946;
  assign n1955 = n1333 & ~n1946;
  assign n1956 = ~n1954 & ~n1955;
  assign n1957 = ~n1952 & ~n1953;
  assign n1958 = n1956 & n1957;
  assign n1959 = ~n1947 & ~n1948;
  assign n1960 = n1951 & n1959;
  assign n1961 = n1958 & n1960;
  assign n1962 = n1933 & n1961;
  assign n1963 = n1268 & ~n1962;
  assign n1964 = REG0_REG_9_ & ~n1268;
  assign n539 = n1963 | n1964;
  assign n1966 = REG3_REG_10_ & n1894;
  assign n1967 = ~REG3_REG_11_ & n1966;
  assign n1968 = REG3_REG_11_ & ~n1966;
  assign n1969 = ~n1967 & ~n1968;
  assign n1970 = n1292_1 & ~n1969;
  assign n1971 = REG0_REG_11_ & n1294;
  assign n1972 = REG1_REG_11_ & n1296;
  assign n1973 = REG2_REG_11_ & n1298;
  assign n1974 = ~n1970 & ~n1971;
  assign n1975 = ~n1972 & n1974;
  assign n1976 = ~n1973 & n1975;
  assign n1977 = n1285 & ~n1976;
  assign n1978 = IR_REG_31_ & n914_1;
  assign n1979 = IR_REG_10_ & ~IR_REG_31_;
  assign n1980 = ~n1978 & ~n1979;
  assign n1981 = n1275 & ~n1980;
  assign n1982 = DATAI_10_ & ~n1275;
  assign n1983 = ~n1981 & ~n1982;
  assign n1984 = n1914 & n1983;
  assign n1985 = ~n1914 & ~n1983;
  assign n1986 = ~n1984 & ~n1985;
  assign n1987 = n1305 & n1986;
  assign n1988 = n1282_1 & ~n1983;
  assign n1989 = ~n1904 & ~n1983;
  assign n1990 = n1904 & n1983;
  assign n1991 = ~n1925 & ~n1990;
  assign n1992 = ~n1989 & n1991;
  assign n1993 = n1923 & ~n1926;
  assign n1994 = n1992 & ~n1993;
  assign n1995 = n1904 & ~n1983;
  assign n1996 = ~n1904 & n1983;
  assign n1997 = ~n1995 & ~n1996;
  assign n1998 = ~n1926 & n1997;
  assign n1999 = ~n1923 & ~n1925;
  assign n2000 = n1998 & ~n1999;
  assign n2001 = ~n1994 & ~n2000;
  assign n2002 = n1318 & n2001;
  assign n2003 = ~n1977 & ~n1987;
  assign n2004 = ~n1988 & n2003;
  assign n2005 = ~n2002 & n2004;
  assign n2006 = ~n1919 & ~n1943;
  assign n2007 = ~n1920 & ~n2006;
  assign n2008 = n1997 & n2007;
  assign n2009 = ~n1997 & ~n2007;
  assign n2010 = ~n2008 & ~n2009;
  assign n2011 = n1342 & ~n2010;
  assign n2012 = n1390 & ~n1835;
  assign n2013 = n1336 & n2001;
  assign n2014 = n1340 & ~n2010;
  assign n2015 = ~n2013 & ~n2014;
  assign n2016 = n1331 & n2001;
  assign n2017 = n1325 & n2001;
  assign n2018 = n1328 & ~n2010;
  assign n2019 = n1333 & ~n2010;
  assign n2020 = ~n2018 & ~n2019;
  assign n2021 = ~n2016 & ~n2017;
  assign n2022 = n2020 & n2021;
  assign n2023 = ~n2011 & ~n2012;
  assign n2024 = n2015 & n2023;
  assign n2025 = n2022 & n2024;
  assign n2026 = n2005 & n2025;
  assign n2027 = n1268 & ~n2026;
  assign n2028 = REG0_REG_10_ & ~n1268;
  assign n544 = n2027 | n2028;
  assign n2030 = REG3_REG_11_ & REG3_REG_10_;
  assign n2031 = n1894 & n2030;
  assign n2032 = ~REG3_REG_12_ & n2031;
  assign n2033 = REG3_REG_12_ & ~n2031;
  assign n2034 = ~n2032 & ~n2033;
  assign n2035 = n1292_1 & ~n2034;
  assign n2036 = REG0_REG_12_ & n1294;
  assign n2037 = REG1_REG_12_ & n1296;
  assign n2038 = REG2_REG_12_ & n1298;
  assign n2039 = ~n2035 & ~n2036;
  assign n2040 = ~n2037 & n2039;
  assign n2041 = ~n2038 & n2040;
  assign n2042 = n1285 & ~n2041;
  assign n2043 = n1913 & n1983;
  assign n2044 = n1907 & n2043;
  assign n2045 = IR_REG_31_ & n923;
  assign n2046 = IR_REG_11_ & ~IR_REG_31_;
  assign n2047 = ~n2045 & ~n2046;
  assign n2048 = n1275 & ~n2047;
  assign n2049 = DATAI_11_ & ~n1275;
  assign n2050 = ~n2048 & ~n2049;
  assign n2051 = n2044 & n2050;
  assign n2052 = ~n2044 & ~n2050;
  assign n2053 = ~n2051 & ~n2052;
  assign n2054 = n1305 & n2053;
  assign n2055 = n1282_1 & ~n2050;
  assign n2056 = ~n1858 & n1991;
  assign n2057 = ~n1851 & n2056;
  assign n2058 = ~n1926 & ~n1989;
  assign n2059 = n1859 & n1991;
  assign n2060 = n2058 & ~n2059;
  assign n2061 = ~n1990 & ~n2060;
  assign n2062 = ~n2057 & ~n2061;
  assign n2063 = n1780 & n2056;
  assign n2064 = ~n1715 & n2063;
  assign n2065 = n2062 & ~n2064;
  assign n2066 = n1976 & ~n2050;
  assign n2067 = ~n1976 & n2050;
  assign n2068 = ~n2066 & ~n2067;
  assign n2069 = n2065 & ~n2068;
  assign n2070 = n1976 & n2050;
  assign n2071 = ~n1976 & ~n2050;
  assign n2072 = ~n2070 & ~n2071;
  assign n2073 = ~n2065 & ~n2072;
  assign n2074 = ~n2069 & ~n2073;
  assign n2075 = n1318 & ~n2074;
  assign n2076 = ~n2042 & ~n2054;
  assign n2077 = ~n2055 & n2076;
  assign n2078 = ~n2075 & n2077;
  assign n2079 = ~n1995 & ~n2068;
  assign n2080 = ~n1996 & n2007;
  assign n2081 = n2079 & ~n2080;
  assign n2082 = ~n1996 & ~n2067;
  assign n2083 = ~n2066 & n2082;
  assign n2084 = ~n1995 & ~n2007;
  assign n2085 = n2083 & ~n2084;
  assign n2086 = ~n2081 & ~n2085;
  assign n2087 = n1342 & ~n2086;
  assign n2088 = n1390 & ~n1904;
  assign n2089 = n1336 & ~n2074;
  assign n2090 = n1340 & ~n2086;
  assign n2091 = ~n2089 & ~n2090;
  assign n2092 = n1331 & ~n2074;
  assign n2093 = n1325 & ~n2074;
  assign n2094 = n1328 & ~n2086;
  assign n2095 = n1333 & ~n2086;
  assign n2096 = ~n2094 & ~n2095;
  assign n2097 = ~n2092 & ~n2093;
  assign n2098 = n2096 & n2097;
  assign n2099 = ~n2087 & ~n2088;
  assign n2100 = n2091 & n2099;
  assign n2101 = n2098 & n2100;
  assign n2102 = n2078 & n2101;
  assign n2103 = n1268 & ~n2102;
  assign n2104 = REG0_REG_11_ & ~n1268;
  assign n549 = n2103 | n2104;
  assign n2106 = REG3_REG_12_ & n2031;
  assign n2107 = ~REG3_REG_13_ & n2106;
  assign n2108 = REG3_REG_13_ & ~n2106;
  assign n2109 = ~n2107 & ~n2108;
  assign n2110 = n1292_1 & ~n2109;
  assign n2111 = REG0_REG_13_ & n1294;
  assign n2112 = REG1_REG_13_ & n1296;
  assign n2113 = REG2_REG_13_ & n1298;
  assign n2114 = ~n2110 & ~n2111;
  assign n2115 = ~n2112 & n2114;
  assign n2116 = ~n2113 & n2115;
  assign n2117 = n1285 & ~n2116;
  assign n2118 = IR_REG_31_ & n931;
  assign n2119 = IR_REG_12_ & ~IR_REG_31_;
  assign n2120 = ~n2118 & ~n2119;
  assign n2121 = n1275 & ~n2120;
  assign n2122 = DATAI_12_ & ~n1275;
  assign n2123 = ~n2121 & ~n2122;
  assign n2124 = n2051 & n2123;
  assign n2125 = ~n2051 & ~n2123;
  assign n2126 = ~n2124 & ~n2125;
  assign n2127 = n1305 & n2126;
  assign n2128 = n1282_1 & ~n2123;
  assign n2129 = n2041 & ~n2123;
  assign n2130 = ~n2041 & n2123;
  assign n2131 = ~n2129 & ~n2130;
  assign n2132 = ~n2065 & ~n2070;
  assign n2133 = ~n2071 & ~n2132;
  assign n2134 = ~n2131 & n2133;
  assign n2135 = n2041 & n2123;
  assign n2136 = ~n2041 & ~n2123;
  assign n2137 = ~n2135 & ~n2136;
  assign n2138 = ~n2133 & ~n2137;
  assign n2139 = ~n2134 & ~n2138;
  assign n2140 = n1318 & ~n2139;
  assign n2141 = ~n2117 & ~n2127;
  assign n2142 = ~n2128 & n2141;
  assign n2143 = ~n2140 & n2142;
  assign n2144 = ~n1995 & ~n2066;
  assign n2145 = ~n1919 & n2144;
  assign n2146 = ~n1943 & n2145;
  assign n2147 = n1920 & n2144;
  assign n2148 = n2082 & ~n2147;
  assign n2149 = ~n2066 & ~n2148;
  assign n2150 = ~n2146 & ~n2149;
  assign n2151 = ~n2131 & ~n2150;
  assign n2152 = n2131 & n2150;
  assign n2153 = ~n2151 & ~n2152;
  assign n2154 = n1342 & ~n2153;
  assign n2155 = n1390 & ~n1976;
  assign n2156 = n1336 & ~n2139;
  assign n2157 = n1340 & ~n2153;
  assign n2158 = ~n2156 & ~n2157;
  assign n2159 = n1331 & ~n2139;
  assign n2160 = n1325 & ~n2139;
  assign n2161 = n1328 & ~n2153;
  assign n2162 = n1333 & ~n2153;
  assign n2163 = ~n2161 & ~n2162;
  assign n2164 = ~n2159 & ~n2160;
  assign n2165 = n2163 & n2164;
  assign n2166 = ~n2154 & ~n2155;
  assign n2167 = n2158 & n2166;
  assign n2168 = n2165 & n2167;
  assign n2169 = n2143 & n2168;
  assign n2170 = n1268 & ~n2169;
  assign n2171 = REG0_REG_12_ & ~n1268;
  assign n554 = n2170 | n2171;
  assign n2173 = REG3_REG_13_ & REG3_REG_12_;
  assign n2174 = n2031 & n2173;
  assign n2175 = ~REG3_REG_14_ & n2174;
  assign n2176 = REG3_REG_14_ & ~n2174;
  assign n2177 = ~n2175 & ~n2176;
  assign n2178 = n1292_1 & ~n2177;
  assign n2179 = REG0_REG_14_ & n1294;
  assign n2180 = REG1_REG_14_ & n1296;
  assign n2181 = REG2_REG_14_ & n1298;
  assign n2182 = ~n2178 & ~n2179;
  assign n2183 = ~n2180 & n2182;
  assign n2184 = ~n2181 & n2183;
  assign n2185 = n1285 & ~n2184;
  assign n2186 = n2050 & n2123;
  assign n2187 = n2044 & n2186;
  assign n2188 = IR_REG_31_ & n948;
  assign n2189 = IR_REG_13_ & ~IR_REG_31_;
  assign n2190 = ~n2188 & ~n2189;
  assign n2191 = n1275 & ~n2190;
  assign n2192 = DATAI_13_ & ~n1275;
  assign n2193 = ~n2191 & ~n2192;
  assign n2194 = n2187 & n2193;
  assign n2195 = ~n2187 & ~n2193;
  assign n2196 = ~n2194 & ~n2195;
  assign n2197 = n1305 & n2196;
  assign n2198 = n1282_1 & ~n2193;
  assign n2199 = ~n2116 & ~n2193;
  assign n2200 = n2116 & n2193;
  assign n2201 = ~n2135 & ~n2200;
  assign n2202 = ~n2199 & n2201;
  assign n2203 = n2133 & ~n2136;
  assign n2204 = n2202 & ~n2203;
  assign n2205 = n2116 & ~n2193;
  assign n2206 = ~n2116 & n2193;
  assign n2207 = ~n2205 & ~n2206;
  assign n2208 = ~n2136 & n2207;
  assign n2209 = ~n2133 & ~n2135;
  assign n2210 = n2208 & ~n2209;
  assign n2211 = ~n2204 & ~n2210;
  assign n2212 = n1318 & n2211;
  assign n2213 = ~n2185 & ~n2197;
  assign n2214 = ~n2198 & n2213;
  assign n2215 = ~n2212 & n2214;
  assign n2216 = ~n2129 & n2145;
  assign n2217 = ~n1943 & n2216;
  assign n2218 = ~n2130 & ~n2149;
  assign n2219 = ~n2129 & ~n2218;
  assign n2220 = ~n2217 & ~n2219;
  assign n2221 = ~n2207 & ~n2220;
  assign n2222 = n2207 & n2220;
  assign n2223 = ~n2221 & ~n2222;
  assign n2224 = n1342 & ~n2223;
  assign n2225 = n1390 & ~n2041;
  assign n2226 = n1336 & n2211;
  assign n2227 = n1340 & ~n2223;
  assign n2228 = ~n2226 & ~n2227;
  assign n2229 = n1331 & n2211;
  assign n2230 = n1325 & n2211;
  assign n2231 = n1328 & ~n2223;
  assign n2232 = n1333 & ~n2223;
  assign n2233 = ~n2231 & ~n2232;
  assign n2234 = ~n2229 & ~n2230;
  assign n2235 = n2233 & n2234;
  assign n2236 = ~n2224 & ~n2225;
  assign n2237 = n2228 & n2236;
  assign n2238 = n2235 & n2237;
  assign n2239 = n2215 & n2238;
  assign n2240 = n1268 & ~n2239;
  assign n2241 = REG0_REG_13_ & ~n1268;
  assign n559 = n2240 | n2241;
  assign n2243 = REG3_REG_14_ & n2174;
  assign n2244 = ~REG3_REG_15_ & n2243;
  assign n2245 = REG3_REG_15_ & ~n2243;
  assign n2246 = ~n2244 & ~n2245;
  assign n2247 = n1292_1 & ~n2246;
  assign n2248 = REG0_REG_15_ & n1294;
  assign n2249 = REG1_REG_15_ & n1296;
  assign n2250 = REG2_REG_15_ & n1298;
  assign n2251 = ~n2247 & ~n2248;
  assign n2252 = ~n2249 & n2251;
  assign n2253 = ~n2250 & n2252;
  assign n2254 = n1285 & ~n2253;
  assign n2255 = IR_REG_31_ & n956;
  assign n2256 = IR_REG_14_ & ~IR_REG_31_;
  assign n2257 = ~n2255 & ~n2256;
  assign n2258 = n1275 & ~n2257;
  assign n2259 = DATAI_14_ & ~n1275;
  assign n2260 = ~n2258 & ~n2259;
  assign n2261 = n2194 & n2260;
  assign n2262 = ~n2194 & ~n2260;
  assign n2263 = ~n2261 & ~n2262;
  assign n2264 = n1305 & n2263;
  assign n2265 = n1282_1 & ~n2260;
  assign n2266 = ~n2136 & ~n2199;
  assign n2267 = n2071 & n2201;
  assign n2268 = n2266 & ~n2267;
  assign n2269 = ~n2200 & ~n2268;
  assign n2270 = ~n2070 & n2201;
  assign n2271 = ~n2065 & n2270;
  assign n2272 = ~n2269 & ~n2271;
  assign n2273 = n2184 & ~n2260;
  assign n2274 = ~n2184 & n2260;
  assign n2275 = ~n2273 & ~n2274;
  assign n2276 = n2272 & ~n2275;
  assign n2277 = ~n2272 & n2275;
  assign n2278 = ~n2276 & ~n2277;
  assign n2279 = n1318 & ~n2278;
  assign n2280 = ~n2254 & ~n2264;
  assign n2281 = ~n2265 & n2280;
  assign n2282 = ~n2279 & n2281;
  assign n2283 = ~n2205 & n2219;
  assign n2284 = ~n2205 & n2216;
  assign n2285 = ~n1943 & n2284;
  assign n2286 = ~n2206 & ~n2283;
  assign n2287 = ~n2285 & n2286;
  assign n2288 = n2275 & n2287;
  assign n2289 = ~n2275 & ~n2287;
  assign n2290 = ~n2288 & ~n2289;
  assign n2291 = n1342 & ~n2290;
  assign n2292 = n1390 & ~n2116;
  assign n2293 = n1336 & ~n2278;
  assign n2294 = n1340 & ~n2290;
  assign n2295 = ~n2293 & ~n2294;
  assign n2296 = n1331 & ~n2278;
  assign n2297 = n1325 & ~n2278;
  assign n2298 = n1328 & ~n2290;
  assign n2299 = n1333 & ~n2290;
  assign n2300 = ~n2298 & ~n2299;
  assign n2301 = ~n2296 & ~n2297;
  assign n2302 = n2300 & n2301;
  assign n2303 = ~n2291 & ~n2292;
  assign n2304 = n2295 & n2303;
  assign n2305 = n2302 & n2304;
  assign n2306 = n2282 & n2305;
  assign n2307 = n1268 & ~n2306;
  assign n2308 = REG0_REG_14_ & ~n1268;
  assign n564 = n2307 | n2308;
  assign n2310 = REG3_REG_15_ & REG3_REG_14_;
  assign n2311 = n2174 & n2310;
  assign n2312 = ~REG3_REG_16_ & n2311;
  assign n2313 = REG3_REG_16_ & ~n2311;
  assign n2314 = ~n2312 & ~n2313;
  assign n2315 = n1292_1 & ~n2314;
  assign n2316 = REG0_REG_16_ & n1294;
  assign n2317 = REG1_REG_16_ & n1296;
  assign n2318 = REG2_REG_16_ & n1298;
  assign n2319 = ~n2315 & ~n2316;
  assign n2320 = ~n2317 & n2319;
  assign n2321 = ~n2318 & n2320;
  assign n2322 = n1285 & ~n2321;
  assign n2323 = n2193 & n2260;
  assign n2324 = n2187 & n2323;
  assign n2325 = IR_REG_31_ & n965;
  assign n2326 = IR_REG_15_ & ~IR_REG_31_;
  assign n2327 = ~n2325 & ~n2326;
  assign n2328 = n1275 & ~n2327;
  assign n2329 = DATAI_15_ & ~n1275;
  assign n2330 = ~n2328 & ~n2329;
  assign n2331 = n2324 & n2330;
  assign n2332 = ~n2324 & ~n2330;
  assign n2333 = ~n2331 & ~n2332;
  assign n2334 = n1305 & n2333;
  assign n2335 = n1282_1 & ~n2330;
  assign n2336 = ~n2184 & ~n2260;
  assign n2337 = ~n2269 & ~n2336;
  assign n2338 = n2184 & n2260;
  assign n2339 = ~n2337 & ~n2338;
  assign n2340 = n2270 & ~n2338;
  assign n2341 = ~n2065 & n2340;
  assign n2342 = ~n2339 & ~n2341;
  assign n2343 = n2253 & ~n2330;
  assign n2344 = ~n2253 & n2330;
  assign n2345 = ~n2343 & ~n2344;
  assign n2346 = n2342 & ~n2345;
  assign n2347 = ~n2342 & n2345;
  assign n2348 = ~n2346 & ~n2347;
  assign n2349 = n1318 & ~n2348;
  assign n2350 = ~n2322 & ~n2334;
  assign n2351 = ~n2335 & n2350;
  assign n2352 = ~n2349 & n2351;
  assign n2353 = ~n2273 & ~n2287;
  assign n2354 = ~n2274 & ~n2353;
  assign n2355 = n2345 & n2354;
  assign n2356 = ~n2345 & ~n2354;
  assign n2357 = ~n2355 & ~n2356;
  assign n2358 = n1342 & ~n2357;
  assign n2359 = n1390 & ~n2184;
  assign n2360 = n1336 & ~n2348;
  assign n2361 = n1340 & ~n2357;
  assign n2362 = ~n2360 & ~n2361;
  assign n2363 = n1331 & ~n2348;
  assign n2364 = n1325 & ~n2348;
  assign n2365 = n1328 & ~n2357;
  assign n2366 = n1333 & ~n2357;
  assign n2367 = ~n2365 & ~n2366;
  assign n2368 = ~n2363 & ~n2364;
  assign n2369 = n2367 & n2368;
  assign n2370 = ~n2358 & ~n2359;
  assign n2371 = n2362 & n2370;
  assign n2372 = n2369 & n2371;
  assign n2373 = n2352 & n2372;
  assign n2374 = n1268 & ~n2373;
  assign n2375 = REG0_REG_15_ & ~n1268;
  assign n569 = n2374 | n2375;
  assign n2377 = REG3_REG_16_ & n2311;
  assign n2378 = ~REG3_REG_17_ & n2377;
  assign n2379 = REG3_REG_17_ & ~n2377;
  assign n2380 = ~n2378 & ~n2379;
  assign n2381 = n1292_1 & ~n2380;
  assign n2382 = REG0_REG_17_ & n1294;
  assign n2383 = REG1_REG_17_ & n1296;
  assign n2384 = REG2_REG_17_ & n1298;
  assign n2385 = ~n2381 & ~n2382;
  assign n2386 = ~n2383 & n2385;
  assign n2387 = ~n2384 & n2386;
  assign n2388 = n1285 & ~n2387;
  assign n2389 = IR_REG_31_ & n973;
  assign n2390 = IR_REG_16_ & ~IR_REG_31_;
  assign n2391 = ~n2389 & ~n2390;
  assign n2392 = n1275 & ~n2391;
  assign n2393 = DATAI_16_ & ~n1275;
  assign n2394 = ~n2392 & ~n2393;
  assign n2395 = n2331 & n2394;
  assign n2396 = ~n2331 & ~n2394;
  assign n2397 = ~n2395 & ~n2396;
  assign n2398 = n1305 & n2397;
  assign n2399 = n1282_1 & ~n2394;
  assign n2400 = n2321 & ~n2394;
  assign n2401 = ~n2321 & n2394;
  assign n2402 = ~n2400 & ~n2401;
  assign n2403 = n2253 & n2330;
  assign n2404 = n2339 & ~n2403;
  assign n2405 = ~n2253 & ~n2330;
  assign n2406 = n2340 & ~n2403;
  assign n2407 = ~n2065 & n2406;
  assign n2408 = ~n2404 & ~n2405;
  assign n2409 = ~n2407 & n2408;
  assign n2410 = ~n2402 & n2409;
  assign n2411 = n2321 & n2394;
  assign n2412 = ~n2321 & ~n2394;
  assign n2413 = ~n2411 & ~n2412;
  assign n2414 = ~n2409 & ~n2413;
  assign n2415 = ~n2410 & ~n2414;
  assign n2416 = n1318 & ~n2415;
  assign n2417 = ~n2388 & ~n2398;
  assign n2418 = ~n2399 & n2417;
  assign n2419 = ~n2416 & n2418;
  assign n2420 = ~n2343 & ~n2402;
  assign n2421 = ~n2344 & n2354;
  assign n2422 = n2420 & ~n2421;
  assign n2423 = ~n2344 & ~n2401;
  assign n2424 = ~n2400 & n2423;
  assign n2425 = ~n2343 & ~n2354;
  assign n2426 = n2424 & ~n2425;
  assign n2427 = ~n2422 & ~n2426;
  assign n2428 = n1342 & ~n2427;
  assign n2429 = n1390 & ~n2253;
  assign n2430 = n1336 & ~n2415;
  assign n2431 = n1340 & ~n2427;
  assign n2432 = ~n2430 & ~n2431;
  assign n2433 = n1331 & ~n2415;
  assign n2434 = n1325 & ~n2415;
  assign n2435 = n1328 & ~n2427;
  assign n2436 = n1333 & ~n2427;
  assign n2437 = ~n2435 & ~n2436;
  assign n2438 = ~n2433 & ~n2434;
  assign n2439 = n2437 & n2438;
  assign n2440 = ~n2428 & ~n2429;
  assign n2441 = n2432 & n2440;
  assign n2442 = n2439 & n2441;
  assign n2443 = n2419 & n2442;
  assign n2444 = n1268 & ~n2443;
  assign n2445 = REG0_REG_16_ & ~n1268;
  assign n574 = n2444 | n2445;
  assign n2447 = REG3_REG_17_ & REG3_REG_16_;
  assign n2448 = n2311 & n2447;
  assign n2449 = ~REG3_REG_18_ & n2448;
  assign n2450 = REG3_REG_18_ & ~n2448;
  assign n2451 = ~n2449 & ~n2450;
  assign n2452 = n1292_1 & ~n2451;
  assign n2453 = REG0_REG_18_ & n1294;
  assign n2454 = REG1_REG_18_ & n1296;
  assign n2455 = REG2_REG_18_ & n1298;
  assign n2456 = ~n2452 & ~n2453;
  assign n2457 = ~n2454 & n2456;
  assign n2458 = ~n2455 & n2457;
  assign n2459 = n1285 & ~n2458;
  assign n2460 = n2330 & n2394;
  assign n2461 = n2324 & n2460;
  assign n2462 = IR_REG_31_ & n983;
  assign n2463 = IR_REG_17_ & ~IR_REG_31_;
  assign n2464 = ~n2462 & ~n2463;
  assign n2465 = n1275 & ~n2464;
  assign n2466 = DATAI_17_ & ~n1275;
  assign n2467 = ~n2465 & ~n2466;
  assign n2468 = n2461 & n2467;
  assign n2469 = ~n2461 & ~n2467;
  assign n2470 = ~n2468 & ~n2469;
  assign n2471 = n1305 & n2470;
  assign n2472 = n1282_1 & ~n2467;
  assign n2473 = n2387 & n2467;
  assign n2474 = ~n2411 & ~n2473;
  assign n2475 = ~n2387 & ~n2467;
  assign n2476 = n2474 & ~n2475;
  assign n2477 = n2409 & ~n2412;
  assign n2478 = n2476 & ~n2477;
  assign n2479 = n2387 & ~n2467;
  assign n2480 = ~n2387 & n2467;
  assign n2481 = ~n2479 & ~n2480;
  assign n2482 = ~n2412 & n2481;
  assign n2483 = ~n2409 & ~n2411;
  assign n2484 = n2482 & ~n2483;
  assign n2485 = ~n2478 & ~n2484;
  assign n2486 = n1318 & n2485;
  assign n2487 = ~n2459 & ~n2471;
  assign n2488 = ~n2472 & n2487;
  assign n2489 = ~n2486 & n2488;
  assign n2490 = ~n2343 & ~n2400;
  assign n2491 = n2274 & n2490;
  assign n2492 = n2423 & ~n2491;
  assign n2493 = ~n2400 & ~n2492;
  assign n2494 = ~n2273 & n2490;
  assign n2495 = ~n2287 & n2494;
  assign n2496 = ~n2493 & ~n2495;
  assign n2497 = ~n2481 & ~n2496;
  assign n2498 = n2481 & n2496;
  assign n2499 = ~n2497 & ~n2498;
  assign n2500 = n1342 & ~n2499;
  assign n2501 = n1390 & ~n2321;
  assign n2502 = n1336 & n2485;
  assign n2503 = n1340 & ~n2499;
  assign n2504 = ~n2502 & ~n2503;
  assign n2505 = n1331 & n2485;
  assign n2506 = n1325 & n2485;
  assign n2507 = n1328 & ~n2499;
  assign n2508 = n1333 & ~n2499;
  assign n2509 = ~n2507 & ~n2508;
  assign n2510 = ~n2505 & ~n2506;
  assign n2511 = n2509 & n2510;
  assign n2512 = ~n2500 & ~n2501;
  assign n2513 = n2504 & n2512;
  assign n2514 = n2511 & n2513;
  assign n2515 = n2489 & n2514;
  assign n2516 = n1268 & ~n2515;
  assign n2517 = REG0_REG_17_ & ~n1268;
  assign n579 = n2516 | n2517;
  assign n2519 = REG3_REG_18_ & n2448;
  assign n2520 = ~REG3_REG_19_ & n2519;
  assign n2521 = REG3_REG_19_ & ~n2519;
  assign n2522 = ~n2520 & ~n2521;
  assign n2523 = n1292_1 & ~n2522;
  assign n2524 = REG0_REG_19_ & n1294;
  assign n2525 = REG1_REG_19_ & n1296;
  assign n2526 = REG2_REG_19_ & n1298;
  assign n2527 = ~n2523 & ~n2524;
  assign n2528 = ~n2525 & n2527;
  assign n2529 = ~n2526 & n2528;
  assign n2530 = n1285 & ~n2529;
  assign n2531 = IR_REG_31_ & n991;
  assign n2532 = IR_REG_18_ & ~IR_REG_31_;
  assign n2533 = ~n2531 & ~n2532;
  assign n2534 = n1275 & ~n2533;
  assign n2535 = DATAI_18_ & ~n1275;
  assign n2536 = ~n2534 & ~n2535;
  assign n2537 = n2468 & n2536;
  assign n2538 = ~n2468 & ~n2536;
  assign n2539 = ~n2537 & ~n2538;
  assign n2540 = n1305 & n2539;
  assign n2541 = n1282_1 & ~n2536;
  assign n2542 = n2412 & ~n2467;
  assign n2543 = ~n2412 & n2467;
  assign n2544 = ~n2387 & ~n2543;
  assign n2545 = ~n2542 & ~n2544;
  assign n2546 = ~n2409 & n2474;
  assign n2547 = n2545 & ~n2546;
  assign n2548 = n2458 & ~n2536;
  assign n2549 = ~n2458 & n2536;
  assign n2550 = ~n2548 & ~n2549;
  assign n2551 = n2547 & ~n2550;
  assign n2552 = n2458 & n2536;
  assign n2553 = ~n2458 & ~n2536;
  assign n2554 = ~n2552 & ~n2553;
  assign n2555 = ~n2547 & ~n2554;
  assign n2556 = ~n2551 & ~n2555;
  assign n2557 = n1318 & ~n2556;
  assign n2558 = ~n2530 & ~n2540;
  assign n2559 = ~n2541 & n2558;
  assign n2560 = ~n2557 & n2559;
  assign n2561 = ~n2479 & n2493;
  assign n2562 = ~n2480 & ~n2561;
  assign n2563 = ~n2479 & n2494;
  assign n2564 = ~n2287 & n2563;
  assign n2565 = n2562 & ~n2564;
  assign n2566 = ~n2550 & ~n2565;
  assign n2567 = n2550 & n2565;
  assign n2568 = ~n2566 & ~n2567;
  assign n2569 = n1342 & ~n2568;
  assign n2570 = n1390 & ~n2387;
  assign n2571 = n1336 & ~n2556;
  assign n2572 = n1340 & ~n2568;
  assign n2573 = ~n2571 & ~n2572;
  assign n2574 = n1331 & ~n2556;
  assign n2575 = n1325 & ~n2556;
  assign n2576 = n1328 & ~n2568;
  assign n2577 = n1333 & ~n2568;
  assign n2578 = ~n2576 & ~n2577;
  assign n2579 = ~n2574 & ~n2575;
  assign n2580 = n2578 & n2579;
  assign n2581 = ~n2569 & ~n2570;
  assign n2582 = n2573 & n2581;
  assign n2583 = n2580 & n2582;
  assign n2584 = n2560 & n2583;
  assign n2585 = n1268 & ~n2584;
  assign n2586 = REG0_REG_18_ & ~n1268;
  assign n584 = n2585 | n2586;
  assign n2588 = REG3_REG_19_ & n2519;
  assign n2589 = ~REG3_REG_20_ & n2588;
  assign n2590 = REG3_REG_20_ & ~n2588;
  assign n2591 = ~n2589 & ~n2590;
  assign n2592 = n1292_1 & ~n2591;
  assign n2593 = REG0_REG_20_ & n1294;
  assign n2594 = REG1_REG_20_ & n1296;
  assign n2595 = REG2_REG_20_ & n1298;
  assign n2596 = ~n2592 & ~n2593;
  assign n2597 = ~n2594 & n2596;
  assign n2598 = ~n2595 & n2597;
  assign n2599 = n1285 & ~n2598;
  assign n2600 = n2467 & n2536;
  assign n2601 = n2461 & n2600;
  assign n2602 = ~n1193 & n1275;
  assign n2603 = DATAI_19_ & ~n1275;
  assign n2604 = ~n2602 & ~n2603;
  assign n2605 = n2601 & n2604;
  assign n2606 = ~n2601 & ~n2604;
  assign n2607 = ~n2605 & ~n2606;
  assign n2608 = n1305 & n2607;
  assign n2609 = n1282_1 & ~n2604;
  assign n2610 = n2529 & ~n2604;
  assign n2611 = ~n2529 & n2604;
  assign n2612 = ~n2610 & ~n2611;
  assign n2613 = ~n2547 & ~n2552;
  assign n2614 = ~n2553 & ~n2613;
  assign n2615 = ~n2612 & n2614;
  assign n2616 = n2529 & n2604;
  assign n2617 = ~n2529 & ~n2604;
  assign n2618 = ~n2616 & ~n2617;
  assign n2619 = ~n2614 & ~n2618;
  assign n2620 = ~n2615 & ~n2619;
  assign n2621 = n1318 & ~n2620;
  assign n2622 = ~n2599 & ~n2608;
  assign n2623 = ~n2609 & n2622;
  assign n2624 = ~n2621 & n2623;
  assign n2625 = ~n2548 & ~n2565;
  assign n2626 = ~n2549 & ~n2625;
  assign n2627 = ~n2612 & ~n2626;
  assign n2628 = n2612 & n2626;
  assign n2629 = ~n2627 & ~n2628;
  assign n2630 = n1342 & ~n2629;
  assign n2631 = n1390 & ~n2458;
  assign n2632 = n1336 & ~n2620;
  assign n2633 = n1340 & ~n2629;
  assign n2634 = ~n2632 & ~n2633;
  assign n2635 = n1331 & ~n2620;
  assign n2636 = n1325 & ~n2620;
  assign n2637 = n1328 & ~n2629;
  assign n2638 = n1333 & ~n2629;
  assign n2639 = ~n2637 & ~n2638;
  assign n2640 = ~n2635 & ~n2636;
  assign n2641 = n2639 & n2640;
  assign n2642 = ~n2630 & ~n2631;
  assign n2643 = n2634 & n2642;
  assign n2644 = n2641 & n2643;
  assign n2645 = n2624 & n2644;
  assign n2646 = n1268 & ~n2645;
  assign n2647 = REG0_REG_19_ & ~n1268;
  assign n589 = n2646 | n2647;
  assign n2649 = REG1_REG_21_ & n1296;
  assign n2650 = REG0_REG_21_ & n1294;
  assign n2651 = REG2_REG_21_ & n1298;
  assign n2652 = REG3_REG_20_ & n2588;
  assign n2653 = ~REG3_REG_21_ & n2652;
  assign n2654 = REG3_REG_21_ & ~n2652;
  assign n2655 = ~n2653 & ~n2654;
  assign n2656 = n1292_1 & ~n2655;
  assign n2657 = ~n2649 & ~n2650;
  assign n2658 = ~n2651 & n2657;
  assign n2659 = ~n2656 & n2658;
  assign n2660 = n1285 & ~n2659;
  assign n2661 = DATAI_20_ & ~n1275;
  assign n2662 = n2605 & ~n2661;
  assign n2663 = ~n2605 & n2661;
  assign n2664 = ~n2662 & ~n2663;
  assign n2665 = n1305 & n2664;
  assign n2666 = n1282_1 & n2661;
  assign n2667 = ~n2598 & n2661;
  assign n2668 = n2598 & ~n2661;
  assign n2669 = ~n2616 & ~n2668;
  assign n2670 = ~n2667 & n2669;
  assign n2671 = n2614 & ~n2617;
  assign n2672 = n2670 & ~n2671;
  assign n2673 = n2598 & n2661;
  assign n2674 = ~n2598 & ~n2661;
  assign n2675 = ~n2673 & ~n2674;
  assign n2676 = ~n2617 & n2675;
  assign n2677 = ~n2614 & ~n2616;
  assign n2678 = n2676 & ~n2677;
  assign n2679 = ~n2672 & ~n2678;
  assign n2680 = n1318 & n2679;
  assign n2681 = ~n2660 & ~n2665;
  assign n2682 = ~n2666 & n2681;
  assign n2683 = ~n2680 & n2682;
  assign n2684 = ~n2610 & ~n2626;
  assign n2685 = ~n2611 & ~n2684;
  assign n2686 = ~n2675 & ~n2685;
  assign n2687 = n2675 & n2685;
  assign n2688 = ~n2686 & ~n2687;
  assign n2689 = n1342 & ~n2688;
  assign n2690 = n1390 & ~n2529;
  assign n2691 = n1336 & n2679;
  assign n2692 = n1340 & ~n2688;
  assign n2693 = ~n2691 & ~n2692;
  assign n2694 = n1331 & n2679;
  assign n2695 = n1325 & n2679;
  assign n2696 = n1328 & ~n2688;
  assign n2697 = n1333 & ~n2688;
  assign n2698 = ~n2696 & ~n2697;
  assign n2699 = ~n2694 & ~n2695;
  assign n2700 = n2698 & n2699;
  assign n2701 = ~n2689 & ~n2690;
  assign n2702 = n2693 & n2701;
  assign n2703 = n2700 & n2702;
  assign n2704 = n2683 & n2703;
  assign n2705 = n1268 & ~n2704;
  assign n2706 = REG0_REG_20_ & ~n1268;
  assign n594 = n2705 | n2706;
  assign n2708 = REG1_REG_22_ & n1296;
  assign n2709 = REG0_REG_22_ & n1294;
  assign n2710 = REG2_REG_22_ & n1298;
  assign n2711 = REG3_REG_21_ & n2652;
  assign n2712 = ~REG3_REG_22_ & n2711;
  assign n2713 = REG3_REG_22_ & ~n2711;
  assign n2714 = ~n2712 & ~n2713;
  assign n2715 = n1292_1 & ~n2714;
  assign n2716 = ~n2708 & ~n2709;
  assign n2717 = ~n2710 & n2716;
  assign n2718 = ~n2715 & n2717;
  assign n2719 = n1285 & ~n2718;
  assign n2720 = n2604 & ~n2661;
  assign n2721 = n2601 & n2720;
  assign n2722 = DATAI_21_ & ~n1275;
  assign n2723 = n2721 & ~n2722;
  assign n2724 = ~n2721 & n2722;
  assign n2725 = ~n2723 & ~n2724;
  assign n2726 = n1305 & n2725;
  assign n2727 = n1282_1 & n2722;
  assign n2728 = n2659 & n2722;
  assign n2729 = ~n2659 & ~n2722;
  assign n2730 = ~n2728 & ~n2729;
  assign n2731 = ~n2614 & n2669;
  assign n2732 = ~n2617 & ~n2661;
  assign n2733 = n2617 & n2661;
  assign n2734 = n2598 & ~n2733;
  assign n2735 = ~n2732 & ~n2734;
  assign n2736 = ~n2731 & ~n2735;
  assign n2737 = ~n2730 & ~n2736;
  assign n2738 = n2730 & ~n2735;
  assign n2739 = ~n2731 & n2738;
  assign n2740 = ~n2737 & ~n2739;
  assign n2741 = n1318 & n2740;
  assign n2742 = ~n2719 & ~n2726;
  assign n2743 = ~n2727 & n2742;
  assign n2744 = ~n2741 & n2743;
  assign n2745 = n2611 & ~n2673;
  assign n2746 = ~n2674 & ~n2745;
  assign n2747 = ~n2610 & ~n2673;
  assign n2748 = ~n2626 & n2747;
  assign n2749 = n2746 & ~n2748;
  assign n2750 = n2730 & n2749;
  assign n2751 = ~n2730 & ~n2749;
  assign n2752 = ~n2750 & ~n2751;
  assign n2753 = n1342 & ~n2752;
  assign n2754 = n1390 & ~n2598;
  assign n2755 = n1336 & n2740;
  assign n2756 = n1340 & ~n2752;
  assign n2757 = ~n2755 & ~n2756;
  assign n2758 = n1331 & n2740;
  assign n2759 = n1325 & n2740;
  assign n2760 = n1328 & ~n2752;
  assign n2761 = n1333 & ~n2752;
  assign n2762 = ~n2760 & ~n2761;
  assign n2763 = ~n2758 & ~n2759;
  assign n2764 = n2762 & n2763;
  assign n2765 = ~n2753 & ~n2754;
  assign n2766 = n2757 & n2765;
  assign n2767 = n2764 & n2766;
  assign n2768 = n2744 & n2767;
  assign n2769 = n1268 & ~n2768;
  assign n2770 = REG0_REG_21_ & ~n1268;
  assign n599 = n2769 | n2770;
  assign n2772 = REG1_REG_23_ & n1296;
  assign n2773 = REG0_REG_23_ & n1294;
  assign n2774 = REG2_REG_23_ & n1298;
  assign n2775 = REG3_REG_22_ & n2711;
  assign n2776 = ~REG3_REG_23_ & n2775;
  assign n2777 = REG3_REG_23_ & ~n2775;
  assign n2778 = ~n2776 & ~n2777;
  assign n2779 = n1292_1 & ~n2778;
  assign n2780 = ~n2772 & ~n2773;
  assign n2781 = ~n2774 & n2780;
  assign n2782 = ~n2779 & n2781;
  assign n2783 = n1285 & ~n2782;
  assign n2784 = DATAI_22_ & ~n1275;
  assign n2785 = n2723 & ~n2784;
  assign n2786 = ~n2723 & n2784;
  assign n2787 = ~n2785 & ~n2786;
  assign n2788 = n1305 & n2787;
  assign n2789 = n1282_1 & n2784;
  assign n2790 = n2659 & ~n2722;
  assign n2791 = n2669 & ~n2790;
  assign n2792 = ~n2552 & n2791;
  assign n2793 = ~n2545 & n2792;
  assign n2794 = n2553 & n2791;
  assign n2795 = ~n2659 & n2722;
  assign n2796 = ~n2735 & ~n2794;
  assign n2797 = ~n2795 & n2796;
  assign n2798 = ~n2790 & ~n2797;
  assign n2799 = ~n2793 & ~n2798;
  assign n2800 = n2474 & n2792;
  assign n2801 = ~n2409 & n2800;
  assign n2802 = n2799 & ~n2801;
  assign n2803 = n2718 & n2784;
  assign n2804 = ~n2718 & ~n2784;
  assign n2805 = ~n2803 & ~n2804;
  assign n2806 = n2802 & ~n2805;
  assign n2807 = ~n2802 & n2805;
  assign n2808 = ~n2806 & ~n2807;
  assign n2809 = n1318 & ~n2808;
  assign n2810 = ~n2783 & ~n2788;
  assign n2811 = ~n2789 & n2810;
  assign n2812 = ~n2809 & n2811;
  assign n2813 = ~n2728 & ~n2749;
  assign n2814 = ~n2729 & ~n2813;
  assign n2815 = n2805 & n2814;
  assign n2816 = ~n2805 & ~n2814;
  assign n2817 = ~n2815 & ~n2816;
  assign n2818 = n1342 & ~n2817;
  assign n2819 = n1390 & ~n2659;
  assign n2820 = n1336 & ~n2808;
  assign n2821 = ~n2728 & ~n2746;
  assign n2822 = ~n2729 & ~n2821;
  assign n2823 = ~n2728 & n2747;
  assign n2824 = ~n2626 & n2823;
  assign n2825 = n2822 & ~n2824;
  assign n2826 = n2805 & n2825;
  assign n2827 = ~n2805 & ~n2825;
  assign n2828 = ~n2826 & ~n2827;
  assign n2829 = n1340 & ~n2828;
  assign n2830 = ~n2820 & ~n2829;
  assign n2831 = n1331 & ~n2808;
  assign n2832 = n1325 & ~n2808;
  assign n2833 = n1328 & ~n2817;
  assign n2834 = n1333 & ~n2817;
  assign n2835 = ~n2833 & ~n2834;
  assign n2836 = ~n2831 & ~n2832;
  assign n2837 = n2835 & n2836;
  assign n2838 = ~n2818 & ~n2819;
  assign n2839 = n2830 & n2838;
  assign n2840 = n2837 & n2839;
  assign n2841 = n2812 & n2840;
  assign n2842 = n1268 & ~n2841;
  assign n2843 = REG0_REG_22_ & ~n1268;
  assign n604 = n2842 | n2843;
  assign n2845 = REG1_REG_24_ & n1296;
  assign n2846 = REG0_REG_24_ & n1294;
  assign n2847 = REG2_REG_24_ & n1298;
  assign n2848 = REG3_REG_23_ & n2775;
  assign n2849 = ~REG3_REG_24_ & n2848;
  assign n2850 = REG3_REG_24_ & ~n2848;
  assign n2851 = ~n2849 & ~n2850;
  assign n2852 = n1292_1 & ~n2851;
  assign n2853 = ~n2845 & ~n2846;
  assign n2854 = ~n2847 & n2853;
  assign n2855 = ~n2852 & n2854;
  assign n2856 = n1285 & ~n2855;
  assign n2857 = ~n2722 & ~n2784;
  assign n2858 = n2721 & n2857;
  assign n2859 = DATAI_23_ & ~n1275;
  assign n2860 = n2858 & ~n2859;
  assign n2861 = ~n2858 & n2859;
  assign n2862 = ~n2860 & ~n2861;
  assign n2863 = n1305 & n2862;
  assign n2864 = n1282_1 & n2859;
  assign n2865 = ~n2718 & n2784;
  assign n2866 = n2718 & ~n2784;
  assign n2867 = ~n2802 & ~n2866;
  assign n2868 = ~n2865 & ~n2867;
  assign n2869 = n2782 & n2859;
  assign n2870 = ~n2782 & ~n2859;
  assign n2871 = ~n2869 & ~n2870;
  assign n2872 = n2868 & ~n2871;
  assign n2873 = ~n2868 & n2871;
  assign n2874 = ~n2872 & ~n2873;
  assign n2875 = n1318 & ~n2874;
  assign n2876 = ~n2856 & ~n2863;
  assign n2877 = ~n2864 & n2876;
  assign n2878 = ~n2875 & n2877;
  assign n2879 = ~n2803 & ~n2871;
  assign n2880 = ~n2804 & n2814;
  assign n2881 = n2879 & ~n2880;
  assign n2882 = ~n2804 & ~n2870;
  assign n2883 = ~n2869 & n2882;
  assign n2884 = ~n2803 & ~n2814;
  assign n2885 = n2883 & ~n2884;
  assign n2886 = ~n2881 & ~n2885;
  assign n2887 = n1342 & ~n2886;
  assign n2888 = n1390 & ~n2718;
  assign n2889 = ~n2799 & ~n2866;
  assign n2890 = ~n2865 & ~n2889;
  assign n2891 = n2800 & ~n2866;
  assign n2892 = ~n2409 & n2891;
  assign n2893 = n2890 & ~n2892;
  assign n2894 = ~n2871 & n2893;
  assign n2895 = n2871 & ~n2893;
  assign n2896 = ~n2894 & ~n2895;
  assign n2897 = n1336 & ~n2896;
  assign n2898 = n2825 & n2883;
  assign n2899 = n2804 & ~n2871;
  assign n2900 = n2803 & n2883;
  assign n2901 = ~n2825 & ~n2871;
  assign n2902 = ~n2803 & n2901;
  assign n2903 = ~n2898 & ~n2899;
  assign n2904 = ~n2900 & n2903;
  assign n2905 = ~n2902 & n2904;
  assign n2906 = n1340 & ~n2905;
  assign n2907 = ~n2897 & ~n2906;
  assign n2908 = n1331 & ~n2896;
  assign n2909 = n1325 & ~n2896;
  assign n2910 = n2729 & n2879;
  assign n2911 = ~n2821 & ~n2869;
  assign n2912 = n2882 & n2911;
  assign n2913 = ~n2824 & n2912;
  assign n2914 = ~n2729 & n2913;
  assign n2915 = n2803 & ~n2869;
  assign n2916 = n2882 & n2915;
  assign n2917 = ~n2728 & n2879;
  assign n2918 = ~n2749 & n2917;
  assign n2919 = ~n2910 & ~n2914;
  assign n2920 = ~n2899 & n2919;
  assign n2921 = ~n2916 & n2920;
  assign n2922 = ~n2918 & n2921;
  assign n2923 = n1328 & ~n2922;
  assign n2924 = n1333 & ~n2922;
  assign n2925 = ~n2923 & ~n2924;
  assign n2926 = ~n2908 & ~n2909;
  assign n2927 = n2925 & n2926;
  assign n2928 = ~n2887 & ~n2888;
  assign n2929 = n2907 & n2928;
  assign n2930 = n2927 & n2929;
  assign n2931 = n2878 & n2930;
  assign n2932 = n1268 & ~n2931;
  assign n2933 = REG0_REG_23_ & ~n1268;
  assign n609 = n2932 | n2933;
  assign n2935 = REG1_REG_25_ & n1296;
  assign n2936 = REG0_REG_25_ & n1294;
  assign n2937 = REG2_REG_25_ & n1298;
  assign n2938 = REG3_REG_24_ & n2848;
  assign n2939 = ~REG3_REG_25_ & n2938;
  assign n2940 = REG3_REG_25_ & ~n2938;
  assign n2941 = ~n2939 & ~n2940;
  assign n2942 = n1292_1 & ~n2941;
  assign n2943 = ~n2935 & ~n2936;
  assign n2944 = ~n2937 & n2943;
  assign n2945 = ~n2942 & n2944;
  assign n2946 = n1285 & ~n2945;
  assign n2947 = DATAI_24_ & ~n1275;
  assign n2948 = n2860 & ~n2947;
  assign n2949 = ~n2860 & n2947;
  assign n2950 = ~n2948 & ~n2949;
  assign n2951 = n1305 & n2950;
  assign n2952 = n1282_1 & n2947;
  assign n2953 = ~n2782 & n2859;
  assign n2954 = n2782 & ~n2859;
  assign n2955 = ~n2868 & ~n2954;
  assign n2956 = ~n2953 & ~n2955;
  assign n2957 = n2855 & n2947;
  assign n2958 = ~n2855 & ~n2947;
  assign n2959 = ~n2957 & ~n2958;
  assign n2960 = n2956 & ~n2959;
  assign n2961 = n2855 & ~n2947;
  assign n2962 = ~n2855 & n2947;
  assign n2963 = ~n2961 & ~n2962;
  assign n2964 = ~n2956 & ~n2963;
  assign n2965 = ~n2960 & ~n2964;
  assign n2966 = n1318 & ~n2965;
  assign n2967 = ~n2946 & ~n2951;
  assign n2968 = ~n2952 & n2967;
  assign n2969 = ~n2966 & n2968;
  assign n2970 = ~n2803 & ~n2869;
  assign n2971 = ~n2728 & n2970;
  assign n2972 = ~n2746 & n2971;
  assign n2973 = n2729 & n2970;
  assign n2974 = n2882 & ~n2973;
  assign n2975 = ~n2869 & ~n2974;
  assign n2976 = ~n2972 & ~n2975;
  assign n2977 = n2747 & n2971;
  assign n2978 = ~n2626 & n2977;
  assign n2979 = n2976 & ~n2978;
  assign n2980 = ~n2959 & ~n2979;
  assign n2981 = n2959 & n2979;
  assign n2982 = ~n2980 & ~n2981;
  assign n2983 = n1342 & ~n2982;
  assign n2984 = n1390 & ~n2782;
  assign n2985 = ~n2893 & ~n2954;
  assign n2986 = ~n2953 & ~n2985;
  assign n2987 = ~n2959 & n2986;
  assign n2988 = ~n2963 & ~n2986;
  assign n2989 = ~n2987 & ~n2988;
  assign n2990 = n1336 & ~n2989;
  assign n2991 = n1340 & ~n2982;
  assign n2992 = ~n2990 & ~n2991;
  assign n2993 = n1331 & ~n2989;
  assign n2994 = n1325 & ~n2989;
  assign n2995 = n1328 & ~n2982;
  assign n2996 = n1333 & ~n2982;
  assign n2997 = ~n2995 & ~n2996;
  assign n2998 = ~n2993 & ~n2994;
  assign n2999 = n2997 & n2998;
  assign n3000 = ~n2983 & ~n2984;
  assign n3001 = n2992 & n3000;
  assign n3002 = n2999 & n3001;
  assign n3003 = n2969 & n3002;
  assign n3004 = n1268 & ~n3003;
  assign n3005 = REG0_REG_24_ & ~n1268;
  assign n614 = n3004 | n3005;
  assign n3007 = REG1_REG_26_ & n1296;
  assign n3008 = REG0_REG_26_ & n1294;
  assign n3009 = REG2_REG_26_ & n1298;
  assign n3010 = REG3_REG_25_ & n2938;
  assign n3011 = ~REG3_REG_26_ & n3010;
  assign n3012 = REG3_REG_26_ & ~n3010;
  assign n3013 = ~n3011 & ~n3012;
  assign n3014 = n1292_1 & ~n3013;
  assign n3015 = ~n3007 & ~n3008;
  assign n3016 = ~n3009 & n3015;
  assign n3017 = ~n3014 & n3016;
  assign n3018 = n1285 & ~n3017;
  assign n3019 = ~n2859 & ~n2947;
  assign n3020 = n2858 & n3019;
  assign n3021 = DATAI_25_ & ~n1275;
  assign n3022 = n3020 & ~n3021;
  assign n3023 = ~n3020 & n3021;
  assign n3024 = ~n3022 & ~n3023;
  assign n3025 = n1305 & n3024;
  assign n3026 = n1282_1 & n3021;
  assign n3027 = n2945 & n3021;
  assign n3028 = ~n2945 & ~n3021;
  assign n3029 = ~n3027 & ~n3028;
  assign n3030 = ~n2956 & ~n2961;
  assign n3031 = ~n2962 & ~n3030;
  assign n3032 = ~n3029 & n3031;
  assign n3033 = n2945 & ~n3021;
  assign n3034 = ~n2945 & n3021;
  assign n3035 = ~n3033 & ~n3034;
  assign n3036 = ~n3031 & ~n3035;
  assign n3037 = ~n3032 & ~n3036;
  assign n3038 = n1318 & ~n3037;
  assign n3039 = ~n3018 & ~n3025;
  assign n3040 = ~n3026 & n3039;
  assign n3041 = ~n3038 & n3040;
  assign n3042 = ~n2957 & ~n2976;
  assign n3043 = ~n2958 & ~n3042;
  assign n3044 = ~n2957 & n2977;
  assign n3045 = ~n2626 & n3044;
  assign n3046 = n3043 & ~n3045;
  assign n3047 = ~n3029 & ~n3046;
  assign n3048 = n3029 & n3046;
  assign n3049 = ~n3047 & ~n3048;
  assign n3050 = n1342 & ~n3049;
  assign n3051 = n1390 & ~n2855;
  assign n3052 = ~n2961 & ~n2986;
  assign n3053 = ~n2962 & ~n3052;
  assign n3054 = ~n3029 & n3053;
  assign n3055 = ~n3035 & ~n3053;
  assign n3056 = ~n3054 & ~n3055;
  assign n3057 = n1336 & ~n3056;
  assign n3058 = n1340 & ~n3049;
  assign n3059 = ~n3057 & ~n3058;
  assign n3060 = n1331 & ~n3056;
  assign n3061 = n1325 & ~n3056;
  assign n3062 = n1328 & ~n3049;
  assign n3063 = n1333 & ~n3049;
  assign n3064 = ~n3062 & ~n3063;
  assign n3065 = ~n3060 & ~n3061;
  assign n3066 = n3064 & n3065;
  assign n3067 = ~n3050 & ~n3051;
  assign n3068 = n3059 & n3067;
  assign n3069 = n3066 & n3068;
  assign n3070 = n3041 & n3069;
  assign n3071 = n1268 & ~n3070;
  assign n3072 = REG0_REG_25_ & ~n1268;
  assign n619 = n3071 | n3072;
  assign n3074 = REG1_REG_27_ & n1296;
  assign n3075 = REG0_REG_27_ & n1294;
  assign n3076 = REG2_REG_27_ & n1298;
  assign n3077 = REG3_REG_26_ & n3010;
  assign n3078 = ~REG3_REG_27_ & n3077;
  assign n3079 = REG3_REG_27_ & ~n3077;
  assign n3080 = ~n3078 & ~n3079;
  assign n3081 = n1292_1 & ~n3080;
  assign n3082 = ~n3074 & ~n3075;
  assign n3083 = ~n3076 & n3082;
  assign n3084 = ~n3081 & n3083;
  assign n3085 = n1285 & ~n3084;
  assign n3086 = DATAI_26_ & ~n1275;
  assign n3087 = n3022 & ~n3086;
  assign n3088 = ~n3022 & n3086;
  assign n3089 = ~n3087 & ~n3088;
  assign n3090 = n1305 & n3089;
  assign n3091 = n1282_1 & n3086;
  assign n3092 = ~n3017 & n3086;
  assign n3093 = n3017 & ~n3086;
  assign n3094 = ~n3033 & ~n3093;
  assign n3095 = ~n3092 & n3094;
  assign n3096 = n3031 & ~n3034;
  assign n3097 = n3095 & ~n3096;
  assign n3098 = n3017 & n3086;
  assign n3099 = ~n3017 & ~n3086;
  assign n3100 = ~n3098 & ~n3099;
  assign n3101 = ~n3034 & n3100;
  assign n3102 = ~n3031 & ~n3033;
  assign n3103 = n3101 & ~n3102;
  assign n3104 = ~n3097 & ~n3103;
  assign n3105 = n1318 & n3104;
  assign n3106 = ~n3085 & ~n3090;
  assign n3107 = ~n3091 & n3106;
  assign n3108 = ~n3105 & n3107;
  assign n3109 = ~n3027 & ~n3043;
  assign n3110 = ~n3028 & ~n3109;
  assign n3111 = ~n3027 & n3044;
  assign n3112 = ~n2626 & n3111;
  assign n3113 = n3110 & ~n3112;
  assign n3114 = n3100 & n3113;
  assign n3115 = ~n3100 & ~n3113;
  assign n3116 = ~n3114 & ~n3115;
  assign n3117 = n1342 & ~n3116;
  assign n3118 = n1390 & ~n2945;
  assign n3119 = ~n3033 & n3086;
  assign n3120 = ~n3017 & ~n3033;
  assign n3121 = ~n3119 & ~n3120;
  assign n3122 = ~n3092 & ~n3121;
  assign n3123 = ~n3034 & n3053;
  assign n3124 = n3122 & ~n3123;
  assign n3125 = ~n3033 & ~n3053;
  assign n3126 = n3101 & ~n3125;
  assign n3127 = ~n3124 & ~n3126;
  assign n3128 = n1336 & n3127;
  assign n3129 = ~n3027 & ~n3046;
  assign n3130 = ~n3028 & ~n3129;
  assign n3131 = n3100 & n3130;
  assign n3132 = ~n3100 & ~n3130;
  assign n3133 = ~n3131 & ~n3132;
  assign n3134 = n1340 & ~n3133;
  assign n3135 = ~n3128 & ~n3134;
  assign n3136 = n1331 & n3127;
  assign n3137 = n1325 & n3127;
  assign n3138 = n1328 & ~n3116;
  assign n3139 = n1333 & ~n3116;
  assign n3140 = ~n3138 & ~n3139;
  assign n3141 = ~n3136 & ~n3137;
  assign n3142 = n3140 & n3141;
  assign n3143 = ~n3117 & ~n3118;
  assign n3144 = n3135 & n3143;
  assign n3145 = n3142 & n3144;
  assign n3146 = n3108 & n3145;
  assign n3147 = n1268 & ~n3146;
  assign n3148 = REG0_REG_26_ & ~n1268;
  assign n624 = n3147 | n3148;
  assign n3150 = REG1_REG_28_ & n1296;
  assign n3151 = REG0_REG_28_ & n1294;
  assign n3152 = REG2_REG_28_ & n1298;
  assign n3153 = REG3_REG_27_ & n3077;
  assign n3154 = ~REG3_REG_28_ & n3153;
  assign n3155 = REG3_REG_28_ & ~n3153;
  assign n3156 = ~n3154 & ~n3155;
  assign n3157 = n1292_1 & ~n3156;
  assign n3158 = ~n3150 & ~n3151;
  assign n3159 = ~n3152 & n3158;
  assign n3160 = ~n3157 & n3159;
  assign n3161 = n1285 & ~n3160;
  assign n3162 = ~n3021 & ~n3086;
  assign n3163 = n3020 & n3162;
  assign n3164 = DATAI_27_ & ~n1275;
  assign n3165 = n3163 & ~n3164;
  assign n3166 = ~n3163 & n3164;
  assign n3167 = ~n3165 & ~n3166;
  assign n3168 = n1305 & n3167;
  assign n3169 = n1282_1 & n3164;
  assign n3170 = ~n3034 & ~n3092;
  assign n3171 = n2962 & n3094;
  assign n3172 = n3170 & ~n3171;
  assign n3173 = ~n3093 & ~n3172;
  assign n3174 = ~n2961 & n3094;
  assign n3175 = ~n2956 & n3174;
  assign n3176 = ~n3173 & ~n3175;
  assign n3177 = n3084 & n3164;
  assign n3178 = ~n3084 & ~n3164;
  assign n3179 = ~n3177 & ~n3178;
  assign n3180 = n3176 & ~n3179;
  assign n3181 = ~n3176 & n3179;
  assign n3182 = ~n3180 & ~n3181;
  assign n3183 = n1318 & ~n3182;
  assign n3184 = ~n3161 & ~n3168;
  assign n3185 = ~n3169 & n3184;
  assign n3186 = ~n3183 & n3185;
  assign n3187 = ~n3098 & ~n3179;
  assign n3188 = ~n3099 & n3113;
  assign n3189 = n3187 & ~n3188;
  assign n3190 = ~n3099 & n3179;
  assign n3191 = ~n3098 & ~n3113;
  assign n3192 = n3190 & ~n3191;
  assign n3193 = ~n3189 & ~n3192;
  assign n3194 = n1342 & ~n3193;
  assign n3195 = n1390 & ~n3017;
  assign n3196 = ~n3034 & ~n3086;
  assign n3197 = n3017 & ~n3034;
  assign n3198 = ~n3093 & ~n3196;
  assign n3199 = ~n3197 & n3198;
  assign n3200 = n2962 & ~n3121;
  assign n3201 = ~n3199 & ~n3200;
  assign n3202 = ~n2954 & ~n2961;
  assign n3203 = ~n3121 & n3202;
  assign n3204 = n2893 & ~n2953;
  assign n3205 = n3203 & ~n3204;
  assign n3206 = n3201 & ~n3205;
  assign n3207 = ~n3179 & n3206;
  assign n3208 = n3179 & ~n3206;
  assign n3209 = ~n3207 & ~n3208;
  assign n3210 = n1336 & ~n3209;
  assign n3211 = ~n3098 & ~n3187;
  assign n3212 = ~n3130 & n3211;
  assign n3213 = n3099 & ~n3179;
  assign n3214 = ~n3190 & ~n3213;
  assign n3215 = ~n3130 & n3187;
  assign n3216 = n3214 & ~n3215;
  assign n3217 = ~n3212 & ~n3216;
  assign n3218 = n1340 & n3217;
  assign n3219 = ~n3210 & ~n3218;
  assign n3220 = n1331 & ~n3209;
  assign n3221 = n1325 & ~n3209;
  assign n3222 = ~n3113 & n3187;
  assign n3223 = n3214 & ~n3222;
  assign n3224 = n3191 & ~n3222;
  assign n3225 = ~n3223 & ~n3224;
  assign n3226 = n1328 & n3225;
  assign n3227 = n1333 & n3225;
  assign n3228 = ~n3226 & ~n3227;
  assign n3229 = ~n3220 & ~n3221;
  assign n3230 = n3228 & n3229;
  assign n3231 = ~n3194 & ~n3195;
  assign n3232 = n3219 & n3231;
  assign n3233 = n3230 & n3232;
  assign n3234 = n3186 & n3233;
  assign n3235 = n1268 & ~n3234;
  assign n3236 = REG0_REG_27_ & ~n1268;
  assign n629 = n3235 | n3236;
  assign n3238 = REG0_REG_29_ & n1294;
  assign n3239 = REG1_REG_29_ & n1296;
  assign n3240 = REG2_REG_29_ & n1298;
  assign n3241 = REG3_REG_28_ & REG3_REG_27_;
  assign n3242 = n3077 & n3241;
  assign n3243 = n1292_1 & n3242;
  assign n3244 = ~n3238 & ~n3239;
  assign n3245 = ~n3240 & n3244;
  assign n3246 = ~n3243 & n3245;
  assign n3247 = n1285 & ~n3246;
  assign n3248 = DATAI_28_ & ~n1275;
  assign n3249 = n3165 & ~n3248;
  assign n3250 = ~n3165 & n3248;
  assign n3251 = ~n3249 & ~n3250;
  assign n3252 = n1305 & n3251;
  assign n3253 = n1282_1 & n3248;
  assign n3254 = ~n3084 & n3164;
  assign n3255 = n3084 & ~n3164;
  assign n3256 = ~n3176 & ~n3255;
  assign n3257 = ~n3254 & ~n3256;
  assign n3258 = n3160 & n3248;
  assign n3259 = ~n3160 & ~n3248;
  assign n3260 = ~n3258 & ~n3259;
  assign n3261 = n3257 & ~n3260;
  assign n3262 = ~n3257 & n3260;
  assign n3263 = ~n3261 & ~n3262;
  assign n3264 = n1318 & ~n3263;
  assign n3265 = ~n3247 & ~n3252;
  assign n3266 = ~n3253 & n3265;
  assign n3267 = ~n3264 & n3266;
  assign n3268 = n3084 & ~n3099;
  assign n3269 = ~n3164 & ~n3268;
  assign n3270 = ~n3084 & n3099;
  assign n3271 = ~n3269 & ~n3270;
  assign n3272 = ~n3098 & ~n3177;
  assign n3273 = ~n3113 & n3272;
  assign n3274 = n3271 & ~n3273;
  assign n3275 = ~n3260 & ~n3274;
  assign n3276 = n3260 & n3274;
  assign n3277 = ~n3275 & ~n3276;
  assign n3278 = n1342 & ~n3277;
  assign n3279 = n1390 & ~n3084;
  assign n3280 = n3200 & ~n3255;
  assign n3281 = n3199 & ~n3255;
  assign n3282 = ~n3254 & ~n3280;
  assign n3283 = ~n3281 & n3282;
  assign n3284 = ~n3121 & ~n3255;
  assign n3285 = n3202 & ~n3204;
  assign n3286 = n3284 & n3285;
  assign n3287 = n3283 & ~n3286;
  assign n3288 = ~n3260 & n3287;
  assign n3289 = n3260 & ~n3287;
  assign n3290 = ~n3288 & ~n3289;
  assign n3291 = n1336 & ~n3290;
  assign n3292 = ~n3130 & n3272;
  assign n3293 = n3271 & ~n3292;
  assign n3294 = ~n3260 & ~n3293;
  assign n3295 = n3260 & n3293;
  assign n3296 = ~n3294 & ~n3295;
  assign n3297 = n1340 & ~n3296;
  assign n3298 = ~n3291 & ~n3297;
  assign n3299 = n1331 & ~n3290;
  assign n3300 = n1325 & ~n3290;
  assign n3301 = n1328 & ~n3277;
  assign n3302 = n1333 & ~n3277;
  assign n3303 = ~n3301 & ~n3302;
  assign n3304 = ~n3299 & ~n3300;
  assign n3305 = n3303 & n3304;
  assign n3306 = ~n3278 & ~n3279;
  assign n3307 = n3298 & n3306;
  assign n3308 = n3305 & n3307;
  assign n3309 = n3267 & n3308;
  assign n3310 = n1268 & ~n3309;
  assign n3311 = REG0_REG_28_ & ~n1268;
  assign n634 = n3310 | n3311;
  assign n3313 = ~n3164 & ~n3248;
  assign n3314 = n3163 & n3313;
  assign n3315 = DATAI_29_ & ~n1275;
  assign n3316 = n3314 & ~n3315;
  assign n3317 = ~n3314 & n3315;
  assign n3318 = ~n3316 & ~n3317;
  assign n3319 = n1305 & n3318;
  assign n3320 = n1282_1 & n3315;
  assign n3321 = n3248 & ~n3257;
  assign n3322 = ~n3160 & ~n3257;
  assign n3323 = ~n3160 & n3248;
  assign n3324 = ~n3321 & ~n3322;
  assign n3325 = ~n3323 & n3324;
  assign n3326 = n3246 & n3315;
  assign n3327 = ~n3246 & ~n3315;
  assign n3328 = ~n3326 & ~n3327;
  assign n3329 = n3325 & ~n3328;
  assign n3330 = ~n3325 & n3328;
  assign n3331 = ~n3329 & ~n3330;
  assign n3332 = n1318 & ~n3331;
  assign n3333 = ~n3319 & ~n3320;
  assign n3334 = ~n3332 & n3333;
  assign n3335 = n1390 & ~n3160;
  assign n3336 = ~B_REG & n1274;
  assign n3337 = ~n1275 & ~n3336;
  assign n3338 = n1284 & ~n3337;
  assign n3339 = REG1_REG_30_ & n1296;
  assign n3340 = REG0_REG_30_ & n1294;
  assign n3341 = REG2_REG_30_ & n1298;
  assign n3342 = ~n3339 & ~n3340;
  assign n3343 = ~n3341 & n3342;
  assign n3344 = n3338 & ~n3343;
  assign n3345 = n3248 & ~n3287;
  assign n3346 = ~n3160 & ~n3287;
  assign n3347 = ~n3345 & ~n3346;
  assign n3348 = ~n3323 & n3347;
  assign n3349 = ~n3328 & n3348;
  assign n3350 = n3328 & ~n3348;
  assign n3351 = ~n3349 & ~n3350;
  assign n3352 = n1336 & ~n3351;
  assign n3353 = n1331 & ~n3351;
  assign n3354 = n1325 & ~n3351;
  assign n3355 = ~n3335 & ~n3344;
  assign n3356 = ~n3352 & n3355;
  assign n3357 = ~n3353 & n3356;
  assign n3358 = ~n3354 & n3357;
  assign n3359 = ~n3248 & ~n3328;
  assign n3360 = ~n3160 & n3359;
  assign n3361 = n3248 & n3328;
  assign n3362 = n3160 & n3361;
  assign n3363 = ~n3360 & ~n3362;
  assign n3364 = ~n3258 & ~n3328;
  assign n3365 = ~n3274 & n3364;
  assign n3366 = ~n3259 & n3328;
  assign n3367 = n3274 & n3366;
  assign n3368 = n3363 & ~n3365;
  assign n3369 = ~n3367 & n3368;
  assign n3370 = n1328 & ~n3369;
  assign n3371 = n1333 & ~n3369;
  assign n3372 = ~n3270 & n3328;
  assign n3373 = ~n3269 & n3372;
  assign n3374 = ~n3259 & n3373;
  assign n3375 = ~n3292 & n3374;
  assign n3376 = n3160 & n3328;
  assign n3377 = n3248 & n3376;
  assign n3378 = ~n3160 & ~n3328;
  assign n3379 = ~n3248 & n3378;
  assign n3380 = ~n3377 & ~n3379;
  assign n3381 = ~n3375 & n3380;
  assign n3382 = ~n3293 & n3364;
  assign n3383 = n3381 & ~n3382;
  assign n3384 = n1340 & ~n3383;
  assign n3385 = ~n3365 & n3380;
  assign n3386 = ~n3367 & n3385;
  assign n3387 = n1342 & ~n3386;
  assign n3388 = ~n3370 & ~n3371;
  assign n3389 = ~n3384 & n3388;
  assign n3390 = ~n3387 & n3389;
  assign n3391 = n3334 & n3358;
  assign n3392 = n3390 & n3391;
  assign n3393 = n1268 & ~n3392;
  assign n3394 = REG0_REG_29_ & ~n1268;
  assign n639 = n3393 | n3394;
  assign n3396 = DATAI_30_ & ~n1275;
  assign n3397 = n1282_1 & n3396;
  assign n3398 = REG1_REG_31_ & n1296;
  assign n3399 = REG0_REG_31_ & n1294;
  assign n3400 = REG2_REG_31_ & n1298;
  assign n3401 = ~n3398 & ~n3399;
  assign n3402 = ~n3400 & n3401;
  assign n3403 = n3338 & ~n3402;
  assign n3404 = n3316 & ~n3396;
  assign n3405 = ~n3316 & n3396;
  assign n3406 = ~n3404 & ~n3405;
  assign n3407 = n1305 & n3406;
  assign n3408 = ~n3397 & ~n3403;
  assign n3409 = ~n3407 & n3408;
  assign n3410 = n1268 & ~n3409;
  assign n3411 = REG0_REG_30_ & ~n1268;
  assign n644 = n3410 | n3411;
  assign n3413 = DATAI_31_ & ~n1275;
  assign n3414 = n1282_1 & n3413;
  assign n3415 = ~n3315 & ~n3396;
  assign n3416 = n3314 & n3415;
  assign n3417 = ~n3413 & n3416;
  assign n3418 = n3413 & ~n3416;
  assign n3419 = ~n3417 & ~n3418;
  assign n3420 = n1305 & n3419;
  assign n3421 = ~n3403 & ~n3414;
  assign n3422 = ~n3420 & n3421;
  assign n3423 = n1268 & ~n3422;
  assign n3424 = REG0_REG_31_ & ~n1268;
  assign n649 = n3423 | n3424;
  assign n3426 = n1134_1 & ~n1183;
  assign n3427 = n1267_1 & n3426;
  assign n3428 = ~n1349 & n3427;
  assign n3429 = REG1_REG_0_ & ~n3427;
  assign n654 = n3428 | n3429;
  assign n3431 = ~n1405 & n3427;
  assign n3432 = REG1_REG_1_ & ~n3427;
  assign n659 = n3431 | n3432;
  assign n3434 = ~n1467 & n3427;
  assign n3435 = REG1_REG_2_ & ~n3427;
  assign n664 = n3434 | n3435;
  assign n3437 = ~n1532 & n3427;
  assign n3438 = REG1_REG_3_ & ~n3427;
  assign n669 = n3437 | n3438;
  assign n3440 = ~n1603 & n3427;
  assign n3441 = REG1_REG_4_ & ~n3427;
  assign n674 = n3440 | n3441;
  assign n3443 = ~n1668 & n3427;
  assign n3444 = REG1_REG_5_ & ~n3427;
  assign n679 = n3443 | n3444;
  assign n3446 = ~n1749 & n3427;
  assign n3447 = REG1_REG_6_ & ~n3427;
  assign n684 = n3446 | n3447;
  assign n3449 = ~n1821 & n3427;
  assign n3450 = REG1_REG_7_ & ~n3427;
  assign n689 = n3449 | n3450;
  assign n3452 = ~n1889 & n3427;
  assign n3453 = REG1_REG_8_ & ~n3427;
  assign n694 = n3452 | n3453;
  assign n3455 = ~n1962 & n3427;
  assign n3456 = REG1_REG_9_ & ~n3427;
  assign n699 = n3455 | n3456;
  assign n3458 = ~n2026 & n3427;
  assign n3459 = REG1_REG_10_ & ~n3427;
  assign n704 = n3458 | n3459;
  assign n3461 = ~n2102 & n3427;
  assign n3462 = REG1_REG_11_ & ~n3427;
  assign n709 = n3461 | n3462;
  assign n3464 = ~n2169 & n3427;
  assign n3465 = REG1_REG_12_ & ~n3427;
  assign n714 = n3464 | n3465;
  assign n3467 = ~n2239 & n3427;
  assign n3468 = REG1_REG_13_ & ~n3427;
  assign n719 = n3467 | n3468;
  assign n3470 = ~n2306 & n3427;
  assign n3471 = REG1_REG_14_ & ~n3427;
  assign n724 = n3470 | n3471;
  assign n3473 = ~n2373 & n3427;
  assign n3474 = REG1_REG_15_ & ~n3427;
  assign n729 = n3473 | n3474;
  assign n3476 = ~n2443 & n3427;
  assign n3477 = REG1_REG_16_ & ~n3427;
  assign n734 = n3476 | n3477;
  assign n3479 = ~n2515 & n3427;
  assign n3480 = REG1_REG_17_ & ~n3427;
  assign n739 = n3479 | n3480;
  assign n3482 = ~n2584 & n3427;
  assign n3483 = REG1_REG_18_ & ~n3427;
  assign n744 = n3482 | n3483;
  assign n3485 = ~n2645 & n3427;
  assign n3486 = REG1_REG_19_ & ~n3427;
  assign n749 = n3485 | n3486;
  assign n3488 = ~n2704 & n3427;
  assign n3489 = REG1_REG_20_ & ~n3427;
  assign n754 = n3488 | n3489;
  assign n3491 = ~n2768 & n3427;
  assign n3492 = REG1_REG_21_ & ~n3427;
  assign n759 = n3491 | n3492;
  assign n3494 = ~n2841 & n3427;
  assign n3495 = REG1_REG_22_ & ~n3427;
  assign n764 = n3494 | n3495;
  assign n3497 = ~n2931 & n3427;
  assign n3498 = REG1_REG_23_ & ~n3427;
  assign n769 = n3497 | n3498;
  assign n3500 = ~n3003 & n3427;
  assign n3501 = REG1_REG_24_ & ~n3427;
  assign n774 = n3500 | n3501;
  assign n3503 = ~n3070 & n3427;
  assign n3504 = REG1_REG_25_ & ~n3427;
  assign n779 = n3503 | n3504;
  assign n3506 = ~n3146 & n3427;
  assign n3507 = REG1_REG_26_ & ~n3427;
  assign n784 = n3506 | n3507;
  assign n3509 = ~n3234 & n3427;
  assign n3510 = REG1_REG_27_ & ~n3427;
  assign n789 = n3509 | n3510;
  assign n3512 = ~n3309 & n3427;
  assign n3513 = REG1_REG_28_ & ~n3427;
  assign n794 = n3512 | n3513;
  assign n3515 = ~n3392 & n3427;
  assign n3516 = REG1_REG_29_ & ~n3427;
  assign n799 = n3515 | n3516;
  assign n3518 = ~n3409 & n3427;
  assign n3519 = REG1_REG_30_ & ~n3427;
  assign n804 = n3518 | n3519;
  assign n3521 = ~n3422 & n3427;
  assign n3522 = REG1_REG_31_ & ~n3427;
  assign n809 = n3521 | n3522;
  assign n3524 = n1193 & n1305;
  assign n3525 = n1197_1 & n1318;
  assign n3526 = ~n1194 & n1284;
  assign n3527 = n1183 & ~n3526;
  assign n3528 = ~n1187_1 & n3527;
  assign n3529 = n1266 & n3528;
  assign n3530 = ~n3525 & ~n3529;
  assign n3531 = n1134_1 & ~n3530;
  assign n3532 = n3524 & n3531;
  assign n3533 = ~n1281 & n3532;
  assign n3534 = n1282_1 & n3531;
  assign n3535 = ~n1281 & n3534;
  assign n3536 = ~n1348 & n3531;
  assign n3537 = REG2_REG_0_ & ~n3531;
  assign n3538 = ~n3536 & ~n3537;
  assign n3539 = ~n3533 & ~n3535;
  assign n3540 = n3538 & n3539;
  assign n3541 = n3525 & n3531;
  assign n3542 = REG3_REG_0_ & n3541;
  assign n3543 = n1285 & n3531;
  assign n3544 = ~n1302_1 & n3543;
  assign n3545 = n1190 & ~n1193;
  assign n3546 = ~n1197_1 & n3545;
  assign n3547 = n3531 & n3546;
  assign n3548 = ~n1316 & n3547;
  assign n3549 = ~n3542 & ~n3544;
  assign n3550 = ~n3548 & n3549;
  assign n814 = ~n3540 | ~n3550;
  assign n3552 = ~n1369 & n3532;
  assign n3553 = ~n1366 & n3534;
  assign n3554 = ~n1404 & n3531;
  assign n3555 = REG2_REG_1_ & ~n3531;
  assign n3556 = ~n3554 & ~n3555;
  assign n3557 = ~n3552 & ~n3553;
  assign n3558 = n3556 & n3557;
  assign n3559 = REG3_REG_1_ & n3541;
  assign n3560 = ~n1359 & n3543;
  assign n3561 = ~n1378 & n3547;
  assign n3562 = ~n3559 & ~n3560;
  assign n3563 = ~n3561 & n3562;
  assign n819 = ~n3558 | ~n3563;
  assign n3565 = n1426 & n3532;
  assign n3566 = ~n1422 & n3534;
  assign n3567 = ~n1466 & n3531;
  assign n3568 = REG2_REG_2_ & ~n3531;
  assign n3569 = ~n3567 & ~n3568;
  assign n3570 = ~n3565 & ~n3566;
  assign n3571 = n3569 & n3570;
  assign n3572 = REG3_REG_2_ & n3541;
  assign n3573 = ~n1415 & n3543;
  assign n3574 = n1440 & n3547;
  assign n3575 = ~n3572 & ~n3573;
  assign n3576 = ~n3574 & n3575;
  assign n824 = ~n3571 | ~n3576;
  assign n3578 = n1490 & n3532;
  assign n3579 = ~n1487 & n3534;
  assign n3580 = ~n1531 & n3531;
  assign n3581 = REG2_REG_3_ & ~n3531;
  assign n3582 = ~n3580 & ~n3581;
  assign n3583 = ~n3578 & ~n3579;
  assign n3584 = n3582 & n3583;
  assign n3585 = ~REG3_REG_3_ & n3541;
  assign n3586 = ~n1480 & n3543;
  assign n3587 = ~n1505 & n3547;
  assign n3588 = ~n3585 & ~n3586;
  assign n3589 = ~n3587 & n3588;
  assign n829 = ~n3584 | ~n3589;
  assign n3591 = n1557 & n3532;
  assign n3592 = ~n1553 & n3534;
  assign n3593 = ~n1602 & n3531;
  assign n3594 = REG2_REG_4_ & ~n3531;
  assign n3595 = ~n3593 & ~n3594;
  assign n3596 = ~n3591 & ~n3592;
  assign n3597 = n3595 & n3596;
  assign n3598 = ~n1473 & n3541;
  assign n3599 = ~n1546 & n3543;
  assign n3600 = ~n1573 & n3547;
  assign n3601 = ~n3598 & ~n3599;
  assign n3602 = ~n3600 & n3601;
  assign n834 = ~n3597 | ~n3602;
  assign n3604 = n1628 & n3532;
  assign n3605 = ~n1625 & n3534;
  assign n3606 = ~n3604 & ~n3605;
  assign n3607 = ~n1539 & n3541;
  assign n3608 = ~n1618 & n3543;
  assign n3609 = n1643 & n3547;
  assign n3610 = ~n3607 & ~n3608;
  assign n3611 = ~n3609 & n3610;
  assign n3612 = ~n1667 & n3531;
  assign n3613 = REG2_REG_5_ & ~n3531;
  assign n3614 = ~n3612 & ~n3613;
  assign n3615 = n3606 & n3611;
  assign n839 = ~n3614 | ~n3615;
  assign n3617 = n1695 & n3532;
  assign n3618 = ~n1691 & n3534;
  assign n3619 = ~n3617 & ~n3618;
  assign n3620 = ~n1611 & n3541;
  assign n3621 = ~n1684 & n3543;
  assign n3622 = ~n1721 & n3547;
  assign n3623 = ~n3620 & ~n3621;
  assign n3624 = ~n3622 & n3623;
  assign n3625 = ~n1748 & n3531;
  assign n3626 = REG2_REG_6_ & ~n3531;
  assign n3627 = ~n3625 & ~n3626;
  assign n3628 = n3619 & n3624;
  assign n844 = ~n3627 | ~n3628;
  assign n3630 = n1776 & n3532;
  assign n3631 = ~n1773 & n3534;
  assign n3632 = ~n3630 & ~n3631;
  assign n3633 = ~n1677 & n3541;
  assign n3634 = ~n1766 & n3543;
  assign n3635 = n1791 & n3547;
  assign n3636 = ~n3633 & ~n3634;
  assign n3637 = ~n3635 & n3636;
  assign n3638 = ~n1820 & n3531;
  assign n3639 = REG2_REG_7_ & ~n3531;
  assign n3640 = ~n3638 & ~n3639;
  assign n3641 = n3632 & n3637;
  assign n849 = ~n3640 | ~n3641;
  assign n3643 = n1845 & n3532;
  assign n3644 = ~n1842 & n3534;
  assign n3645 = ~n3643 & ~n3644;
  assign n3646 = ~n1759 & n3541;
  assign n3647 = ~n1835 & n3543;
  assign n3648 = ~n1862 & n3547;
  assign n3649 = ~n3646 & ~n3647;
  assign n3650 = ~n3648 & n3649;
  assign n3651 = ~n1888 & n3531;
  assign n3652 = REG2_REG_8_ & ~n3531;
  assign n3653 = ~n3651 & ~n3652;
  assign n3654 = n3645 & n3650;
  assign n854 = ~n3653 | ~n3654;
  assign n3656 = n1916 & n3532;
  assign n3657 = ~n1913 & n3534;
  assign n3658 = ~n3656 & ~n3657;
  assign n3659 = ~n1828 & n3541;
  assign n3660 = ~n1904 & n3543;
  assign n3661 = ~n1929 & n3547;
  assign n3662 = ~n3659 & ~n3660;
  assign n3663 = ~n3661 & n3662;
  assign n3664 = ~n1961 & n3531;
  assign n3665 = REG2_REG_9_ & ~n3531;
  assign n3666 = ~n3664 & ~n3665;
  assign n3667 = n3658 & n3663;
  assign n859 = ~n3666 | ~n3667;
  assign n3669 = n1986 & n3532;
  assign n3670 = ~n1983 & n3534;
  assign n3671 = ~n3669 & ~n3670;
  assign n3672 = ~n1897 & n3541;
  assign n3673 = ~n1976 & n3543;
  assign n3674 = n2001 & n3547;
  assign n3675 = ~n3672 & ~n3673;
  assign n3676 = ~n3674 & n3675;
  assign n3677 = ~n2025 & n3531;
  assign n3678 = REG2_REG_10_ & ~n3531;
  assign n3679 = ~n3677 & ~n3678;
  assign n3680 = n3671 & n3676;
  assign n864 = ~n3679 | ~n3680;
  assign n3682 = n2053 & n3532;
  assign n3683 = ~n2050 & n3534;
  assign n3684 = ~n3682 & ~n3683;
  assign n3685 = ~n1969 & n3541;
  assign n3686 = ~n2041 & n3543;
  assign n3687 = ~n2074 & n3547;
  assign n3688 = ~n3685 & ~n3686;
  assign n3689 = ~n3687 & n3688;
  assign n3690 = ~n2101 & n3531;
  assign n3691 = REG2_REG_11_ & ~n3531;
  assign n3692 = ~n3690 & ~n3691;
  assign n3693 = n3684 & n3689;
  assign n869 = ~n3692 | ~n3693;
  assign n3695 = n2126 & n3532;
  assign n3696 = ~n2123 & n3534;
  assign n3697 = ~n3695 & ~n3696;
  assign n3698 = ~n2034 & n3541;
  assign n3699 = ~n2116 & n3543;
  assign n3700 = ~n2139 & n3547;
  assign n3701 = ~n3698 & ~n3699;
  assign n3702 = ~n3700 & n3701;
  assign n3703 = ~n2168 & n3531;
  assign n3704 = REG2_REG_12_ & ~n3531;
  assign n3705 = ~n3703 & ~n3704;
  assign n3706 = n3697 & n3702;
  assign n874 = ~n3705 | ~n3706;
  assign n3708 = ~n2109 & n3541;
  assign n3709 = ~n2184 & n3543;
  assign n3710 = ~n3708 & ~n3709;
  assign n3711 = n2196 & n3532;
  assign n3712 = ~n2193 & n3534;
  assign n3713 = ~n3711 & ~n3712;
  assign n3714 = n2211 & n3547;
  assign n3715 = ~n2238 & n3531;
  assign n3716 = REG2_REG_13_ & ~n3531;
  assign n3717 = ~n3715 & ~n3716;
  assign n3718 = n3710 & n3713;
  assign n3719 = ~n3714 & n3718;
  assign n879 = ~n3717 | ~n3719;
  assign n3721 = n2263 & n3532;
  assign n3722 = ~n2260 & n3534;
  assign n3723 = ~n3721 & ~n3722;
  assign n3724 = ~n2177 & n3541;
  assign n3725 = ~n2253 & n3543;
  assign n3726 = ~n2278 & n3547;
  assign n3727 = ~n3724 & ~n3725;
  assign n3728 = ~n3726 & n3727;
  assign n3729 = ~n2305 & n3531;
  assign n3730 = REG2_REG_14_ & ~n3531;
  assign n3731 = ~n3729 & ~n3730;
  assign n3732 = n3723 & n3728;
  assign n884 = ~n3731 | ~n3732;
  assign n3734 = ~n2246 & n3541;
  assign n3735 = ~n2321 & n3543;
  assign n3736 = ~n3734 & ~n3735;
  assign n3737 = n2333 & n3532;
  assign n3738 = ~n2330 & n3534;
  assign n3739 = ~n3737 & ~n3738;
  assign n3740 = ~n2348 & n3547;
  assign n3741 = ~n2372 & n3531;
  assign n3742 = REG2_REG_15_ & ~n3531;
  assign n3743 = ~n3741 & ~n3742;
  assign n3744 = n3736 & n3739;
  assign n3745 = ~n3740 & n3744;
  assign n889 = ~n3743 | ~n3745;
  assign n3747 = ~n2314 & n3541;
  assign n3748 = ~n2387 & n3543;
  assign n3749 = ~n3747 & ~n3748;
  assign n3750 = n2397 & n3532;
  assign n3751 = ~n2394 & n3534;
  assign n3752 = ~n3750 & ~n3751;
  assign n3753 = ~n2415 & n3547;
  assign n3754 = ~n2442 & n3531;
  assign n3755 = REG2_REG_16_ & ~n3531;
  assign n3756 = ~n3754 & ~n3755;
  assign n3757 = n3749 & n3752;
  assign n3758 = ~n3753 & n3757;
  assign n894 = ~n3756 | ~n3758;
  assign n3760 = ~n2380 & n3541;
  assign n3761 = ~n2458 & n3543;
  assign n3762 = ~n3760 & ~n3761;
  assign n3763 = n2470 & n3532;
  assign n3764 = ~n2467 & n3534;
  assign n3765 = ~n3763 & ~n3764;
  assign n3766 = n2485 & n3547;
  assign n3767 = ~n2514 & n3531;
  assign n3768 = REG2_REG_17_ & ~n3531;
  assign n3769 = ~n3767 & ~n3768;
  assign n3770 = n3762 & n3765;
  assign n3771 = ~n3766 & n3770;
  assign n899 = ~n3769 | ~n3771;
  assign n3773 = ~n2451 & n3541;
  assign n3774 = ~n2529 & n3543;
  assign n3775 = ~n3773 & ~n3774;
  assign n3776 = n2539 & n3532;
  assign n3777 = ~n2536 & n3534;
  assign n3778 = ~n3776 & ~n3777;
  assign n3779 = ~n2556 & n3547;
  assign n3780 = ~n2583 & n3531;
  assign n3781 = REG2_REG_18_ & ~n3531;
  assign n3782 = ~n3780 & ~n3781;
  assign n3783 = n3775 & n3778;
  assign n3784 = ~n3779 & n3783;
  assign n904 = ~n3782 | ~n3784;
  assign n3786 = ~n2522 & n3541;
  assign n3787 = ~n2598 & n3543;
  assign n3788 = ~n3786 & ~n3787;
  assign n3789 = n2607 & n3532;
  assign n3790 = ~n2604 & n3534;
  assign n3791 = ~n3789 & ~n3790;
  assign n3792 = ~n2620 & n3547;
  assign n3793 = ~n2644 & n3531;
  assign n3794 = REG2_REG_19_ & ~n3531;
  assign n3795 = ~n3793 & ~n3794;
  assign n3796 = n3788 & n3791;
  assign n3797 = ~n3792 & n3796;
  assign n909 = ~n3795 | ~n3797;
  assign n3799 = ~n2591 & n3541;
  assign n3800 = ~n2659 & n3543;
  assign n3801 = ~n3799 & ~n3800;
  assign n3802 = n2664 & n3532;
  assign n3803 = n2661 & n3534;
  assign n3804 = ~n3802 & ~n3803;
  assign n3805 = n2679 & n3547;
  assign n3806 = ~n2703 & n3531;
  assign n3807 = REG2_REG_20_ & ~n3531;
  assign n3808 = ~n3806 & ~n3807;
  assign n3809 = n3801 & n3804;
  assign n3810 = ~n3805 & n3809;
  assign n914 = ~n3808 | ~n3810;
  assign n3812 = ~n2655 & n3541;
  assign n3813 = ~n2718 & n3543;
  assign n3814 = ~n3812 & ~n3813;
  assign n3815 = n2725 & n3532;
  assign n3816 = n2722 & n3534;
  assign n3817 = ~n3815 & ~n3816;
  assign n3818 = n2740 & n3547;
  assign n3819 = ~n2767 & n3531;
  assign n3820 = REG2_REG_21_ & ~n3531;
  assign n3821 = ~n3819 & ~n3820;
  assign n3822 = n3814 & n3817;
  assign n3823 = ~n3818 & n3822;
  assign n919 = ~n3821 | ~n3823;
  assign n3825 = ~n2714 & n3541;
  assign n3826 = ~n2782 & n3543;
  assign n3827 = ~n3825 & ~n3826;
  assign n3828 = n2787 & n3532;
  assign n3829 = n2784 & n3534;
  assign n3830 = ~n3828 & ~n3829;
  assign n3831 = ~n2808 & n3547;
  assign n3832 = ~n2840 & n3531;
  assign n3833 = REG2_REG_22_ & ~n3531;
  assign n3834 = ~n3832 & ~n3833;
  assign n3835 = n3827 & n3830;
  assign n3836 = ~n3831 & n3835;
  assign n924 = ~n3834 | ~n3836;
  assign n3838 = ~n2778 & n3541;
  assign n3839 = ~n2855 & n3543;
  assign n3840 = ~n3838 & ~n3839;
  assign n3841 = n2862 & n3532;
  assign n3842 = n2859 & n3534;
  assign n3843 = ~n3841 & ~n3842;
  assign n3844 = ~n2874 & n3547;
  assign n3845 = ~n2930 & n3531;
  assign n3846 = REG2_REG_23_ & ~n3531;
  assign n3847 = ~n3845 & ~n3846;
  assign n3848 = n3840 & n3843;
  assign n3849 = ~n3844 & n3848;
  assign n929 = ~n3847 | ~n3849;
  assign n3851 = ~n2851 & n3541;
  assign n3852 = ~n2945 & n3543;
  assign n3853 = ~n3851 & ~n3852;
  assign n3854 = n2950 & n3532;
  assign n3855 = n2947 & n3534;
  assign n3856 = ~n3854 & ~n3855;
  assign n3857 = ~n2965 & n3547;
  assign n3858 = ~n3002 & n3531;
  assign n3859 = REG2_REG_24_ & ~n3531;
  assign n3860 = ~n3858 & ~n3859;
  assign n3861 = n3853 & n3856;
  assign n3862 = ~n3857 & n3861;
  assign n934 = ~n3860 | ~n3862;
  assign n3864 = ~n2941 & n3541;
  assign n3865 = ~n3017 & n3543;
  assign n3866 = ~n3864 & ~n3865;
  assign n3867 = n3024 & n3532;
  assign n3868 = n3021 & n3534;
  assign n3869 = ~n3867 & ~n3868;
  assign n3870 = ~n3037 & n3547;
  assign n3871 = ~n3069 & n3531;
  assign n3872 = REG2_REG_25_ & ~n3531;
  assign n3873 = ~n3871 & ~n3872;
  assign n3874 = n3866 & n3869;
  assign n3875 = ~n3870 & n3874;
  assign n939 = ~n3873 | ~n3875;
  assign n3877 = ~n3013 & n3541;
  assign n3878 = ~n3084 & n3543;
  assign n3879 = ~n3877 & ~n3878;
  assign n3880 = n3089 & n3532;
  assign n3881 = n3086 & n3534;
  assign n3882 = ~n3880 & ~n3881;
  assign n3883 = n3104 & n3547;
  assign n3884 = ~n3145 & n3531;
  assign n3885 = REG2_REG_26_ & ~n3531;
  assign n3886 = ~n3884 & ~n3885;
  assign n3887 = n3879 & n3882;
  assign n3888 = ~n3883 & n3887;
  assign n944 = ~n3886 | ~n3888;
  assign n3890 = ~n3080 & n3541;
  assign n3891 = ~n3160 & n3543;
  assign n3892 = ~n3890 & ~n3891;
  assign n3893 = n3167 & n3532;
  assign n3894 = n3164 & n3534;
  assign n3895 = ~n3893 & ~n3894;
  assign n3896 = ~n3182 & n3547;
  assign n3897 = ~n3233 & n3531;
  assign n3898 = REG2_REG_27_ & ~n3531;
  assign n3899 = ~n3897 & ~n3898;
  assign n3900 = n3892 & n3895;
  assign n3901 = ~n3896 & n3900;
  assign n949 = ~n3899 | ~n3901;
  assign n3903 = ~n3156 & n3541;
  assign n3904 = ~n3246 & n3543;
  assign n3905 = ~n3903 & ~n3904;
  assign n3906 = n3251 & n3532;
  assign n3907 = n3248 & n3534;
  assign n3908 = ~n3906 & ~n3907;
  assign n3909 = ~n3263 & n3547;
  assign n3910 = ~n3308 & n3531;
  assign n3911 = REG2_REG_28_ & ~n3531;
  assign n3912 = ~n3910 & ~n3911;
  assign n3913 = n3905 & n3908;
  assign n3914 = ~n3909 & n3913;
  assign n954 = ~n3912 | ~n3914;
  assign n3916 = n3315 & n3534;
  assign n3917 = n3242 & n3541;
  assign n3918 = n3318 & n3532;
  assign n3919 = ~n3331 & n3547;
  assign n3920 = ~n3387 & n3388;
  assign n3921 = n3358 & ~n3384;
  assign n3922 = n3920 & n3921;
  assign n3923 = n3531 & ~n3922;
  assign n3924 = REG2_REG_29_ & ~n3531;
  assign n3925 = ~n3923 & ~n3924;
  assign n3926 = ~n3916 & ~n3917;
  assign n3927 = ~n3918 & n3926;
  assign n3928 = ~n3919 & n3927;
  assign n959 = ~n3925 | ~n3928;
  assign n3930 = n3406 & n3532;
  assign n3931 = n3396 & n3534;
  assign n3932 = n3403 & n3531;
  assign n3933 = REG2_REG_30_ & ~n3531;
  assign n3934 = ~n3932 & ~n3933;
  assign n3935 = ~n3930 & ~n3931;
  assign n964 = ~n3934 | ~n3935;
  assign n3937 = n3419 & n3532;
  assign n3938 = n3413 & n3534;
  assign n3939 = REG2_REG_31_ & ~n3531;
  assign n3940 = ~n3932 & ~n3939;
  assign n3941 = ~n3937 & ~n3938;
  assign n969 = ~n3940 | ~n3941;
  assign n3943 = STATE_REG & ~n1121;
  assign n3944 = n1121 & n1132;
  assign n3945 = n1133 & ~n1284;
  assign n3946 = n1121 & ~n3945;
  assign n3947 = ~n1275 & ~n3946;
  assign n1337 = ~STATE_REG | n3947;
  assign n3949 = ~n3944 & ~n1337;
  assign n3950 = n3943 & ~n3949;
  assign n3951 = n1274 & n3950;
  assign n3952 = ~n1193 & n3951;
  assign n3953 = ADDR_REG_19_ & n3949;
  assign n3954 = REG3_REG_19_ & ~STATE_REG;
  assign n3955 = ~n3953 & ~n3954;
  assign n3956 = n1271 & n3950;
  assign n3957 = ~REG1_REG_18_ & n2533;
  assign n3958 = REG1_REG_19_ & n1193;
  assign n3959 = ~REG1_REG_19_ & ~n1193;
  assign n3960 = ~n3958 & ~n3959;
  assign n3961 = ~n3957 & ~n3960;
  assign n3962 = REG1_REG_17_ & ~n2464;
  assign n3963 = ~REG1_REG_17_ & n2464;
  assign n3964 = REG1_REG_16_ & ~n2391;
  assign n3965 = ~REG1_REG_16_ & n2391;
  assign n3966 = REG1_REG_12_ & ~n2120;
  assign n3967 = ~REG1_REG_12_ & n2120;
  assign n3968 = REG1_REG_11_ & ~n2047;
  assign n3969 = ~REG1_REG_11_ & n2047;
  assign n3970 = REG1_REG_9_ & ~n1910;
  assign n3971 = ~REG1_REG_9_ & n1910;
  assign n3972 = REG1_REG_7_ & ~n1770;
  assign n3973 = ~REG1_REG_7_ & n1770;
  assign n3974 = REG1_REG_6_ & ~n1688;
  assign n3975 = ~REG1_REG_6_ & n1688;
  assign n3976 = REG1_REG_4_ & ~n1550;
  assign n3977 = ~REG1_REG_4_ & n1550;
  assign n3978 = REG1_REG_2_ & ~n1419;
  assign n3979 = ~REG1_REG_2_ & n1419;
  assign n3980 = REG1_REG_0_ & ~n1278;
  assign n3981 = REG1_REG_1_ & n3980;
  assign n3982 = ~REG1_REG_1_ & ~n3980;
  assign n3983 = ~n1363 & ~n3982;
  assign n3984 = ~n3981 & ~n3983;
  assign n3985 = ~n3979 & ~n3984;
  assign n3986 = ~n3978 & ~n3985;
  assign n3987 = REG1_REG_3_ & ~n3986;
  assign n3988 = ~REG1_REG_3_ & n3986;
  assign n3989 = ~n1484 & ~n3988;
  assign n3990 = ~n3987 & ~n3989;
  assign n3991 = ~n3977 & ~n3990;
  assign n3992 = ~n3976 & ~n3991;
  assign n3993 = REG1_REG_5_ & ~n3992;
  assign n3994 = ~REG1_REG_5_ & n3992;
  assign n3995 = ~n1622 & ~n3994;
  assign n3996 = ~n3993 & ~n3995;
  assign n3997 = ~n3975 & ~n3996;
  assign n3998 = ~n3974 & ~n3997;
  assign n3999 = ~n3973 & ~n3998;
  assign n4000 = ~n3972 & ~n3999;
  assign n4001 = REG1_REG_8_ & ~n4000;
  assign n4002 = ~REG1_REG_8_ & n4000;
  assign n4003 = ~n1839 & ~n4002;
  assign n4004 = ~n4001 & ~n4003;
  assign n4005 = ~n3971 & ~n4004;
  assign n4006 = ~n3970 & ~n4005;
  assign n4007 = REG1_REG_10_ & ~n4006;
  assign n4008 = ~REG1_REG_10_ & n4006;
  assign n4009 = ~n1980 & ~n4008;
  assign n4010 = ~n4007 & ~n4009;
  assign n4011 = ~n3969 & ~n4010;
  assign n4012 = ~n3968 & ~n4011;
  assign n4013 = ~n3967 & ~n4012;
  assign n4014 = ~n3966 & ~n4013;
  assign n4015 = REG1_REG_13_ & ~n4014;
  assign n4016 = ~REG1_REG_13_ & n4014;
  assign n4017 = ~n2190 & ~n4016;
  assign n4018 = ~n4015 & ~n4017;
  assign n4019 = REG1_REG_14_ & ~n4018;
  assign n4020 = ~REG1_REG_14_ & n4018;
  assign n4021 = ~n2257 & ~n4020;
  assign n4022 = ~n4019 & ~n4021;
  assign n4023 = REG1_REG_15_ & ~n4022;
  assign n4024 = ~REG1_REG_15_ & n4022;
  assign n4025 = ~n2327 & ~n4024;
  assign n4026 = ~n4023 & ~n4025;
  assign n4027 = ~n3965 & ~n4026;
  assign n4028 = ~n3964 & ~n4027;
  assign n4029 = ~n3963 & ~n4028;
  assign n4030 = ~n3962 & ~n4029;
  assign n4031 = REG1_REG_18_ & ~n2533;
  assign n4032 = n4030 & ~n4031;
  assign n4033 = n3961 & ~n4032;
  assign n4034 = n3960 & ~n4031;
  assign n4035 = ~n3957 & ~n4030;
  assign n4036 = n4034 & ~n4035;
  assign n4037 = ~n4033 & ~n4036;
  assign n4038 = n3956 & n4037;
  assign n4039 = ~n3952 & n3955;
  assign n4040 = ~n4038 & n4039;
  assign n4041 = ~n1282_1 & ~n3525;
  assign n4042 = ~n1336 & ~n1340;
  assign n4043 = ~n3524 & n4042;
  assign n4044 = ~n1324 & ~n1342;
  assign n4045 = ~n1333 & n4044;
  assign n4046 = ~n1330 & ~n3546;
  assign n4047 = ~n1328 & n4046;
  assign n4048 = n4041 & n4043;
  assign n4049 = n4045 & n4048;
  assign n4050 = n4047 & n4049;
  assign n4051 = n1274 & ~n4050;
  assign n4052 = ~n1193 & n4051;
  assign n4053 = n1134_1 & ~n3949;
  assign n4054 = n4052 & n4053;
  assign n4055 = ~n1271 & ~n1274;
  assign n4056 = ~n4050 & n4055;
  assign n4057 = ~REG2_REG_18_ & n2533;
  assign n4058 = REG2_REG_19_ & n1193;
  assign n4059 = ~REG2_REG_19_ & ~n1193;
  assign n4060 = ~n4058 & ~n4059;
  assign n4061 = ~n4057 & ~n4060;
  assign n4062 = REG2_REG_17_ & ~n2464;
  assign n4063 = ~REG2_REG_17_ & n2464;
  assign n4064 = REG2_REG_16_ & ~n2391;
  assign n4065 = ~REG2_REG_16_ & n2391;
  assign n4066 = REG2_REG_15_ & ~n2327;
  assign n4067 = ~REG2_REG_15_ & n2327;
  assign n4068 = REG2_REG_14_ & ~n2257;
  assign n4069 = ~REG2_REG_14_ & n2257;
  assign n4070 = REG2_REG_13_ & ~n2190;
  assign n4071 = ~REG2_REG_13_ & n2190;
  assign n4072 = REG2_REG_12_ & ~n2120;
  assign n4073 = ~REG2_REG_12_ & n2120;
  assign n4074 = REG2_REG_11_ & ~n2047;
  assign n4075 = ~REG2_REG_11_ & n2047;
  assign n4076 = REG2_REG_10_ & ~n1980;
  assign n4077 = ~REG2_REG_10_ & n1980;
  assign n4078 = REG2_REG_9_ & ~n1910;
  assign n4079 = ~REG2_REG_9_ & n1910;
  assign n4080 = REG2_REG_8_ & ~n1839;
  assign n4081 = ~REG2_REG_8_ & n1839;
  assign n4082 = REG2_REG_7_ & ~n1770;
  assign n4083 = ~REG2_REG_7_ & n1770;
  assign n4084 = REG2_REG_6_ & ~n1688;
  assign n4085 = ~REG2_REG_6_ & n1688;
  assign n4086 = REG2_REG_5_ & ~n1622;
  assign n4087 = ~REG2_REG_5_ & n1622;
  assign n4088 = REG2_REG_4_ & ~n1550;
  assign n4089 = ~REG2_REG_4_ & n1550;
  assign n4090 = REG2_REG_3_ & ~n1484;
  assign n4091 = ~REG2_REG_3_ & n1484;
  assign n4092 = REG2_REG_2_ & ~n1419;
  assign n4093 = ~REG2_REG_2_ & n1419;
  assign n4094 = REG2_REG_0_ & ~n1278;
  assign n4095 = ~n1363 & n4094;
  assign n4096 = n1363 & ~n4094;
  assign n4097 = REG2_REG_1_ & ~n4096;
  assign n4098 = ~n4095 & ~n4097;
  assign n4099 = ~n4093 & ~n4098;
  assign n4100 = ~n4092 & ~n4099;
  assign n4101 = ~n4091 & ~n4100;
  assign n4102 = ~n4090 & ~n4101;
  assign n4103 = ~n4089 & ~n4102;
  assign n4104 = ~n4088 & ~n4103;
  assign n4105 = ~n4087 & ~n4104;
  assign n4106 = ~n4086 & ~n4105;
  assign n4107 = ~n4085 & ~n4106;
  assign n4108 = ~n4084 & ~n4107;
  assign n4109 = ~n4083 & ~n4108;
  assign n4110 = ~n4082 & ~n4109;
  assign n4111 = ~n4081 & ~n4110;
  assign n4112 = ~n4080 & ~n4111;
  assign n4113 = ~n4079 & ~n4112;
  assign n4114 = ~n4078 & ~n4113;
  assign n4115 = ~n4077 & ~n4114;
  assign n4116 = ~n4076 & ~n4115;
  assign n4117 = ~n4075 & ~n4116;
  assign n4118 = ~n4074 & ~n4117;
  assign n4119 = ~n4073 & ~n4118;
  assign n4120 = ~n4072 & ~n4119;
  assign n4121 = ~n4071 & ~n4120;
  assign n4122 = ~n4070 & ~n4121;
  assign n4123 = ~n4069 & ~n4122;
  assign n4124 = ~n4068 & ~n4123;
  assign n4125 = ~n4067 & ~n4124;
  assign n4126 = ~n4066 & ~n4125;
  assign n4127 = ~n4065 & ~n4126;
  assign n4128 = ~n4064 & ~n4127;
  assign n4129 = ~n4063 & ~n4128;
  assign n4130 = ~n4062 & ~n4129;
  assign n4131 = REG2_REG_18_ & ~n2533;
  assign n4132 = n4130 & ~n4131;
  assign n4133 = n4061 & ~n4132;
  assign n4134 = n4060 & ~n4131;
  assign n4135 = ~n4057 & ~n4130;
  assign n4136 = n4134 & ~n4135;
  assign n4137 = ~n4133 & ~n4136;
  assign n4138 = n4053 & n4056;
  assign n4139 = n4137 & n4138;
  assign n4140 = n3950 & n4055;
  assign n4141 = n4137 & n4140;
  assign n4142 = n1271 & ~n4050;
  assign n4143 = n4053 & n4142;
  assign n4144 = n4037 & n4143;
  assign n4145 = ~n4054 & ~n4139;
  assign n4146 = ~n4141 & n4145;
  assign n4147 = ~n4144 & n4146;
  assign n974 = ~n4040 | ~n4147;
  assign n4149 = ~n2533 & n3951;
  assign n4150 = ADDR_REG_18_ & n3949;
  assign n4151 = REG3_REG_18_ & ~STATE_REG;
  assign n4152 = ~n4150 & ~n4151;
  assign n4153 = REG1_REG_18_ & n2533;
  assign n4154 = ~REG1_REG_18_ & ~n2533;
  assign n4155 = ~n4153 & ~n4154;
  assign n4156 = n4030 & ~n4155;
  assign n4157 = ~n4030 & n4155;
  assign n4158 = ~n4156 & ~n4157;
  assign n4159 = n3956 & ~n4158;
  assign n4160 = ~n4149 & n4152;
  assign n4161 = ~n4159 & n4160;
  assign n4162 = ~n2533 & n4051;
  assign n4163 = n4053 & n4162;
  assign n4164 = REG2_REG_18_ & n2533;
  assign n4165 = ~REG2_REG_18_ & ~n2533;
  assign n4166 = ~n4164 & ~n4165;
  assign n4167 = n4130 & ~n4166;
  assign n4168 = ~n4130 & n4166;
  assign n4169 = ~n4167 & ~n4168;
  assign n4170 = n4138 & ~n4169;
  assign n4171 = n4140 & ~n4169;
  assign n4172 = n4143 & ~n4158;
  assign n4173 = ~n4163 & ~n4170;
  assign n4174 = ~n4171 & n4173;
  assign n4175 = ~n4172 & n4174;
  assign n978 = ~n4161 | ~n4175;
  assign n4177 = ADDR_REG_17_ & n3949;
  assign n4178 = ~n2464 & n3951;
  assign n4179 = ~n4177 & ~n4178;
  assign n4180 = REG2_REG_17_ & n2464;
  assign n4181 = ~REG2_REG_17_ & ~n2464;
  assign n4182 = ~n4180 & ~n4181;
  assign n4183 = n4128 & ~n4182;
  assign n4184 = ~n4128 & n4182;
  assign n4185 = ~n4183 & ~n4184;
  assign n4186 = n4140 & ~n4185;
  assign n4187 = REG3_REG_17_ & ~STATE_REG;
  assign n4188 = ~n4186 & ~n4187;
  assign n4189 = REG1_REG_17_ & n2464;
  assign n4190 = ~REG1_REG_17_ & ~n2464;
  assign n4191 = ~n4189 & ~n4190;
  assign n4192 = n4028 & ~n4191;
  assign n4193 = ~n4028 & n4191;
  assign n4194 = ~n4192 & ~n4193;
  assign n4195 = n3956 & ~n4194;
  assign n4196 = ~n2464 & n4051;
  assign n4197 = n4056 & ~n4185;
  assign n4198 = n4142 & ~n4194;
  assign n4199 = ~n4196 & ~n4197;
  assign n4200 = ~n4198 & n4199;
  assign n4201 = n4053 & ~n4200;
  assign n4202 = n4179 & n4188;
  assign n4203 = ~n4195 & n4202;
  assign n982 = n4201 | ~n4203;
  assign n4205 = ADDR_REG_16_ & n3949;
  assign n4206 = ~n2391 & n3951;
  assign n4207 = ~n4205 & ~n4206;
  assign n4208 = REG2_REG_16_ & n2391;
  assign n4209 = ~REG2_REG_16_ & ~n2391;
  assign n4210 = ~n4208 & ~n4209;
  assign n4211 = n4126 & ~n4210;
  assign n4212 = ~n4126 & n4210;
  assign n4213 = ~n4211 & ~n4212;
  assign n4214 = n4140 & ~n4213;
  assign n4215 = REG3_REG_16_ & ~STATE_REG;
  assign n4216 = ~n4214 & ~n4215;
  assign n4217 = REG1_REG_16_ & n2391;
  assign n4218 = ~REG1_REG_16_ & ~n2391;
  assign n4219 = ~n4217 & ~n4218;
  assign n4220 = n4026 & ~n4219;
  assign n4221 = ~n4026 & n4219;
  assign n4222 = ~n4220 & ~n4221;
  assign n4223 = n3956 & ~n4222;
  assign n4224 = ~n2391 & n4051;
  assign n4225 = n4056 & ~n4213;
  assign n4226 = n4142 & ~n4222;
  assign n4227 = ~n4224 & ~n4225;
  assign n4228 = ~n4226 & n4227;
  assign n4229 = n4053 & ~n4228;
  assign n4230 = n4207 & n4216;
  assign n4231 = ~n4223 & n4230;
  assign n986 = n4229 | ~n4231;
  assign n4233 = ADDR_REG_15_ & n3949;
  assign n4234 = ~n2327 & n3951;
  assign n4235 = ~n4233 & ~n4234;
  assign n4236 = REG2_REG_15_ & n2327;
  assign n4237 = ~REG2_REG_15_ & ~n2327;
  assign n4238 = ~n4236 & ~n4237;
  assign n4239 = n4124 & ~n4238;
  assign n4240 = ~n4124 & n4238;
  assign n4241 = ~n4239 & ~n4240;
  assign n4242 = n4140 & ~n4241;
  assign n4243 = REG3_REG_15_ & ~STATE_REG;
  assign n4244 = ~n4242 & ~n4243;
  assign n4245 = ~n4023 & ~n4024;
  assign n4246 = ~n2327 & ~n4245;
  assign n4247 = n2327 & n4245;
  assign n4248 = ~n4246 & ~n4247;
  assign n4249 = n3956 & ~n4248;
  assign n4250 = ~n2327 & n4051;
  assign n4251 = n4056 & ~n4241;
  assign n4252 = n4142 & ~n4248;
  assign n4253 = ~n4250 & ~n4251;
  assign n4254 = ~n4252 & n4253;
  assign n4255 = n4053 & ~n4254;
  assign n4256 = n4235 & n4244;
  assign n4257 = ~n4249 & n4256;
  assign n990 = n4255 | ~n4257;
  assign n4259 = ADDR_REG_14_ & n3949;
  assign n4260 = ~n2257 & n3951;
  assign n4261 = ~n4259 & ~n4260;
  assign n4262 = REG2_REG_14_ & n2257;
  assign n4263 = ~REG2_REG_14_ & ~n2257;
  assign n4264 = ~n4262 & ~n4263;
  assign n4265 = n4122 & ~n4264;
  assign n4266 = ~n4122 & n4264;
  assign n4267 = ~n4265 & ~n4266;
  assign n4268 = n4140 & ~n4267;
  assign n4269 = REG3_REG_14_ & ~STATE_REG;
  assign n4270 = ~n4268 & ~n4269;
  assign n4271 = ~n4019 & ~n4020;
  assign n4272 = ~n2257 & ~n4271;
  assign n4273 = n2257 & n4271;
  assign n4274 = ~n4272 & ~n4273;
  assign n4275 = n3956 & ~n4274;
  assign n4276 = ~n2257 & n4051;
  assign n4277 = n4056 & ~n4267;
  assign n4278 = n4142 & ~n4274;
  assign n4279 = ~n4276 & ~n4277;
  assign n4280 = ~n4278 & n4279;
  assign n4281 = n4053 & ~n4280;
  assign n4282 = n4261 & n4270;
  assign n4283 = ~n4275 & n4282;
  assign n994 = n4281 | ~n4283;
  assign n4285 = ADDR_REG_13_ & n3949;
  assign n4286 = ~n2190 & n3951;
  assign n4287 = ~n4285 & ~n4286;
  assign n4288 = REG2_REG_13_ & n2190;
  assign n4289 = ~REG2_REG_13_ & ~n2190;
  assign n4290 = ~n4288 & ~n4289;
  assign n4291 = n4120 & ~n4290;
  assign n4292 = ~n4120 & n4290;
  assign n4293 = ~n4291 & ~n4292;
  assign n4294 = n4140 & ~n4293;
  assign n4295 = REG3_REG_13_ & ~STATE_REG;
  assign n4296 = ~n4294 & ~n4295;
  assign n4297 = ~n4015 & ~n4016;
  assign n4298 = ~n2190 & ~n4297;
  assign n4299 = n2190 & n4297;
  assign n4300 = ~n4298 & ~n4299;
  assign n4301 = n3956 & ~n4300;
  assign n4302 = ~n2190 & n4051;
  assign n4303 = n4056 & ~n4293;
  assign n4304 = n4142 & ~n4300;
  assign n4305 = ~n4302 & ~n4303;
  assign n4306 = ~n4304 & n4305;
  assign n4307 = n4053 & ~n4306;
  assign n4308 = n4287 & n4296;
  assign n4309 = ~n4301 & n4308;
  assign n998 = n4307 | ~n4309;
  assign n4311 = ADDR_REG_12_ & n3949;
  assign n4312 = ~n2120 & n3951;
  assign n4313 = ~n4311 & ~n4312;
  assign n4314 = REG2_REG_12_ & n2120;
  assign n4315 = ~REG2_REG_12_ & ~n2120;
  assign n4316 = ~n4314 & ~n4315;
  assign n4317 = n4118 & ~n4316;
  assign n4318 = ~n4118 & n4316;
  assign n4319 = ~n4317 & ~n4318;
  assign n4320 = n4140 & ~n4319;
  assign n4321 = REG3_REG_12_ & ~STATE_REG;
  assign n4322 = ~n4320 & ~n4321;
  assign n4323 = REG1_REG_12_ & n2120;
  assign n4324 = ~REG1_REG_12_ & ~n2120;
  assign n4325 = ~n4323 & ~n4324;
  assign n4326 = n4012 & ~n4325;
  assign n4327 = ~n4012 & n4325;
  assign n4328 = ~n4326 & ~n4327;
  assign n4329 = n3956 & ~n4328;
  assign n4330 = ~n2120 & n4051;
  assign n4331 = n4056 & ~n4319;
  assign n4332 = n4142 & ~n4328;
  assign n4333 = ~n4330 & ~n4331;
  assign n4334 = ~n4332 & n4333;
  assign n4335 = n4053 & ~n4334;
  assign n4336 = n4313 & n4322;
  assign n4337 = ~n4329 & n4336;
  assign n1002 = n4335 | ~n4337;
  assign n4339 = ADDR_REG_11_ & n3949;
  assign n4340 = ~n2047 & n3951;
  assign n4341 = ~n4339 & ~n4340;
  assign n4342 = REG2_REG_11_ & n2047;
  assign n4343 = ~REG2_REG_11_ & ~n2047;
  assign n4344 = ~n4342 & ~n4343;
  assign n4345 = n4116 & ~n4344;
  assign n4346 = ~n4116 & n4344;
  assign n4347 = ~n4345 & ~n4346;
  assign n4348 = n4140 & ~n4347;
  assign n4349 = REG3_REG_11_ & ~STATE_REG;
  assign n4350 = ~n4348 & ~n4349;
  assign n4351 = REG1_REG_11_ & n2047;
  assign n4352 = ~REG1_REG_11_ & ~n2047;
  assign n4353 = ~n4351 & ~n4352;
  assign n4354 = n4010 & ~n4353;
  assign n4355 = ~n4010 & n4353;
  assign n4356 = ~n4354 & ~n4355;
  assign n4357 = n3956 & ~n4356;
  assign n4358 = ~n2047 & n4051;
  assign n4359 = n4056 & ~n4347;
  assign n4360 = n4142 & ~n4356;
  assign n4361 = ~n4358 & ~n4359;
  assign n4362 = ~n4360 & n4361;
  assign n4363 = n4053 & ~n4362;
  assign n4364 = n4341 & n4350;
  assign n4365 = ~n4357 & n4364;
  assign n1006 = n4363 | ~n4365;
  assign n4367 = ADDR_REG_10_ & n3949;
  assign n4368 = ~n1980 & n3951;
  assign n4369 = ~n4367 & ~n4368;
  assign n4370 = REG2_REG_10_ & n1980;
  assign n4371 = ~REG2_REG_10_ & ~n1980;
  assign n4372 = ~n4370 & ~n4371;
  assign n4373 = n4114 & ~n4372;
  assign n4374 = ~n4114 & n4372;
  assign n4375 = ~n4373 & ~n4374;
  assign n4376 = n4140 & ~n4375;
  assign n4377 = REG3_REG_10_ & ~STATE_REG;
  assign n4378 = ~n4376 & ~n4377;
  assign n4379 = ~n4007 & ~n4008;
  assign n4380 = ~n1980 & ~n4379;
  assign n4381 = n1980 & n4379;
  assign n4382 = ~n4380 & ~n4381;
  assign n4383 = n3956 & ~n4382;
  assign n4384 = ~n1980 & n4051;
  assign n4385 = n4056 & ~n4375;
  assign n4386 = n4142 & ~n4382;
  assign n4387 = ~n4384 & ~n4385;
  assign n4388 = ~n4386 & n4387;
  assign n4389 = n4053 & ~n4388;
  assign n4390 = n4369 & n4378;
  assign n4391 = ~n4383 & n4390;
  assign n1010 = n4389 | ~n4391;
  assign n4393 = ADDR_REG_9_ & n3949;
  assign n4394 = ~n1910 & n3951;
  assign n4395 = ~n4393 & ~n4394;
  assign n4396 = REG2_REG_9_ & n1910;
  assign n4397 = ~REG2_REG_9_ & ~n1910;
  assign n4398 = ~n4396 & ~n4397;
  assign n4399 = n4112 & ~n4398;
  assign n4400 = ~n4112 & n4398;
  assign n4401 = ~n4399 & ~n4400;
  assign n4402 = n4140 & ~n4401;
  assign n4403 = REG3_REG_9_ & ~STATE_REG;
  assign n4404 = ~n4402 & ~n4403;
  assign n4405 = REG1_REG_9_ & n1910;
  assign n4406 = ~REG1_REG_9_ & ~n1910;
  assign n4407 = ~n4405 & ~n4406;
  assign n4408 = n4004 & ~n4407;
  assign n4409 = ~n4004 & n4407;
  assign n4410 = ~n4408 & ~n4409;
  assign n4411 = n3956 & ~n4410;
  assign n4412 = ~n1910 & n4051;
  assign n4413 = n4056 & ~n4401;
  assign n4414 = n4142 & ~n4410;
  assign n4415 = ~n4412 & ~n4413;
  assign n4416 = ~n4414 & n4415;
  assign n4417 = n4053 & ~n4416;
  assign n4418 = n4395 & n4404;
  assign n4419 = ~n4411 & n4418;
  assign n1014 = n4417 | ~n4419;
  assign n4421 = ADDR_REG_8_ & n3949;
  assign n4422 = ~n1839 & n3951;
  assign n4423 = ~n4421 & ~n4422;
  assign n4424 = REG2_REG_8_ & n1839;
  assign n4425 = ~REG2_REG_8_ & ~n1839;
  assign n4426 = ~n4424 & ~n4425;
  assign n4427 = n4110 & ~n4426;
  assign n4428 = ~n4110 & n4426;
  assign n4429 = ~n4427 & ~n4428;
  assign n4430 = n4140 & ~n4429;
  assign n4431 = REG3_REG_8_ & ~STATE_REG;
  assign n4432 = ~n4430 & ~n4431;
  assign n4433 = ~n4001 & ~n4002;
  assign n4434 = ~n1839 & ~n4433;
  assign n4435 = n1839 & n4433;
  assign n4436 = ~n4434 & ~n4435;
  assign n4437 = n3956 & ~n4436;
  assign n4438 = ~n1839 & n4051;
  assign n4439 = n4056 & ~n4429;
  assign n4440 = n4142 & ~n4436;
  assign n4441 = ~n4438 & ~n4439;
  assign n4442 = ~n4440 & n4441;
  assign n4443 = n4053 & ~n4442;
  assign n4444 = n4423 & n4432;
  assign n4445 = ~n4437 & n4444;
  assign n1018 = n4443 | ~n4445;
  assign n4447 = REG1_REG_7_ & n1770;
  assign n4448 = ~REG1_REG_7_ & ~n1770;
  assign n4449 = ~n4447 & ~n4448;
  assign n4450 = n3998 & ~n4449;
  assign n4451 = ~n3998 & n4449;
  assign n4452 = ~n4450 & ~n4451;
  assign n4453 = n3956 & ~n4452;
  assign n4454 = ~n1770 & n3951;
  assign n4455 = ADDR_REG_7_ & n3949;
  assign n4456 = ~n4453 & ~n4454;
  assign n4457 = ~n4455 & n4456;
  assign n4458 = REG2_REG_7_ & n1770;
  assign n4459 = ~REG2_REG_7_ & ~n1770;
  assign n4460 = ~n4458 & ~n4459;
  assign n4461 = n4108 & ~n4460;
  assign n4462 = ~n4108 & n4460;
  assign n4463 = ~n4461 & ~n4462;
  assign n4464 = n4140 & ~n4463;
  assign n4465 = REG3_REG_7_ & ~STATE_REG;
  assign n4466 = ~n1770 & n4051;
  assign n4467 = n4056 & ~n4463;
  assign n4468 = n4142 & ~n4452;
  assign n4469 = ~n4466 & ~n4467;
  assign n4470 = ~n4468 & n4469;
  assign n4471 = n4053 & ~n4470;
  assign n4472 = ~n4464 & ~n4465;
  assign n4473 = ~n4471 & n4472;
  assign n1022 = ~n4457 | ~n4473;
  assign n4475 = REG1_REG_6_ & n1688;
  assign n4476 = ~REG1_REG_6_ & ~n1688;
  assign n4477 = ~n4475 & ~n4476;
  assign n4478 = n3996 & ~n4477;
  assign n4479 = ~n3996 & n4477;
  assign n4480 = ~n4478 & ~n4479;
  assign n4481 = n3956 & ~n4480;
  assign n4482 = ~n1688 & n3951;
  assign n4483 = ADDR_REG_6_ & n3949;
  assign n4484 = ~n4481 & ~n4482;
  assign n4485 = ~n4483 & n4484;
  assign n4486 = REG2_REG_6_ & n1688;
  assign n4487 = ~REG2_REG_6_ & ~n1688;
  assign n4488 = ~n4486 & ~n4487;
  assign n4489 = n4106 & ~n4488;
  assign n4490 = ~n4106 & n4488;
  assign n4491 = ~n4489 & ~n4490;
  assign n4492 = n4140 & ~n4491;
  assign n4493 = REG3_REG_6_ & ~STATE_REG;
  assign n4494 = ~n1688 & n4051;
  assign n4495 = n4056 & ~n4491;
  assign n4496 = n4142 & ~n4480;
  assign n4497 = ~n4494 & ~n4495;
  assign n4498 = ~n4496 & n4497;
  assign n4499 = n4053 & ~n4498;
  assign n4500 = ~n4492 & ~n4493;
  assign n4501 = ~n4499 & n4500;
  assign n1026 = ~n4485 | ~n4501;
  assign n4503 = ~n3993 & ~n3994;
  assign n4504 = ~n1622 & ~n4503;
  assign n4505 = n1622 & n4503;
  assign n4506 = ~n4504 & ~n4505;
  assign n4507 = n3956 & ~n4506;
  assign n4508 = ~n1622 & n3951;
  assign n4509 = ADDR_REG_5_ & n3949;
  assign n4510 = ~n4507 & ~n4508;
  assign n4511 = ~n4509 & n4510;
  assign n4512 = REG2_REG_5_ & n1622;
  assign n4513 = ~REG2_REG_5_ & ~n1622;
  assign n4514 = ~n4512 & ~n4513;
  assign n4515 = n4104 & ~n4514;
  assign n4516 = ~n4104 & n4514;
  assign n4517 = ~n4515 & ~n4516;
  assign n4518 = n4140 & ~n4517;
  assign n4519 = REG3_REG_5_ & ~STATE_REG;
  assign n4520 = ~n1622 & n4051;
  assign n4521 = n4056 & ~n4517;
  assign n4522 = n4142 & ~n4506;
  assign n4523 = ~n4520 & ~n4521;
  assign n4524 = ~n4522 & n4523;
  assign n4525 = n4053 & ~n4524;
  assign n4526 = ~n4518 & ~n4519;
  assign n4527 = ~n4525 & n4526;
  assign n1030 = ~n4511 | ~n4527;
  assign n4529 = REG1_REG_4_ & n1550;
  assign n4530 = ~REG1_REG_4_ & ~n1550;
  assign n4531 = ~n4529 & ~n4530;
  assign n4532 = n3990 & ~n4531;
  assign n4533 = ~n3990 & n4531;
  assign n4534 = ~n4532 & ~n4533;
  assign n4535 = n3956 & ~n4534;
  assign n4536 = ~n1550 & n3951;
  assign n4537 = ADDR_REG_4_ & n3949;
  assign n4538 = ~n4535 & ~n4536;
  assign n4539 = ~n4537 & n4538;
  assign n4540 = REG3_REG_4_ & ~STATE_REG;
  assign n4541 = REG2_REG_4_ & n1550;
  assign n4542 = ~REG2_REG_4_ & ~n1550;
  assign n4543 = ~n4541 & ~n4542;
  assign n4544 = n4102 & ~n4543;
  assign n4545 = ~n4102 & n4543;
  assign n4546 = ~n4544 & ~n4545;
  assign n4547 = n4140 & ~n4546;
  assign n4548 = ~n1550 & n4051;
  assign n4549 = n4056 & ~n4546;
  assign n4550 = n4142 & ~n4534;
  assign n4551 = ~n4548 & ~n4549;
  assign n4552 = ~n4550 & n4551;
  assign n4553 = n4053 & ~n4552;
  assign n1341 = STATE_REG & n3944;
  assign n4555 = REG2_REG_0_ & n4055;
  assign n4556 = n1278 & n4555;
  assign n4557 = ~REG2_REG_0_ & ~n1271;
  assign n4558 = ~n1274 & ~n4557;
  assign n4559 = ~n1278 & ~n4558;
  assign n4560 = ~n1193 & n1197_1;
  assign n4561 = ~n1327_1 & ~n4560;
  assign n4562 = n1197_1 & n1201;
  assign n4563 = ~n1132 & n4562;
  assign n4564 = n4561 & ~n4563;
  assign n4565 = ~n1132 & ~n4564;
  assign n4566 = n1132 & ~n1278;
  assign n4567 = ~n1132 & ~n4046;
  assign n4568 = ~n1281 & n4567;
  assign n4569 = ~n4566 & ~n4568;
  assign n4570 = ~n1132 & n4560;
  assign n4571 = ~n1198 & ~n1324;
  assign n4572 = ~n1333 & n4571;
  assign n4573 = ~n1328 & n4572;
  assign n4574 = ~n1132 & ~n4573;
  assign n4575 = ~n4570 & ~n4574;
  assign n4576 = ~n1313 & ~n4575;
  assign n4577 = n4569 & ~n4576;
  assign n4578 = n4565 & n4577;
  assign n4579 = ~n4565 & ~n4577;
  assign n4580 = ~n4578 & ~n4579;
  assign n4581 = ~n1313 & n4567;
  assign n4582 = REG1_REG_0_ & n1132;
  assign n4583 = ~n4581 & ~n4582;
  assign n4584 = ~n4563 & ~n4570;
  assign n4585 = ~n4574 & n4584;
  assign n4586 = ~n1281 & ~n4585;
  assign n4587 = n4583 & ~n4586;
  assign n4588 = ~n4565 & ~n4587;
  assign n4589 = n4565 & n4587;
  assign n4590 = ~n4588 & ~n4589;
  assign n4591 = ~n4580 & n4590;
  assign n4592 = n4580 & ~n4590;
  assign n4593 = ~n4591 & ~n4592;
  assign n4594 = n1271 & ~n1274;
  assign n4595 = ~n4593 & n4594;
  assign n4596 = ~n4556 & ~n4559;
  assign n4597 = ~n4595 & n4596;
  assign n4598 = n1341 & ~n4597;
  assign n4599 = ~n4553 & ~n4598;
  assign n4600 = ~n4540 & ~n4547;
  assign n4601 = n4599 & n4600;
  assign n1034 = ~n4539 | ~n4601;
  assign n4603 = ~n3987 & ~n3988;
  assign n4604 = ~n1484 & ~n4603;
  assign n4605 = n1484 & n4603;
  assign n4606 = ~n4604 & ~n4605;
  assign n4607 = n3956 & ~n4606;
  assign n4608 = ~n1484 & n3951;
  assign n4609 = ADDR_REG_3_ & n3949;
  assign n4610 = ~n4607 & ~n4608;
  assign n4611 = ~n4609 & n4610;
  assign n4612 = REG2_REG_3_ & n1484;
  assign n4613 = ~REG2_REG_3_ & ~n1484;
  assign n4614 = ~n4612 & ~n4613;
  assign n4615 = n4100 & ~n4614;
  assign n4616 = ~n4100 & n4614;
  assign n4617 = ~n4615 & ~n4616;
  assign n4618 = n4140 & ~n4617;
  assign n4619 = REG3_REG_3_ & ~STATE_REG;
  assign n4620 = ~n1484 & n4051;
  assign n4621 = n4056 & ~n4617;
  assign n4622 = n4142 & ~n4606;
  assign n4623 = ~n4620 & ~n4621;
  assign n4624 = ~n4622 & n4623;
  assign n4625 = n4053 & ~n4624;
  assign n4626 = ~n4618 & ~n4619;
  assign n4627 = ~n4625 & n4626;
  assign n1038 = ~n4611 | ~n4627;
  assign n4629 = REG1_REG_2_ & n1419;
  assign n4630 = ~REG1_REG_2_ & ~n1419;
  assign n4631 = ~n4629 & ~n4630;
  assign n4632 = n3984 & ~n4631;
  assign n4633 = ~n3984 & n4631;
  assign n4634 = ~n4632 & ~n4633;
  assign n4635 = n3956 & ~n4634;
  assign n4636 = ~n1419 & n3951;
  assign n4637 = ADDR_REG_2_ & n3949;
  assign n4638 = ~n4635 & ~n4636;
  assign n4639 = ~n4637 & n4638;
  assign n4640 = REG3_REG_2_ & ~STATE_REG;
  assign n4641 = REG2_REG_2_ & n1419;
  assign n4642 = ~REG2_REG_2_ & ~n1419;
  assign n4643 = ~n4641 & ~n4642;
  assign n4644 = n4098 & ~n4643;
  assign n4645 = ~n4098 & n4643;
  assign n4646 = ~n4644 & ~n4645;
  assign n4647 = n4140 & ~n4646;
  assign n4648 = ~n1419 & n4051;
  assign n4649 = n4056 & ~n4646;
  assign n4650 = n4142 & ~n4634;
  assign n4651 = ~n4648 & ~n4649;
  assign n4652 = ~n4650 & n4651;
  assign n4653 = n4053 & ~n4652;
  assign n4654 = ~n4598 & ~n4653;
  assign n4655 = ~n4640 & ~n4647;
  assign n4656 = n4654 & n4655;
  assign n1042 = ~n4639 | ~n4656;
  assign n4658 = ~n1363 & n3981;
  assign n4659 = REG1_REG_1_ & ~n3980;
  assign n4660 = n1363 & n4659;
  assign n4661 = ~n4658 & ~n4660;
  assign n4662 = n1363 & n3980;
  assign n4663 = ~n1363 & ~n3980;
  assign n4664 = ~n4662 & ~n4663;
  assign n4665 = ~REG1_REG_1_ & ~n4664;
  assign n4666 = n4661 & ~n4665;
  assign n4667 = n3956 & ~n4666;
  assign n4668 = ~n1363 & n3951;
  assign n4669 = ADDR_REG_1_ & n3949;
  assign n4670 = ~n4667 & ~n4668;
  assign n4671 = ~n4669 & n4670;
  assign n4672 = REG2_REG_1_ & n4095;
  assign n4673 = ~n1363 & ~n4094;
  assign n4674 = ~REG2_REG_1_ & n4673;
  assign n4675 = ~n4672 & ~n4674;
  assign n4676 = ~REG2_REG_1_ & n4094;
  assign n4677 = REG2_REG_1_ & ~n4094;
  assign n4678 = ~n4676 & ~n4677;
  assign n4679 = n1363 & ~n4678;
  assign n4680 = n4675 & ~n4679;
  assign n4681 = n4140 & ~n4680;
  assign n4682 = REG3_REG_1_ & ~STATE_REG;
  assign n4683 = ~n1363 & n4051;
  assign n4684 = n4056 & ~n4680;
  assign n4685 = n4142 & ~n4666;
  assign n4686 = ~n4683 & ~n4684;
  assign n4687 = ~n4685 & n4686;
  assign n4688 = n4053 & ~n4687;
  assign n4689 = ~n4681 & ~n4682;
  assign n4690 = ~n4688 & n4689;
  assign n1046 = ~n4671 | ~n4690;
  assign n4692 = REG1_REG_0_ & n1278;
  assign n4693 = ~REG1_REG_0_ & ~n1278;
  assign n4694 = ~n4692 & ~n4693;
  assign n4695 = n3956 & ~n4694;
  assign n4696 = ~n1278 & n3951;
  assign n4697 = ADDR_REG_0_ & n3949;
  assign n4698 = ~n4695 & ~n4696;
  assign n4699 = ~n4697 & n4698;
  assign n4700 = REG2_REG_0_ & n1278;
  assign n4701 = ~REG2_REG_0_ & ~n1278;
  assign n4702 = ~n4700 & ~n4701;
  assign n4703 = n4140 & ~n4702;
  assign n4704 = REG3_REG_0_ & ~STATE_REG;
  assign n4705 = ~n1278 & n4051;
  assign n4706 = n4056 & ~n4702;
  assign n4707 = n4142 & ~n4694;
  assign n4708 = ~n4705 & ~n4706;
  assign n4709 = ~n4707 & n4708;
  assign n4710 = n4053 & ~n4709;
  assign n4711 = ~n4703 & ~n4704;
  assign n4712 = ~n4710 & n4711;
  assign n1050 = ~n4699 | ~n4712;
  assign n4714 = ~n1313 & n1341;
  assign n4715 = DATAO_REG_0_ & ~n1341;
  assign n1054 = n4714 | n4715;
  assign n4717 = ~n1302_1 & n1341;
  assign n4718 = DATAO_REG_1_ & ~n1341;
  assign n1058 = n4717 | n4718;
  assign n4720 = ~n1359 & n1341;
  assign n4721 = DATAO_REG_2_ & ~n1341;
  assign n1062 = n4720 | n4721;
  assign n4723 = ~n1415 & n1341;
  assign n4724 = DATAO_REG_3_ & ~n1341;
  assign n1066 = n4723 | n4724;
  assign n4726 = ~n1480 & n1341;
  assign n4727 = DATAO_REG_4_ & ~n1341;
  assign n1070 = n4726 | n4727;
  assign n4729 = ~n1546 & n1341;
  assign n4730 = DATAO_REG_5_ & ~n1341;
  assign n1074 = n4729 | n4730;
  assign n4732 = ~n1618 & n1341;
  assign n4733 = DATAO_REG_6_ & ~n1341;
  assign n1078 = n4732 | n4733;
  assign n4735 = ~n1684 & n1341;
  assign n4736 = DATAO_REG_7_ & ~n1341;
  assign n1082 = n4735 | n4736;
  assign n4738 = ~n1766 & n1341;
  assign n4739 = DATAO_REG_8_ & ~n1341;
  assign n1086 = n4738 | n4739;
  assign n4741 = ~n1835 & n1341;
  assign n4742 = DATAO_REG_9_ & ~n1341;
  assign n1090 = n4741 | n4742;
  assign n4744 = ~n1904 & n1341;
  assign n4745 = DATAO_REG_10_ & ~n1341;
  assign n1094 = n4744 | n4745;
  assign n4747 = ~n1976 & n1341;
  assign n4748 = DATAO_REG_11_ & ~n1341;
  assign n1098 = n4747 | n4748;
  assign n4750 = ~n2041 & n1341;
  assign n4751 = DATAO_REG_12_ & ~n1341;
  assign n1102 = n4750 | n4751;
  assign n4753 = ~n2116 & n1341;
  assign n4754 = DATAO_REG_13_ & ~n1341;
  assign n1106 = n4753 | n4754;
  assign n4756 = ~n2184 & n1341;
  assign n4757 = DATAO_REG_14_ & ~n1341;
  assign n1110 = n4756 | n4757;
  assign n4759 = ~n2253 & n1341;
  assign n4760 = DATAO_REG_15_ & ~n1341;
  assign n1114 = n4759 | n4760;
  assign n4762 = ~n2321 & n1341;
  assign n4763 = DATAO_REG_16_ & ~n1341;
  assign n1118 = n4762 | n4763;
  assign n4765 = ~n2387 & n1341;
  assign n4766 = DATAO_REG_17_ & ~n1341;
  assign n1122 = n4765 | n4766;
  assign n4768 = ~n2458 & n1341;
  assign n4769 = DATAO_REG_18_ & ~n1341;
  assign n1126 = n4768 | n4769;
  assign n4771 = ~n2529 & n1341;
  assign n4772 = DATAO_REG_19_ & ~n1341;
  assign n1130 = n4771 | n4772;
  assign n4774 = ~n2598 & n1341;
  assign n4775 = DATAO_REG_20_ & ~n1341;
  assign n1134 = n4774 | n4775;
  assign n4777 = ~n2659 & n1341;
  assign n4778 = DATAO_REG_21_ & ~n1341;
  assign n1138 = n4777 | n4778;
  assign n4780 = ~n2718 & n1341;
  assign n4781 = DATAO_REG_22_ & ~n1341;
  assign n1142 = n4780 | n4781;
  assign n4783 = ~n2782 & n1341;
  assign n4784 = DATAO_REG_23_ & ~n1341;
  assign n1146 = n4783 | n4784;
  assign n4786 = ~n2855 & n1341;
  assign n4787 = DATAO_REG_24_ & ~n1341;
  assign n1150 = n4786 | n4787;
  assign n4789 = ~n2945 & n1341;
  assign n4790 = DATAO_REG_25_ & ~n1341;
  assign n1154 = n4789 | n4790;
  assign n4792 = ~n3017 & n1341;
  assign n4793 = DATAO_REG_26_ & ~n1341;
  assign n1158 = n4792 | n4793;
  assign n4795 = ~n3084 & n1341;
  assign n4796 = DATAO_REG_27_ & ~n1341;
  assign n1162 = n4795 | n4796;
  assign n4798 = ~n3160 & n1341;
  assign n4799 = DATAO_REG_28_ & ~n1341;
  assign n1166 = n4798 | n4799;
  assign n4801 = ~n3246 & n1341;
  assign n4802 = DATAO_REG_29_ & ~n1341;
  assign n1170 = n4801 | n4802;
  assign n4804 = ~n3343 & n1341;
  assign n4805 = DATAO_REG_30_ & ~n1341;
  assign n1174 = n4804 | n4805;
  assign n4807 = ~n3402 & n1341;
  assign n4808 = DATAO_REG_31_ & ~n1341;
  assign n1178 = n4807 | n4808;
  assign n4810 = ~n1121 & ~n1201;
  assign n4811 = ~n1201 & n1330;
  assign n4812 = n4055 & n4811;
  assign n4813 = n1121 & ~n4812;
  assign n4814 = STATE_REG & ~n3944;
  assign n4815 = ~n4810 & ~n4813;
  assign n4816 = n4814 & n4815;
  assign n4817 = B_REG & ~n4816;
  assign n4818 = n1121 & n1323;
  assign n4819 = ~n1121 & n1323;
  assign n4820 = n3413 & n4819;
  assign n4821 = n1201 & ~n3402;
  assign n4822 = ~n4820 & ~n4821;
  assign n4823 = ~n3343 & n3402;
  assign n4824 = ~n3402 & ~n4823;
  assign n4825 = n3343 & ~n3402;
  assign n4826 = ~n4823 & ~n4825;
  assign n4827 = n4823 & n4826;
  assign n4828 = ~n4824 & ~n4827;
  assign n4829 = ~n1190 & ~n4828;
  assign n4830 = n4822 & ~n4829;
  assign n4831 = ~n3402 & n4819;
  assign n4832 = ~n1323 & n3413;
  assign n4833 = ~n4831 & ~n4832;
  assign n4834 = n4818 & n4830;
  assign n4835 = ~n4833 & n4834;
  assign n4836 = ~n4818 & ~n4830;
  assign n4837 = n4833 & n4836;
  assign n4838 = ~n4835 & ~n4837;
  assign n4839 = n4830 & ~n4833;
  assign n4840 = ~n4830 & n4833;
  assign n4841 = n3396 & n4819;
  assign n4842 = n1201 & ~n3343;
  assign n4843 = ~n4841 & ~n4842;
  assign n4844 = ~n3343 & ~n4823;
  assign n4845 = n3343 & n4823;
  assign n4846 = ~n4844 & ~n4845;
  assign n4847 = ~n1190 & ~n4846;
  assign n4848 = n4843 & ~n4847;
  assign n4849 = ~n3343 & n4819;
  assign n4850 = ~n1323 & n3396;
  assign n4851 = ~n4849 & ~n4850;
  assign n4852 = ~n4848 & n4851;
  assign n4853 = ~n4839 & ~n4840;
  assign n4854 = ~n4852 & n4853;
  assign n4855 = ~n3246 & n4819;
  assign n4856 = ~n1323 & n3315;
  assign n4857 = n1121 & ~n3160;
  assign n4858 = ~n4855 & ~n4856;
  assign n4859 = ~n4857 & n4858;
  assign n4860 = ~n3246 & ~n4823;
  assign n4861 = ~n3246 & n4823;
  assign n4862 = ~n4860 & ~n4861;
  assign n4863 = ~n1190 & ~n4862;
  assign n4864 = n1201 & ~n3246;
  assign n4865 = n3315 & n4819;
  assign n4866 = ~n1121 & ~n4865;
  assign n4867 = ~n4864 & n4866;
  assign n4868 = ~n4863 & n4867;
  assign n4869 = ~n4859 & n4868;
  assign n4870 = n4848 & ~n4851;
  assign n4871 = ~n4869 & ~n4870;
  assign n4872 = ~n3160 & ~n4823;
  assign n4873 = ~n3160 & n4823;
  assign n4874 = ~n4872 & ~n4873;
  assign n4875 = ~n1190 & ~n4874;
  assign n4876 = n1201 & ~n3160;
  assign n4877 = n3248 & n4819;
  assign n4878 = ~n1121 & ~n4877;
  assign n4879 = ~n4876 & n4878;
  assign n4880 = ~n4875 & n4879;
  assign n4881 = ~n3160 & n4819;
  assign n4882 = ~n1323 & n3248;
  assign n4883 = n1121 & ~n3084;
  assign n4884 = ~n4881 & ~n4882;
  assign n4885 = ~n4883 & n4884;
  assign n4886 = ~n4880 & n4885;
  assign n4887 = n4859 & ~n4868;
  assign n4888 = ~n4886 & ~n4887;
  assign n4889 = n1121 & ~n3017;
  assign n4890 = ~n1323 & n3164;
  assign n4891 = ~n3084 & n4819;
  assign n4892 = ~n4889 & ~n4890;
  assign n4893 = ~n4891 & n4892;
  assign n4894 = ~n3084 & ~n4823;
  assign n4895 = ~n3084 & n4823;
  assign n4896 = ~n4894 & ~n4895;
  assign n4897 = ~n1190 & ~n4896;
  assign n4898 = n1201 & ~n3084;
  assign n4899 = n3164 & n4819;
  assign n4900 = ~n1121 & ~n4899;
  assign n4901 = ~n4898 & n4900;
  assign n4902 = ~n4897 & n4901;
  assign n4903 = ~n4893 & n4902;
  assign n4904 = n4880 & ~n4885;
  assign n4905 = ~n4903 & ~n4904;
  assign n4906 = ~n3017 & ~n4823;
  assign n4907 = ~n3017 & n4823;
  assign n4908 = ~n4906 & ~n4907;
  assign n4909 = ~n1190 & ~n4908;
  assign n4910 = n1201 & ~n3017;
  assign n4911 = n3086 & n4819;
  assign n4912 = ~n1121 & ~n4911;
  assign n4913 = ~n4910 & n4912;
  assign n4914 = ~n4909 & n4913;
  assign n4915 = ~n3017 & n4819;
  assign n4916 = ~n1323 & n3086;
  assign n4917 = n1121 & ~n2945;
  assign n4918 = ~n4915 & ~n4916;
  assign n4919 = ~n4917 & n4918;
  assign n4920 = ~n4914 & n4919;
  assign n4921 = n4893 & ~n4902;
  assign n4922 = ~n4920 & ~n4921;
  assign n4923 = n1121 & ~n2855;
  assign n4924 = ~n1323 & n3021;
  assign n4925 = ~n2945 & n4819;
  assign n4926 = ~n4923 & ~n4924;
  assign n4927 = ~n4925 & n4926;
  assign n4928 = ~n2945 & ~n4823;
  assign n4929 = ~n2945 & n4823;
  assign n4930 = ~n4928 & ~n4929;
  assign n4931 = ~n1190 & ~n4930;
  assign n4932 = n1201 & ~n2945;
  assign n4933 = n3021 & n4819;
  assign n4934 = ~n1121 & ~n4933;
  assign n4935 = ~n4932 & n4934;
  assign n4936 = ~n4931 & n4935;
  assign n4937 = ~n4927 & n4936;
  assign n4938 = n4914 & ~n4919;
  assign n4939 = ~n4937 & ~n4938;
  assign n4940 = ~n2855 & ~n4823;
  assign n4941 = ~n2855 & n4823;
  assign n4942 = ~n4940 & ~n4941;
  assign n4943 = ~n1190 & ~n4942;
  assign n4944 = n1201 & ~n2855;
  assign n4945 = n2947 & n4819;
  assign n4946 = ~n1121 & ~n4945;
  assign n4947 = ~n4944 & n4946;
  assign n4948 = ~n4943 & n4947;
  assign n4949 = ~n2855 & n4819;
  assign n4950 = ~n1323 & n2947;
  assign n4951 = n1121 & ~n2782;
  assign n4952 = ~n4949 & ~n4950;
  assign n4953 = ~n4951 & n4952;
  assign n4954 = ~n4948 & n4953;
  assign n4955 = n4927 & ~n4936;
  assign n4956 = ~n4954 & ~n4955;
  assign n4957 = n1121 & ~n2718;
  assign n4958 = ~n1323 & n2859;
  assign n4959 = ~n2782 & n4819;
  assign n4960 = ~n4957 & ~n4958;
  assign n4961 = ~n4959 & n4960;
  assign n4962 = ~n2782 & ~n4823;
  assign n4963 = ~n2782 & n4823;
  assign n4964 = ~n4962 & ~n4963;
  assign n4965 = ~n1190 & ~n4964;
  assign n4966 = n1201 & ~n2782;
  assign n4967 = n2859 & n4819;
  assign n4968 = ~n1121 & ~n4967;
  assign n4969 = ~n4966 & n4968;
  assign n4970 = ~n4965 & n4969;
  assign n4971 = ~n4961 & n4970;
  assign n4972 = n4948 & ~n4953;
  assign n4973 = ~n4971 & ~n4972;
  assign n4974 = ~n2718 & ~n4823;
  assign n4975 = ~n2718 & n4823;
  assign n4976 = ~n4974 & ~n4975;
  assign n4977 = ~n1190 & ~n4976;
  assign n4978 = n1201 & ~n2718;
  assign n4979 = n2784 & n4819;
  assign n4980 = ~n1121 & ~n4979;
  assign n4981 = ~n4978 & n4980;
  assign n4982 = ~n4977 & n4981;
  assign n4983 = ~n2718 & n4819;
  assign n4984 = ~n1323 & n2784;
  assign n4985 = n1121 & ~n2659;
  assign n4986 = ~n4983 & ~n4984;
  assign n4987 = ~n4985 & n4986;
  assign n4988 = ~n4982 & n4987;
  assign n4989 = n4961 & ~n4970;
  assign n4990 = ~n4988 & ~n4989;
  assign n4991 = n1121 & ~n2598;
  assign n4992 = ~n1323 & n2722;
  assign n4993 = ~n2659 & n4819;
  assign n4994 = ~n4991 & ~n4992;
  assign n4995 = ~n4993 & n4994;
  assign n4996 = ~n2659 & ~n4823;
  assign n4997 = ~n2659 & n4823;
  assign n4998 = ~n4996 & ~n4997;
  assign n4999 = ~n1190 & ~n4998;
  assign n5000 = n1201 & ~n2659;
  assign n5001 = n2722 & n4819;
  assign n5002 = ~n1121 & ~n5001;
  assign n5003 = ~n5000 & n5002;
  assign n5004 = ~n4999 & n5003;
  assign n5005 = ~n4995 & n5004;
  assign n5006 = n4982 & ~n4987;
  assign n5007 = ~n5005 & ~n5006;
  assign n5008 = ~n2598 & ~n4823;
  assign n5009 = ~n2598 & n4823;
  assign n5010 = ~n5008 & ~n5009;
  assign n5011 = ~n1190 & ~n5010;
  assign n5012 = n1201 & ~n2598;
  assign n5013 = n2661 & n4819;
  assign n5014 = ~n1121 & ~n5013;
  assign n5015 = ~n5012 & n5014;
  assign n5016 = ~n5011 & n5015;
  assign n5017 = ~n2598 & n4819;
  assign n5018 = ~n1323 & n2661;
  assign n5019 = n1121 & ~n2529;
  assign n5020 = ~n5017 & ~n5018;
  assign n5021 = ~n5019 & n5020;
  assign n5022 = ~n5016 & n5021;
  assign n5023 = n4995 & ~n5004;
  assign n5024 = ~n5022 & ~n5023;
  assign n5025 = n1121 & ~n2458;
  assign n5026 = ~n1323 & ~n2604;
  assign n5027 = ~n2529 & n4819;
  assign n5028 = ~n5025 & ~n5026;
  assign n5029 = ~n5027 & n5028;
  assign n5030 = ~n2529 & ~n4823;
  assign n5031 = ~n2529 & n4823;
  assign n5032 = ~n5030 & ~n5031;
  assign n5033 = ~n1190 & ~n5032;
  assign n5034 = ~n2604 & n4819;
  assign n5035 = n1201 & ~n2529;
  assign n5036 = ~n1121 & ~n5034;
  assign n5037 = ~n5035 & n5036;
  assign n5038 = ~n5033 & n5037;
  assign n5039 = ~n5029 & n5038;
  assign n5040 = n5016 & ~n5021;
  assign n5041 = ~n5039 & ~n5040;
  assign n5042 = ~n2458 & ~n4823;
  assign n5043 = ~n2458 & n4823;
  assign n5044 = ~n5042 & ~n5043;
  assign n5045 = ~n1190 & ~n5044;
  assign n5046 = ~n2536 & n4819;
  assign n5047 = n1201 & ~n2458;
  assign n5048 = ~n1121 & ~n5046;
  assign n5049 = ~n5047 & n5048;
  assign n5050 = ~n5045 & n5049;
  assign n5051 = ~n2458 & n4819;
  assign n5052 = ~n1323 & ~n2536;
  assign n5053 = n1121 & ~n2387;
  assign n5054 = ~n5051 & ~n5052;
  assign n5055 = ~n5053 & n5054;
  assign n5056 = ~n5050 & n5055;
  assign n5057 = n5029 & ~n5038;
  assign n5058 = ~n5056 & ~n5057;
  assign n5059 = ~n2387 & n4819;
  assign n5060 = ~n1323 & ~n2467;
  assign n5061 = n1121 & ~n2321;
  assign n5062 = ~n5059 & ~n5060;
  assign n5063 = ~n5061 & n5062;
  assign n5064 = ~n2387 & ~n4823;
  assign n5065 = ~n2387 & n4823;
  assign n5066 = ~n5064 & ~n5065;
  assign n5067 = ~n1190 & ~n5066;
  assign n5068 = ~n2467 & n4819;
  assign n5069 = n1201 & ~n2387;
  assign n5070 = ~n1121 & ~n5068;
  assign n5071 = ~n5069 & n5070;
  assign n5072 = ~n5067 & n5071;
  assign n5073 = ~n5063 & n5072;
  assign n5074 = n5050 & ~n5055;
  assign n5075 = ~n5073 & ~n5074;
  assign n5076 = ~n2321 & ~n4823;
  assign n5077 = ~n2321 & n4823;
  assign n5078 = ~n5076 & ~n5077;
  assign n5079 = ~n1190 & ~n5078;
  assign n5080 = ~n2394 & n4819;
  assign n5081 = n1201 & ~n2321;
  assign n5082 = ~n1121 & ~n5080;
  assign n5083 = ~n5081 & n5082;
  assign n5084 = ~n5079 & n5083;
  assign n5085 = ~n2321 & n4819;
  assign n5086 = ~n1323 & ~n2394;
  assign n5087 = n1121 & ~n2253;
  assign n5088 = ~n5085 & ~n5086;
  assign n5089 = ~n5087 & n5088;
  assign n5090 = ~n5084 & n5089;
  assign n5091 = n5063 & ~n5072;
  assign n5092 = ~n5090 & ~n5091;
  assign n5093 = ~n2253 & n4819;
  assign n5094 = ~n1323 & ~n2330;
  assign n5095 = n1121 & ~n2184;
  assign n5096 = ~n5093 & ~n5094;
  assign n5097 = ~n5095 & n5096;
  assign n5098 = ~n2253 & ~n4823;
  assign n5099 = ~n2253 & n4823;
  assign n5100 = ~n5098 & ~n5099;
  assign n5101 = ~n1190 & ~n5100;
  assign n5102 = ~n2330 & n4819;
  assign n5103 = n1201 & ~n2253;
  assign n5104 = ~n1121 & ~n5102;
  assign n5105 = ~n5103 & n5104;
  assign n5106 = ~n5101 & n5105;
  assign n5107 = ~n5097 & n5106;
  assign n5108 = n5084 & ~n5089;
  assign n5109 = ~n5107 & ~n5108;
  assign n5110 = ~n2184 & ~n4823;
  assign n5111 = ~n2184 & n4823;
  assign n5112 = ~n5110 & ~n5111;
  assign n5113 = ~n1190 & ~n5112;
  assign n5114 = ~n2260 & n4819;
  assign n5115 = n1201 & ~n2184;
  assign n5116 = ~n1121 & ~n5114;
  assign n5117 = ~n5115 & n5116;
  assign n5118 = ~n5113 & n5117;
  assign n5119 = ~n2184 & n4819;
  assign n5120 = ~n1323 & ~n2260;
  assign n5121 = n1121 & ~n2116;
  assign n5122 = ~n5119 & ~n5120;
  assign n5123 = ~n5121 & n5122;
  assign n5124 = ~n5118 & n5123;
  assign n5125 = n5097 & ~n5106;
  assign n5126 = ~n5124 & ~n5125;
  assign n5127 = ~n1480 & n4819;
  assign n5128 = ~n1323 & ~n1553;
  assign n5129 = n1121 & ~n1415;
  assign n5130 = ~n5127 & ~n5128;
  assign n5131 = ~n5129 & n5130;
  assign n5132 = ~n1480 & ~n4823;
  assign n5133 = ~n1480 & n4823;
  assign n5134 = ~n5132 & ~n5133;
  assign n5135 = ~n1190 & ~n5134;
  assign n5136 = ~n1553 & n4819;
  assign n5137 = n1201 & ~n1480;
  assign n5138 = ~n1121 & ~n5136;
  assign n5139 = ~n5137 & n5138;
  assign n5140 = ~n5135 & n5139;
  assign n5141 = ~n5131 & n5140;
  assign n5142 = ~n1415 & n4819;
  assign n5143 = ~n1323 & ~n1487;
  assign n5144 = n1121 & ~n1359;
  assign n5145 = ~n5142 & ~n5143;
  assign n5146 = ~n5144 & n5145;
  assign n5147 = ~n1415 & ~n4823;
  assign n5148 = ~n1415 & n4823;
  assign n5149 = ~n5147 & ~n5148;
  assign n5150 = ~n1190 & ~n5149;
  assign n5151 = ~n1487 & n4819;
  assign n5152 = n1201 & ~n1415;
  assign n5153 = ~n1121 & ~n5151;
  assign n5154 = ~n5152 & n5153;
  assign n5155 = ~n5150 & n5154;
  assign n5156 = ~n5146 & n5155;
  assign n5157 = ~n1313 & n4819;
  assign n5158 = ~n1281 & ~n1323;
  assign n5159 = ~n5157 & ~n5158;
  assign n5160 = ~n1302_1 & n4819;
  assign n5161 = ~n1323 & ~n1366;
  assign n5162 = n1121 & ~n1313;
  assign n5163 = ~n5160 & ~n5161;
  assign n5164 = ~n5162 & n5163;
  assign n5165 = ~n1313 & ~n4823;
  assign n5166 = ~n1313 & n4823;
  assign n5167 = ~n5165 & ~n5166;
  assign n5168 = ~n1190 & ~n5167;
  assign n5169 = ~n1281 & n4819;
  assign n5170 = n1201 & ~n1313;
  assign n5171 = ~n1121 & ~n5169;
  assign n5172 = ~n5170 & n5171;
  assign n5173 = ~n5168 & n5172;
  assign n5174 = ~n5159 & ~n5164;
  assign n5175 = n5173 & n5174;
  assign n5176 = ~n5141 & ~n5156;
  assign n5177 = ~n5175 & n5176;
  assign n5178 = ~n1302_1 & ~n4823;
  assign n5179 = ~n1302_1 & n4823;
  assign n5180 = ~n5178 & ~n5179;
  assign n5181 = ~n1190 & ~n5180;
  assign n5182 = ~n1366 & n4819;
  assign n5183 = n1201 & ~n1302_1;
  assign n5184 = ~n1121 & ~n5182;
  assign n5185 = ~n5183 & n5184;
  assign n5186 = ~n5181 & n5185;
  assign n5187 = ~n5164 & n5186;
  assign n5188 = ~n1359 & n4819;
  assign n5189 = ~n1323 & ~n1422;
  assign n5190 = n1121 & ~n1302_1;
  assign n5191 = ~n5188 & ~n5189;
  assign n5192 = ~n5190 & n5191;
  assign n5193 = ~n1359 & ~n4823;
  assign n5194 = ~n1359 & n4823;
  assign n5195 = ~n5193 & ~n5194;
  assign n5196 = ~n1190 & ~n5195;
  assign n5197 = ~n1422 & n4819;
  assign n5198 = n1201 & ~n1359;
  assign n5199 = ~n1121 & ~n5197;
  assign n5200 = ~n5198 & n5199;
  assign n5201 = ~n5196 & n5200;
  assign n5202 = ~n5192 & n5201;
  assign n5203 = n5173 & n5186;
  assign n5204 = ~n5159 & n5203;
  assign n5205 = ~n5187 & ~n5202;
  assign n5206 = ~n5204 & n5205;
  assign n5207 = n5177 & n5206;
  assign n5208 = ~n1618 & ~n4823;
  assign n5209 = ~n1618 & n4823;
  assign n5210 = ~n5208 & ~n5209;
  assign n5211 = ~n1190 & ~n5210;
  assign n5212 = ~n1691 & n4819;
  assign n5213 = n1201 & ~n1618;
  assign n5214 = ~n1121 & ~n5212;
  assign n5215 = ~n5213 & n5214;
  assign n5216 = ~n5211 & n5215;
  assign n5217 = ~n1618 & n4819;
  assign n5218 = ~n1323 & ~n1691;
  assign n5219 = n1121 & ~n1546;
  assign n5220 = ~n5217 & ~n5218;
  assign n5221 = ~n5219 & n5220;
  assign n5222 = ~n5216 & n5221;
  assign n5223 = ~n1546 & ~n4823;
  assign n5224 = ~n1546 & n4823;
  assign n5225 = ~n5223 & ~n5224;
  assign n5226 = ~n1190 & ~n5225;
  assign n5227 = ~n1625 & n4819;
  assign n5228 = n1201 & ~n1546;
  assign n5229 = ~n1121 & ~n5227;
  assign n5230 = ~n5228 & n5229;
  assign n5231 = ~n5226 & n5230;
  assign n5232 = ~n1546 & n4819;
  assign n5233 = ~n1323 & ~n1625;
  assign n5234 = n1121 & ~n1480;
  assign n5235 = ~n5232 & ~n5233;
  assign n5236 = ~n5234 & n5235;
  assign n5237 = ~n5231 & n5236;
  assign n5238 = ~n1684 & ~n4823;
  assign n5239 = ~n1684 & n4823;
  assign n5240 = ~n5238 & ~n5239;
  assign n5241 = ~n1190 & ~n5240;
  assign n5242 = ~n1773 & n4819;
  assign n5243 = n1201 & ~n1684;
  assign n5244 = ~n1121 & ~n5242;
  assign n5245 = ~n5243 & n5244;
  assign n5246 = ~n5241 & n5245;
  assign n5247 = ~n1684 & n4819;
  assign n5248 = ~n1323 & ~n1773;
  assign n5249 = n1121 & ~n1618;
  assign n5250 = ~n5247 & ~n5248;
  assign n5251 = ~n5249 & n5250;
  assign n5252 = ~n5246 & n5251;
  assign n5253 = ~n5222 & ~n5237;
  assign n5254 = ~n5252 & n5253;
  assign n5255 = n5131 & ~n5140;
  assign n5256 = n5146 & ~n5155;
  assign n5257 = ~n5141 & n5256;
  assign n5258 = ~n5141 & ~n5201;
  assign n5259 = ~n5156 & n5258;
  assign n5260 = n5192 & n5259;
  assign n5261 = ~n5255 & ~n5257;
  assign n5262 = ~n5260 & n5261;
  assign n5263 = ~n5207 & n5254;
  assign n5264 = n5262 & n5263;
  assign n5265 = n5246 & ~n5251;
  assign n5266 = n5216 & ~n5221;
  assign n5267 = ~n5252 & n5266;
  assign n5268 = ~n5236 & ~n5252;
  assign n5269 = ~n5222 & n5268;
  assign n5270 = n5231 & n5269;
  assign n5271 = ~n1835 & n4819;
  assign n5272 = ~n1323 & ~n1913;
  assign n5273 = n1121 & ~n1766;
  assign n5274 = ~n5271 & ~n5272;
  assign n5275 = ~n5273 & n5274;
  assign n5276 = ~n1835 & ~n4823;
  assign n5277 = ~n1835 & n4823;
  assign n5278 = ~n5276 & ~n5277;
  assign n5279 = ~n1190 & ~n5278;
  assign n5280 = ~n1913 & n4819;
  assign n5281 = n1201 & ~n1835;
  assign n5282 = ~n1121 & ~n5280;
  assign n5283 = ~n5281 & n5282;
  assign n5284 = ~n5279 & n5283;
  assign n5285 = ~n5275 & n5284;
  assign n5286 = ~n1766 & n4819;
  assign n5287 = ~n1323 & ~n1842;
  assign n5288 = n1121 & ~n1684;
  assign n5289 = ~n5286 & ~n5287;
  assign n5290 = ~n5288 & n5289;
  assign n5291 = ~n1766 & ~n4823;
  assign n5292 = ~n1766 & n4823;
  assign n5293 = ~n5291 & ~n5292;
  assign n5294 = ~n1190 & ~n5293;
  assign n5295 = ~n1842 & n4819;
  assign n5296 = n1201 & ~n1766;
  assign n5297 = ~n1121 & ~n5295;
  assign n5298 = ~n5296 & n5297;
  assign n5299 = ~n5294 & n5298;
  assign n5300 = ~n5290 & n5299;
  assign n5301 = ~n1904 & n4819;
  assign n5302 = ~n1323 & ~n1983;
  assign n5303 = n1121 & ~n1835;
  assign n5304 = ~n5301 & ~n5302;
  assign n5305 = ~n5303 & n5304;
  assign n5306 = ~n1904 & ~n4823;
  assign n5307 = ~n1904 & n4823;
  assign n5308 = ~n5306 & ~n5307;
  assign n5309 = ~n1190 & ~n5308;
  assign n5310 = ~n1983 & n4819;
  assign n5311 = n1201 & ~n1904;
  assign n5312 = ~n1121 & ~n5310;
  assign n5313 = ~n5311 & n5312;
  assign n5314 = ~n5309 & n5313;
  assign n5315 = ~n5305 & n5314;
  assign n5316 = ~n5285 & ~n5300;
  assign n5317 = ~n5315 & n5316;
  assign n5318 = ~n5265 & ~n5267;
  assign n5319 = ~n5270 & n5318;
  assign n5320 = n5317 & n5319;
  assign n5321 = ~n5264 & n5320;
  assign n5322 = n5305 & ~n5314;
  assign n5323 = n5275 & ~n5284;
  assign n5324 = ~n5315 & n5323;
  assign n5325 = ~n5299 & ~n5315;
  assign n5326 = ~n5285 & n5325;
  assign n5327 = n5290 & n5326;
  assign n5328 = ~n2041 & ~n4823;
  assign n5329 = ~n2041 & n4823;
  assign n5330 = ~n5328 & ~n5329;
  assign n5331 = ~n1190 & ~n5330;
  assign n5332 = ~n2123 & n4819;
  assign n5333 = n1201 & ~n2041;
  assign n5334 = ~n1121 & ~n5332;
  assign n5335 = ~n5333 & n5334;
  assign n5336 = ~n5331 & n5335;
  assign n5337 = ~n2041 & n4819;
  assign n5338 = ~n1323 & ~n2123;
  assign n5339 = n1121 & ~n1976;
  assign n5340 = ~n5337 & ~n5338;
  assign n5341 = ~n5339 & n5340;
  assign n5342 = ~n5336 & n5341;
  assign n5343 = ~n1976 & ~n4823;
  assign n5344 = ~n1976 & n4823;
  assign n5345 = ~n5343 & ~n5344;
  assign n5346 = ~n1190 & ~n5345;
  assign n5347 = ~n2050 & n4819;
  assign n5348 = n1201 & ~n1976;
  assign n5349 = ~n1121 & ~n5347;
  assign n5350 = ~n5348 & n5349;
  assign n5351 = ~n5346 & n5350;
  assign n5352 = ~n1976 & n4819;
  assign n5353 = ~n1323 & ~n2050;
  assign n5354 = n1121 & ~n1904;
  assign n5355 = ~n5352 & ~n5353;
  assign n5356 = ~n5354 & n5355;
  assign n5357 = ~n5351 & n5356;
  assign n5358 = ~n2116 & ~n4823;
  assign n5359 = ~n2116 & n4823;
  assign n5360 = ~n5358 & ~n5359;
  assign n5361 = ~n1190 & ~n5360;
  assign n5362 = ~n2193 & n4819;
  assign n5363 = n1201 & ~n2116;
  assign n5364 = ~n1121 & ~n5362;
  assign n5365 = ~n5363 & n5364;
  assign n5366 = ~n5361 & n5365;
  assign n5367 = ~n2116 & n4819;
  assign n5368 = ~n1323 & ~n2193;
  assign n5369 = n1121 & ~n2041;
  assign n5370 = ~n5367 & ~n5368;
  assign n5371 = ~n5369 & n5370;
  assign n5372 = ~n5366 & n5371;
  assign n5373 = ~n5342 & ~n5357;
  assign n5374 = ~n5372 & n5373;
  assign n5375 = ~n5322 & ~n5324;
  assign n5376 = ~n5327 & n5375;
  assign n5377 = n5374 & n5376;
  assign n5378 = ~n5321 & n5377;
  assign n5379 = n5118 & ~n5123;
  assign n5380 = n5366 & ~n5371;
  assign n5381 = ~n5379 & ~n5380;
  assign n5382 = n5336 & ~n5341;
  assign n5383 = ~n5372 & n5382;
  assign n5384 = ~n5356 & ~n5372;
  assign n5385 = ~n5342 & n5384;
  assign n5386 = n5351 & n5385;
  assign n5387 = n5381 & ~n5383;
  assign n5388 = ~n5386 & n5387;
  assign n5389 = ~n5378 & n5388;
  assign n5390 = n5126 & ~n5389;
  assign n5391 = n5109 & ~n5390;
  assign n5392 = n5092 & ~n5391;
  assign n5393 = n5075 & ~n5392;
  assign n5394 = n5058 & ~n5393;
  assign n5395 = n5041 & ~n5394;
  assign n5396 = n5024 & ~n5395;
  assign n5397 = n5007 & ~n5396;
  assign n5398 = n4990 & ~n5397;
  assign n5399 = n4973 & ~n5398;
  assign n5400 = n4956 & ~n5399;
  assign n5401 = n4939 & ~n5400;
  assign n5402 = n4922 & ~n5401;
  assign n5403 = n4905 & ~n5402;
  assign n5404 = n4888 & ~n5403;
  assign n5405 = n4871 & ~n5404;
  assign n5406 = n4854 & ~n5405;
  assign n5407 = n4838 & ~n5406;
  assign n5408 = n1134_1 & n4812;
  assign n5409 = ~n5407 & n5408;
  assign n5410 = ~n4817 & ~n5409;
  assign n5411 = ~n1631 & ~n1632;
  assign n5412 = ~n2473 & ~n2475;
  assign n5413 = ~n1503 & ~n5411;
  assign n5414 = ~n1431 & n5413;
  assign n5415 = ~n5412 & n5414;
  assign n5416 = ~n1779 & ~n1781;
  assign n5417 = ~n1719 & ~n5416;
  assign n5418 = ~n2137 & n5417;
  assign n5419 = ~n2413 & n5418;
  assign n5420 = ~n2403 & ~n2405;
  assign n5421 = n1281 & n1313;
  assign n5422 = ~n1375 & ~n5421;
  assign n5423 = ~n2336 & ~n2338;
  assign n5424 = ~n5420 & ~n5422;
  assign n5425 = ~n1374 & n5424;
  assign n5426 = ~n5423 & n5425;
  assign n5427 = ~n2199 & ~n2200;
  assign n5428 = ~n2554 & ~n5427;
  assign n5429 = ~n1927 & n5428;
  assign n5430 = ~n1860 & n5429;
  assign n5431 = n3160 & ~n3248;
  assign n5432 = ~n3323 & ~n5431;
  assign n5433 = ~n3254 & ~n3255;
  assign n5434 = ~n5432 & ~n5433;
  assign n5435 = n5415 & n5419;
  assign n5436 = n5426 & n5435;
  assign n5437 = n5430 & n5436;
  assign n5438 = n5434 & n5437;
  assign n5439 = ~n1989 & ~n1990;
  assign n5440 = ~n1571 & ~n2618;
  assign n5441 = ~n5439 & n5440;
  assign n5442 = ~n2072 & n5441;
  assign n5443 = n3343 & ~n3396;
  assign n5444 = ~n3343 & n3396;
  assign n5445 = ~n5443 & ~n5444;
  assign n5446 = n3402 & ~n3413;
  assign n5447 = ~n3402 & n3413;
  assign n5448 = ~n5446 & ~n5447;
  assign n5449 = ~n2667 & ~n2668;
  assign n5450 = ~n5445 & ~n5448;
  assign n5451 = ~n5449 & n5450;
  assign n5452 = n3246 & ~n3315;
  assign n5453 = ~n3246 & n3315;
  assign n5454 = ~n5452 & ~n5453;
  assign n5455 = ~n2953 & ~n2954;
  assign n5456 = ~n2865 & ~n2866;
  assign n5457 = ~n2790 & ~n2795;
  assign n5458 = ~n2963 & ~n5455;
  assign n5459 = ~n5456 & n5458;
  assign n5460 = ~n5457 & n5459;
  assign n5461 = ~n3092 & ~n3093;
  assign n5462 = ~n3035 & ~n5461;
  assign n5463 = n5442 & n5451;
  assign n5464 = ~n5454 & n5463;
  assign n5465 = n5460 & n5464;
  assign n5466 = n5462 & n5465;
  assign n5467 = n5438 & n5466;
  assign n5468 = n1198 & ~n5467;
  assign n5469 = ~n1193 & n5468;
  assign n5470 = n1284 & ~n5407;
  assign n5471 = ~n1190 & n5470;
  assign n5472 = n2870 & ~n2957;
  assign n5473 = ~n2958 & ~n5472;
  assign n5474 = ~n3028 & n5473;
  assign n5475 = ~n3099 & n5474;
  assign n5476 = ~n2130 & ~n2206;
  assign n5477 = ~n2274 & ~n2344;
  assign n5478 = ~n2549 & ~n2611;
  assign n5479 = ~n2674 & ~n2729;
  assign n5480 = n2480 & ~n2548;
  assign n5481 = ~n2401 & n5478;
  assign n5482 = n5479 & n5481;
  assign n5483 = ~n5480 & n5482;
  assign n5484 = n5477 & n5483;
  assign n5485 = n5476 & n5484;
  assign n5486 = ~n1855 & ~n1920;
  assign n5487 = n2067 & ~n2129;
  assign n5488 = ~n1786 & n5486;
  assign n5489 = ~n1996 & n5488;
  assign n5490 = ~n5487 & n5489;
  assign n5491 = ~n1699 & n5490;
  assign n5492 = ~n2869 & ~n2957;
  assign n5493 = n2804 & n5492;
  assign n5494 = n1638 & ~n1698;
  assign n5495 = ~n5493 & ~n5494;
  assign n5496 = n5485 & n5491;
  assign n5497 = n5495 & n5496;
  assign n5498 = n5475 & n5497;
  assign n5499 = ~n3343 & ~n3396;
  assign n5500 = n3402 & n3413;
  assign n5501 = ~n5499 & ~n5500;
  assign n5502 = ~n3327 & n5501;
  assign n5503 = ~n3178 & n5502;
  assign n5504 = n1480 & n5503;
  assign n5505 = ~n1553 & n5498;
  assign n5506 = ~n3259 & n5505;
  assign n5507 = n5504 & n5506;
  assign n5508 = ~n5487 & ~n5493;
  assign n5509 = ~n3099 & n5508;
  assign n5510 = ~n1996 & n5485;
  assign n5511 = n5474 & n5510;
  assign n5512 = n5509 & n5511;
  assign n5513 = n1766 & ~n1920;
  assign n5514 = ~n3259 & n5513;
  assign n5515 = ~n1842 & n5512;
  assign n5516 = n5503 & n5515;
  assign n5517 = n5514 & n5516;
  assign n5518 = ~n1498 & ~n1561;
  assign n5519 = n1359 & n5518;
  assign n5520 = ~n3259 & n5519;
  assign n5521 = ~n1422 & n5497;
  assign n5522 = n5475 & n5521;
  assign n5523 = n5503 & n5522;
  assign n5524 = n5520 & n5523;
  assign n5525 = ~n5507 & ~n5517;
  assign n5526 = ~n5524 & n5525;
  assign n5527 = n1904 & ~n3259;
  assign n5528 = n5485 & ~n5493;
  assign n5529 = ~n1983 & n5528;
  assign n5530 = n5475 & n5529;
  assign n5531 = ~n5487 & n5530;
  assign n5532 = n5503 & n5531;
  assign n5533 = n5527 & n5532;
  assign n5534 = ~n2260 & n5483;
  assign n5535 = n5475 & ~n5493;
  assign n5536 = ~n2344 & n5503;
  assign n5537 = n2184 & ~n3259;
  assign n5538 = n5534 & n5535;
  assign n5539 = n5536 & n5538;
  assign n5540 = n5537 & n5539;
  assign n5541 = ~n2394 & n5478;
  assign n5542 = ~n2674 & ~n5493;
  assign n5543 = ~n3099 & n5542;
  assign n5544 = n5474 & n5543;
  assign n5545 = ~n2729 & n5544;
  assign n5546 = ~n5480 & n5503;
  assign n5547 = n2321 & ~n3259;
  assign n5548 = n5541 & n5545;
  assign n5549 = n5546 & n5548;
  assign n5550 = n5547 & n5549;
  assign n5551 = n2598 & ~n2729;
  assign n5552 = ~n3259 & n5551;
  assign n5553 = n2661 & n5535;
  assign n5554 = n5503 & n5553;
  assign n5555 = n5552 & n5554;
  assign n5556 = ~n5550 & ~n5555;
  assign n5557 = ~n5533 & ~n5540;
  assign n5558 = n5556 & n5557;
  assign n5559 = n2458 & ~n2611;
  assign n5560 = ~n3259 & n5559;
  assign n5561 = ~n2536 & n5545;
  assign n5562 = n5503 & n5561;
  assign n5563 = n5560 & n5562;
  assign n5564 = ~n2728 & ~n2803;
  assign n5565 = n5492 & n5564;
  assign n5566 = ~n3259 & ~n5565;
  assign n5567 = n5503 & n5535;
  assign n5568 = n5566 & n5567;
  assign n5569 = ~n2467 & n5478;
  assign n5570 = n2387 & n5503;
  assign n5571 = n5545 & n5569;
  assign n5572 = ~n3259 & n5571;
  assign n5573 = n5570 & n5572;
  assign n5574 = n3248 & ~n5499;
  assign n5575 = ~n3327 & n5574;
  assign n5576 = n3160 & n5575;
  assign n5577 = ~n5500 & n5576;
  assign n5578 = n3343 & n3396;
  assign n5579 = n3315 & ~n5499;
  assign n5580 = n3246 & n5579;
  assign n5581 = ~n5578 & ~n5580;
  assign n5582 = ~n5500 & ~n5581;
  assign n5583 = n3164 & ~n3327;
  assign n5584 = ~n5499 & n5583;
  assign n5585 = n3084 & n5584;
  assign n5586 = ~n5500 & n5585;
  assign n5587 = ~n3259 & n5586;
  assign n5588 = ~n5577 & ~n5582;
  assign n5589 = ~n5587 & n5588;
  assign n5590 = ~n5563 & ~n5568;
  assign n5591 = ~n5573 & n5590;
  assign n5592 = n5589 & n5591;
  assign n5593 = n1415 & ~n1561;
  assign n5594 = ~n3259 & n5593;
  assign n5595 = ~n1487 & n5498;
  assign n5596 = n5503 & n5595;
  assign n5597 = n5594 & n5596;
  assign n5598 = n1546 & ~n3259;
  assign n5599 = ~n1625 & n5528;
  assign n5600 = n5475 & n5599;
  assign n5601 = n5491 & n5600;
  assign n5602 = n5503 & n5601;
  assign n5603 = n5598 & n5602;
  assign n5604 = ~n1691 & n5503;
  assign n5605 = n1618 & ~n3259;
  assign n5606 = n5485 & n5490;
  assign n5607 = n5535 & n5606;
  assign n5608 = n5604 & n5607;
  assign n5609 = n5605 & n5608;
  assign n5610 = ~n2330 & n5483;
  assign n5611 = n2253 & n5503;
  assign n5612 = n5535 & n5610;
  assign n5613 = ~n3259 & n5612;
  assign n5614 = n5611 & n5613;
  assign n5615 = ~n5609 & ~n5614;
  assign n5616 = n2116 & n5503;
  assign n5617 = ~n2193 & n5484;
  assign n5618 = n5535 & n5617;
  assign n5619 = ~n3259 & n5618;
  assign n5620 = n5616 & n5619;
  assign n5621 = n2529 & n5503;
  assign n5622 = ~n2604 & n5545;
  assign n5623 = ~n3259 & n5622;
  assign n5624 = n5621 & n5623;
  assign n5625 = ~n5620 & ~n5624;
  assign n5626 = ~n1773 & n5486;
  assign n5627 = n1684 & n5503;
  assign n5628 = n5512 & n5626;
  assign n5629 = ~n3259 & n5628;
  assign n5630 = n5627 & n5629;
  assign n5631 = ~n5597 & ~n5603;
  assign n5632 = n5615 & n5631;
  assign n5633 = n5625 & n5632;
  assign n5634 = ~n5630 & n5633;
  assign n5635 = ~n1436 & n5518;
  assign n5636 = ~n1366 & n5635;
  assign n5637 = n1302_1 & n5503;
  assign n5638 = n5498 & n5636;
  assign n5639 = ~n3259 & n5638;
  assign n5640 = n5637 & n5639;
  assign n5641 = n3027 & ~n3099;
  assign n5642 = ~n3098 & ~n5641;
  assign n5643 = n5503 & ~n5642;
  assign n5644 = ~n3259 & n5643;
  assign n5645 = ~n3402 & ~n3413;
  assign n5646 = ~n2804 & ~n3259;
  assign n5647 = n1197_1 & ~n1317_1;
  assign n5648 = n1281 & n5647;
  assign n5649 = ~n1281 & ~n5647;
  assign n5650 = ~n1313 & ~n5649;
  assign n5651 = ~n1383 & ~n5650;
  assign n5652 = n5635 & ~n5648;
  assign n5653 = n5651 & n5652;
  assign n5654 = ~n5494 & n5653;
  assign n5655 = n5485 & n5654;
  assign n5656 = n5475 & n5655;
  assign n5657 = n5491 & n5656;
  assign n5658 = n5503 & n5657;
  assign n5659 = n5646 & n5658;
  assign n5660 = ~n5645 & ~n5659;
  assign n5661 = n1976 & n5503;
  assign n5662 = ~n2050 & n5528;
  assign n5663 = n5475 & n5662;
  assign n5664 = ~n3259 & n5663;
  assign n5665 = n5661 & n5664;
  assign n5666 = n1835 & n5503;
  assign n5667 = ~n1913 & n5512;
  assign n5668 = ~n3259 & n5667;
  assign n5669 = n5666 & n5668;
  assign n5670 = ~n2206 & n5503;
  assign n5671 = n2041 & ~n3259;
  assign n5672 = ~n2123 & n5484;
  assign n5673 = n5535 & n5672;
  assign n5674 = n5670 & n5673;
  assign n5675 = n5671 & n5674;
  assign n5676 = ~n5665 & ~n5669;
  assign n5677 = ~n5675 & n5676;
  assign n5678 = ~n5640 & ~n5644;
  assign n5679 = n5660 & n5678;
  assign n5680 = n5677 & n5679;
  assign n5681 = n5526 & n5558;
  assign n5682 = n5592 & n5681;
  assign n5683 = n5634 & n5682;
  assign n5684 = n5680 & n5683;
  assign n5685 = ~n1284 & ~n5684;
  assign n5686 = n1284 & n5407;
  assign n5687 = ~n5685 & ~n5686;
  assign n5688 = n1190 & ~n5687;
  assign n5689 = ~n5471 & ~n5688;
  assign n5690 = n1198 & n5467;
  assign n5691 = n5689 & ~n5690;
  assign n5692 = n1193 & ~n5691;
  assign n5693 = n1201 & n1328;
  assign n5694 = n3021 & n4930;
  assign n5695 = n2859 & n4964;
  assign n5696 = ~n2947 & ~n4942;
  assign n5697 = n5695 & ~n5696;
  assign n5698 = n2947 & n4942;
  assign n5699 = ~n5697 & ~n5698;
  assign n5700 = ~n1842 & n5293;
  assign n5701 = ~n1773 & n5240;
  assign n5702 = ~n1913 & n5278;
  assign n5703 = ~n1983 & n5308;
  assign n5704 = ~n5700 & ~n5701;
  assign n5705 = ~n5702 & n5704;
  assign n5706 = ~n5703 & n5705;
  assign n5707 = n1691 & ~n5210;
  assign n5708 = n1773 & ~n5240;
  assign n5709 = ~n5707 & ~n5708;
  assign n5710 = ~n1625 & n5225;
  assign n5711 = ~n1691 & n5210;
  assign n5712 = ~n5710 & ~n5711;
  assign n5713 = n1625 & ~n5225;
  assign n5714 = n1553 & ~n5134;
  assign n5715 = ~n5713 & ~n5714;
  assign n5716 = n5712 & ~n5715;
  assign n5717 = n5709 & ~n5716;
  assign n5718 = n5706 & ~n5717;
  assign n5719 = ~n2330 & n5100;
  assign n5720 = ~n2394 & n5078;
  assign n5721 = ~n5719 & ~n5720;
  assign n5722 = ~n2123 & n5330;
  assign n5723 = n2193 & ~n5360;
  assign n5724 = n5722 & ~n5723;
  assign n5725 = n5721 & ~n5724;
  assign n5726 = ~n2050 & n5345;
  assign n5727 = n2123 & ~n5330;
  assign n5728 = ~n5723 & ~n5727;
  assign n5729 = n5726 & n5728;
  assign n5730 = ~n2260 & n5112;
  assign n5731 = ~n2193 & n5360;
  assign n5732 = ~n5730 & ~n5731;
  assign n5733 = n5725 & ~n5729;
  assign n5734 = n5732 & n5733;
  assign n5735 = ~n2604 & n5032;
  assign n5736 = ~n2536 & n5044;
  assign n5737 = n2604 & ~n5032;
  assign n5738 = n5736 & ~n5737;
  assign n5739 = ~n5735 & ~n5738;
  assign n5740 = ~n2467 & n5066;
  assign n5741 = n2536 & ~n5044;
  assign n5742 = ~n5737 & ~n5741;
  assign n5743 = n5740 & n5742;
  assign n5744 = n2784 & n4976;
  assign n5745 = n2722 & n4998;
  assign n5746 = ~n5744 & ~n5745;
  assign n5747 = n2661 & n5010;
  assign n5748 = n5746 & ~n5747;
  assign n5749 = n5739 & ~n5743;
  assign n5750 = n5748 & n5749;
  assign n5751 = n5734 & n5750;
  assign n5752 = n5718 & n5751;
  assign n5753 = ~n1553 & n5134;
  assign n5754 = n5712 & ~n5753;
  assign n5755 = n5706 & n5754;
  assign n5756 = n1487 & ~n5149;
  assign n5757 = n5755 & n5756;
  assign n5758 = n5751 & n5757;
  assign n5759 = ~n5752 & ~n5758;
  assign n5760 = ~n1487 & n5149;
  assign n5761 = n5755 & ~n5760;
  assign n5762 = ~n1422 & n5195;
  assign n5763 = ~n1366 & n5180;
  assign n5764 = ~n5762 & ~n5763;
  assign n5765 = ~n1281 & n5167;
  assign n5766 = n1366 & ~n5180;
  assign n5767 = n5765 & ~n5766;
  assign n5768 = n5764 & ~n5767;
  assign n5769 = n5761 & n5768;
  assign n5770 = n5751 & n5769;
  assign n5771 = ~n5195 & n5761;
  assign n5772 = n5751 & n5771;
  assign n5773 = n1422 & n5772;
  assign n5774 = ~n5696 & ~n5770;
  assign n5775 = ~n5773 & n5774;
  assign n5776 = n2260 & ~n5720;
  assign n5777 = ~n5112 & n5776;
  assign n5778 = ~n5719 & n5777;
  assign n5779 = n5750 & n5778;
  assign n5780 = n2050 & ~n5345;
  assign n5781 = n5751 & n5780;
  assign n5782 = n1983 & ~n5308;
  assign n5783 = n5751 & n5782;
  assign n5784 = ~n5702 & ~n5703;
  assign n5785 = n1913 & ~n5278;
  assign n5786 = n1842 & ~n5293;
  assign n5787 = ~n5785 & ~n5786;
  assign n5788 = n5784 & ~n5787;
  assign n5789 = n5751 & n5788;
  assign n5790 = ~n5779 & ~n5781;
  assign n5791 = ~n5783 & n5790;
  assign n5792 = ~n5789 & n5791;
  assign n5793 = ~n2859 & ~n4964;
  assign n5794 = ~n2784 & ~n4976;
  assign n5795 = ~n5793 & ~n5794;
  assign n5796 = ~n5742 & n5750;
  assign n5797 = n5795 & ~n5796;
  assign n5798 = ~n5728 & n5751;
  assign n5799 = n2394 & ~n5078;
  assign n5800 = n5750 & n5799;
  assign n5801 = n2330 & ~n5100;
  assign n5802 = ~n5720 & n5801;
  assign n5803 = n5750 & n5802;
  assign n5804 = ~n5800 & ~n5803;
  assign n5805 = ~n2722 & ~n4998;
  assign n5806 = ~n5744 & n5805;
  assign n5807 = ~n2661 & ~n5010;
  assign n5808 = n5746 & n5807;
  assign n5809 = ~n5806 & ~n5808;
  assign n5810 = n2467 & ~n5066;
  assign n5811 = n5750 & n5810;
  assign n5812 = n5809 & ~n5811;
  assign n5813 = n5797 & ~n5798;
  assign n5814 = n5804 & n5813;
  assign n5815 = n5812 & n5814;
  assign n5816 = n5759 & n5775;
  assign n5817 = n5792 & n5816;
  assign n5818 = n5815 & n5817;
  assign n5819 = n5699 & ~n5818;
  assign n5820 = n3021 & ~n5819;
  assign n5821 = n3396 & n4846;
  assign n5822 = ~n3413 & ~n4828;
  assign n5823 = ~n3315 & ~n5821;
  assign n5824 = ~n5822 & n5823;
  assign n5825 = ~n5821 & ~n5822;
  assign n5826 = ~n4862 & n5825;
  assign n5827 = ~n5824 & ~n5826;
  assign n5828 = n3164 & n4896;
  assign n5829 = ~n5827 & ~n5828;
  assign n5830 = n3086 & n4908;
  assign n5831 = n5829 & ~n5830;
  assign n5832 = ~n3248 & ~n5828;
  assign n5833 = ~n5827 & n5832;
  assign n5834 = n4874 & ~n5833;
  assign n5835 = n5831 & ~n5834;
  assign n5836 = n4930 & ~n5819;
  assign n5837 = ~n5694 & ~n5820;
  assign n5838 = n5835 & n5837;
  assign n5839 = ~n5836 & n5838;
  assign n5840 = ~n4874 & n5829;
  assign n5841 = ~n5833 & ~n5840;
  assign n5842 = ~n3086 & ~n4908;
  assign n5843 = ~n3164 & ~n4896;
  assign n5844 = ~n5842 & ~n5843;
  assign n5845 = ~n5841 & ~n5844;
  assign n5846 = ~n3396 & ~n4846;
  assign n5847 = ~n5822 & n5846;
  assign n5848 = ~n4862 & n5824;
  assign n5849 = n3413 & n4828;
  assign n5850 = ~n5847 & ~n5848;
  assign n5851 = ~n5849 & n5850;
  assign n5852 = ~n3248 & ~n5827;
  assign n5853 = ~n4874 & n5852;
  assign n5854 = n5851 & ~n5853;
  assign n5855 = ~n5845 & n5854;
  assign n5856 = ~n5839 & n5855;
  assign n5857 = n5693 & n5856;
  assign n5858 = n1333 & ~n5856;
  assign n5859 = n3546 & n5684;
  assign n5860 = n3525 & n5407;
  assign n5861 = ~n5857 & ~n5858;
  assign n5862 = ~n5859 & n5861;
  assign n5863 = ~n5860 & n5862;
  assign n5864 = ~n5469 & ~n5692;
  assign n5865 = n5863 & n5864;
  assign n5866 = ~n1121 & ~n5865;
  assign n5867 = ~n1193 & n4819;
  assign n5868 = n5684 & n5867;
  assign n5869 = ~n5866 & ~n5868;
  assign n5870 = STATE_REG & ~n5869;
  assign n1182 = ~n5410 | n5870;
  assign n5872 = n1134_1 & n1282_1;
  assign n5873 = ~n1183 & ~n1187_1;
  assign n5874 = n1266 & n5873;
  assign n5875 = n5872 & ~n5874;
  assign n5876 = ~n3526 & ~n3944;
  assign n5877 = n1121 & n5876;
  assign n5878 = ~n1342 & n4042;
  assign n5879 = n1197_1 & ~n5878;
  assign n5880 = ~n1333 & ~n3546;
  assign n5881 = n1201 & ~n5880;
  assign n5882 = ~n1331 & ~n3524;
  assign n5883 = ~n5693 & n5882;
  assign n5884 = ~n1325 & ~n5879;
  assign n5885 = ~n5881 & n5884;
  assign n5886 = n5883 & n5885;
  assign n5887 = ~n5874 & ~n5886;
  assign n5888 = n5877 & ~n5887;
  assign n5889 = STATE_REG & ~n5888;
  assign n5890 = ~n5875 & ~n5889;
  assign n5891 = ~n2246 & ~n5890;
  assign n5892 = n5872 & n5874;
  assign n5893 = n1134_1 & n3525;
  assign n5894 = ~n5892 & ~n5893;
  assign n5895 = ~n2330 & ~n5894;
  assign n5896 = n1134_1 & n4811;
  assign n5897 = n1274 & n5874;
  assign n5898 = ~n2321 & n5897;
  assign n5899 = ~n1274 & n5874;
  assign n5900 = ~n2184 & n5899;
  assign n5901 = ~n2246 & ~n5874;
  assign n5902 = ~n5898 & ~n5900;
  assign n5903 = ~n5901 & n5902;
  assign n5904 = n5896 & ~n5903;
  assign n5905 = ~n2184 & ~n4575;
  assign n5906 = ~n2260 & n4567;
  assign n5907 = ~n5905 & ~n5906;
  assign n5908 = ~n2184 & n4567;
  assign n5909 = ~n2260 & ~n4585;
  assign n5910 = ~n5908 & ~n5909;
  assign n5911 = ~n4565 & ~n5910;
  assign n5912 = n4565 & n5910;
  assign n5913 = ~n5911 & ~n5912;
  assign n5914 = ~n5907 & ~n5913;
  assign n5915 = n5907 & n5913;
  assign n5916 = ~n1904 & ~n4575;
  assign n5917 = ~n1983 & n4567;
  assign n5918 = ~n5916 & ~n5917;
  assign n5919 = ~n1904 & n4567;
  assign n5920 = ~n1983 & ~n4585;
  assign n5921 = ~n5919 & ~n5920;
  assign n5922 = ~n4565 & ~n5921;
  assign n5923 = n4565 & n5921;
  assign n5924 = ~n5922 & ~n5923;
  assign n5925 = ~n5918 & ~n5924;
  assign n5926 = ~n2041 & n4567;
  assign n5927 = ~n2123 & ~n4585;
  assign n5928 = ~n5926 & ~n5927;
  assign n5929 = ~n4565 & ~n5928;
  assign n5930 = n4565 & n5928;
  assign n5931 = ~n5929 & ~n5930;
  assign n5932 = ~n2041 & ~n4575;
  assign n5933 = ~n2123 & n4567;
  assign n5934 = ~n5932 & ~n5933;
  assign n5935 = n5931 & n5934;
  assign n5936 = ~n2116 & n4567;
  assign n5937 = ~n2193 & ~n4585;
  assign n5938 = ~n5936 & ~n5937;
  assign n5939 = ~n4565 & ~n5938;
  assign n5940 = n4565 & n5938;
  assign n5941 = ~n5939 & ~n5940;
  assign n5942 = ~n2116 & ~n4575;
  assign n5943 = ~n2193 & n4567;
  assign n5944 = ~n5942 & ~n5943;
  assign n5945 = n5941 & n5944;
  assign n5946 = ~n5935 & ~n5945;
  assign n5947 = ~n1976 & n4567;
  assign n5948 = ~n2050 & ~n4585;
  assign n5949 = ~n5947 & ~n5948;
  assign n5950 = ~n4565 & ~n5949;
  assign n5951 = n4565 & n5949;
  assign n5952 = ~n5950 & ~n5951;
  assign n5953 = ~n1976 & ~n4575;
  assign n5954 = ~n2050 & n4567;
  assign n5955 = ~n5953 & ~n5954;
  assign n5956 = n5952 & n5955;
  assign n5957 = n5946 & ~n5956;
  assign n5958 = n5925 & n5957;
  assign n5959 = ~n5941 & ~n5944;
  assign n5960 = ~n5931 & ~n5934;
  assign n5961 = ~n5959 & ~n5960;
  assign n5962 = ~n5952 & ~n5955;
  assign n5963 = n5946 & n5962;
  assign n5964 = n5961 & ~n5963;
  assign n5965 = ~n5945 & ~n5964;
  assign n5966 = ~n5958 & ~n5965;
  assign n5967 = n5918 & n5924;
  assign n5968 = n5957 & ~n5967;
  assign n5969 = ~n1835 & ~n4575;
  assign n5970 = ~n1913 & n4567;
  assign n5971 = ~n5969 & ~n5970;
  assign n5972 = ~n1684 & ~n4575;
  assign n5973 = ~n1773 & n4567;
  assign n5974 = ~n5972 & ~n5973;
  assign n5975 = ~n1618 & ~n4575;
  assign n5976 = ~n1691 & n4567;
  assign n5977 = ~n5975 & ~n5976;
  assign n5978 = ~n1618 & n4567;
  assign n5979 = ~n1691 & ~n4585;
  assign n5980 = ~n5978 & ~n5979;
  assign n5981 = ~n4565 & ~n5980;
  assign n5982 = n4565 & n5980;
  assign n5983 = ~n5981 & ~n5982;
  assign n5984 = ~n5977 & ~n5983;
  assign n5985 = ~n5974 & n5984;
  assign n5986 = ~n1684 & n4567;
  assign n5987 = ~n1773 & ~n4585;
  assign n5988 = ~n5986 & ~n5987;
  assign n5989 = ~n4565 & ~n5988;
  assign n5990 = n4565 & n5988;
  assign n5991 = ~n5989 & ~n5990;
  assign n5992 = n5974 & ~n5984;
  assign n5993 = ~n5991 & ~n5992;
  assign n5994 = ~n1546 & ~n4575;
  assign n5995 = ~n1625 & n4567;
  assign n5996 = ~n5994 & ~n5995;
  assign n5997 = ~n1546 & n4567;
  assign n5998 = ~n1625 & ~n4585;
  assign n5999 = ~n5997 & ~n5998;
  assign n6000 = ~n4565 & ~n5999;
  assign n6001 = n4565 & n5999;
  assign n6002 = ~n6000 & ~n6001;
  assign n6003 = ~n5996 & ~n6002;
  assign n6004 = n5977 & n5983;
  assign n6005 = n5974 & n5991;
  assign n6006 = ~n6004 & ~n6005;
  assign n6007 = n6003 & n6006;
  assign n6008 = ~n5985 & ~n5993;
  assign n6009 = ~n6007 & n6008;
  assign n6010 = ~n1766 & n4567;
  assign n6011 = ~n1842 & ~n4585;
  assign n6012 = ~n6010 & ~n6011;
  assign n6013 = ~n4565 & ~n6012;
  assign n6014 = n4565 & n6012;
  assign n6015 = ~n6013 & ~n6014;
  assign n6016 = ~n1766 & ~n4575;
  assign n6017 = ~n1842 & n4567;
  assign n6018 = ~n6016 & ~n6017;
  assign n6019 = n6015 & n6018;
  assign n6020 = ~n6009 & ~n6019;
  assign n6021 = ~n6015 & ~n6018;
  assign n6022 = ~n6020 & ~n6021;
  assign n6023 = n5996 & n6002;
  assign n6024 = n6006 & ~n6023;
  assign n6025 = ~n6019 & n6024;
  assign n6026 = ~n1480 & n4567;
  assign n6027 = ~n1553 & ~n4585;
  assign n6028 = ~n6026 & ~n6027;
  assign n6029 = ~n4565 & ~n6028;
  assign n6030 = n4565 & n6028;
  assign n6031 = ~n6029 & ~n6030;
  assign n6032 = ~n1480 & ~n4575;
  assign n6033 = ~n1553 & n4567;
  assign n6034 = ~n6032 & ~n6033;
  assign n6035 = n6031 & n6034;
  assign n6036 = ~n1415 & ~n4575;
  assign n6037 = ~n1487 & n4567;
  assign n6038 = ~n6036 & ~n6037;
  assign n6039 = ~n1359 & ~n4575;
  assign n6040 = ~n1422 & n4567;
  assign n6041 = ~n6039 & ~n6040;
  assign n6042 = ~n1359 & n4567;
  assign n6043 = ~n1422 & ~n4585;
  assign n6044 = ~n6042 & ~n6043;
  assign n6045 = ~n4565 & ~n6044;
  assign n6046 = n4565 & n6044;
  assign n6047 = ~n6045 & ~n6046;
  assign n6048 = ~n6041 & ~n6047;
  assign n6049 = ~n6038 & n6048;
  assign n6050 = ~n1415 & n4567;
  assign n6051 = ~n1487 & ~n4585;
  assign n6052 = ~n6050 & ~n6051;
  assign n6053 = ~n4565 & ~n6052;
  assign n6054 = n4565 & n6052;
  assign n6055 = ~n6053 & ~n6054;
  assign n6056 = n6038 & ~n6048;
  assign n6057 = ~n6055 & ~n6056;
  assign n6058 = ~n6049 & ~n6057;
  assign n6059 = n6041 & n6047;
  assign n6060 = n6038 & n6055;
  assign n6061 = ~n6059 & ~n6060;
  assign n6062 = n4565 & ~n4577;
  assign n6063 = ~n1302_1 & n4567;
  assign n6064 = ~n1366 & ~n4585;
  assign n6065 = ~n6063 & ~n6064;
  assign n6066 = ~n4565 & ~n6065;
  assign n6067 = n4565 & n6065;
  assign n6068 = ~n6066 & ~n6067;
  assign n6069 = ~n1302_1 & ~n4575;
  assign n6070 = ~n1366 & n4567;
  assign n6071 = ~n6069 & ~n6070;
  assign n6072 = n6068 & n6071;
  assign n6073 = n6062 & ~n6072;
  assign n6074 = ~n6068 & ~n6071;
  assign n6075 = ~n4565 & n4577;
  assign n6076 = ~n4590 & ~n6075;
  assign n6077 = ~n6072 & n6076;
  assign n6078 = ~n6073 & ~n6074;
  assign n6079 = ~n6077 & n6078;
  assign n6080 = n6061 & ~n6079;
  assign n6081 = n6058 & ~n6080;
  assign n6082 = ~n6035 & ~n6081;
  assign n6083 = ~n6031 & ~n6034;
  assign n6084 = ~n6082 & ~n6083;
  assign n6085 = n6025 & ~n6084;
  assign n6086 = n6022 & ~n6085;
  assign n6087 = ~n5971 & ~n6086;
  assign n6088 = ~n1835 & n4567;
  assign n6089 = ~n1913 & ~n4585;
  assign n6090 = ~n6088 & ~n6089;
  assign n6091 = ~n4565 & ~n6090;
  assign n6092 = n4565 & n6090;
  assign n6093 = ~n6091 & ~n6092;
  assign n6094 = ~n6086 & ~n6093;
  assign n6095 = ~n5971 & ~n6093;
  assign n6096 = ~n6087 & ~n6094;
  assign n6097 = ~n6095 & n6096;
  assign n6098 = n5968 & ~n6097;
  assign n6099 = n5966 & ~n6098;
  assign n6100 = ~n5915 & ~n6099;
  assign n6101 = ~n5914 & ~n6100;
  assign n6102 = ~n2253 & n4567;
  assign n6103 = ~n2330 & ~n4585;
  assign n6104 = ~n6102 & ~n6103;
  assign n6105 = ~n4565 & ~n6104;
  assign n6106 = n4565 & n6104;
  assign n6107 = ~n6105 & ~n6106;
  assign n6108 = ~n2253 & ~n4575;
  assign n6109 = ~n2330 & n4567;
  assign n6110 = ~n6108 & ~n6109;
  assign n6111 = ~n6107 & n6110;
  assign n6112 = n6107 & ~n6110;
  assign n6113 = ~n6111 & ~n6112;
  assign n6114 = n6101 & ~n6113;
  assign n6115 = ~n6101 & n6113;
  assign n6116 = ~n6114 & ~n6115;
  assign n6117 = n1134_1 & ~n5886;
  assign n6118 = n5874 & n6117;
  assign n6119 = ~n6116 & n6118;
  assign n6120 = ~n5891 & ~n5895;
  assign n6121 = ~n4243 & n6120;
  assign n6122 = ~n5904 & n6121;
  assign n1187 = n6119 | ~n6122;
  assign n6124 = n1282_1 & ~n5874;
  assign n6125 = n5888 & ~n6124;
  assign n6126 = STATE_REG & ~n6125;
  assign n6127 = ~n3013 & n6126;
  assign n6128 = n1282_1 & n5874;
  assign n6129 = ~n3525 & ~n6128;
  assign n6130 = n1134_1 & ~n6129;
  assign n6131 = n3086 & n6130;
  assign n6132 = REG3_REG_26_ & ~STATE_REG;
  assign n6133 = ~n3084 & n5897;
  assign n6134 = ~n2945 & n5899;
  assign n6135 = ~n3013 & ~n5874;
  assign n6136 = ~n6133 & ~n6134;
  assign n6137 = ~n6135 & n6136;
  assign n6138 = n5896 & ~n6137;
  assign n6139 = ~n3017 & ~n4575;
  assign n6140 = n3086 & n4567;
  assign n6141 = ~n6139 & ~n6140;
  assign n6142 = ~n3017 & n4567;
  assign n6143 = n3086 & ~n4585;
  assign n6144 = ~n6142 & ~n6143;
  assign n6145 = ~n4565 & ~n6144;
  assign n6146 = n4565 & n6144;
  assign n6147 = ~n6145 & ~n6146;
  assign n6148 = ~n6141 & ~n6147;
  assign n6149 = ~n2945 & n4567;
  assign n6150 = n3021 & ~n4585;
  assign n6151 = ~n6149 & ~n6150;
  assign n6152 = ~n4565 & ~n6151;
  assign n6153 = n4565 & n6151;
  assign n6154 = ~n6152 & ~n6153;
  assign n6155 = ~n2945 & ~n4575;
  assign n6156 = n3021 & n4567;
  assign n6157 = ~n6155 & ~n6156;
  assign n6158 = n6154 & n6157;
  assign n6159 = n6141 & n6147;
  assign n6160 = ~n6158 & ~n6159;
  assign n6161 = ~n6148 & n6160;
  assign n6162 = ~n2855 & ~n4575;
  assign n6163 = n2947 & n4567;
  assign n6164 = ~n6162 & ~n6163;
  assign n6165 = ~n2855 & n4567;
  assign n6166 = n2947 & ~n4585;
  assign n6167 = ~n6165 & ~n6166;
  assign n6168 = ~n4565 & ~n6167;
  assign n6169 = n4565 & n6167;
  assign n6170 = ~n6168 & ~n6169;
  assign n6171 = ~n6164 & ~n6170;
  assign n6172 = ~n6154 & ~n6157;
  assign n6173 = ~n6171 & ~n6172;
  assign n6174 = n6164 & n6170;
  assign n6175 = ~n2782 & ~n4575;
  assign n6176 = n2859 & n4567;
  assign n6177 = ~n6175 & ~n6176;
  assign n6178 = ~n2782 & n4567;
  assign n6179 = n2859 & ~n4585;
  assign n6180 = ~n6178 & ~n6179;
  assign n6181 = ~n4565 & ~n6180;
  assign n6182 = n4565 & n6180;
  assign n6183 = ~n6181 & ~n6182;
  assign n6184 = ~n6177 & ~n6183;
  assign n6185 = n6177 & n6183;
  assign n6186 = ~n2718 & ~n4575;
  assign n6187 = n2784 & n4567;
  assign n6188 = ~n6186 & ~n6187;
  assign n6189 = ~n2718 & n4567;
  assign n6190 = n2784 & ~n4585;
  assign n6191 = ~n6189 & ~n6190;
  assign n6192 = ~n4565 & ~n6191;
  assign n6193 = n4565 & n6191;
  assign n6194 = ~n6192 & ~n6193;
  assign n6195 = ~n6188 & ~n6194;
  assign n6196 = n6188 & n6194;
  assign n6197 = ~n2659 & n4567;
  assign n6198 = n2722 & ~n4585;
  assign n6199 = ~n6197 & ~n6198;
  assign n6200 = ~n4565 & ~n6199;
  assign n6201 = n4565 & n6199;
  assign n6202 = ~n6200 & ~n6201;
  assign n6203 = ~n2659 & ~n4575;
  assign n6204 = n2722 & n4567;
  assign n6205 = ~n6203 & ~n6204;
  assign n6206 = n6202 & n6205;
  assign n6207 = ~n6202 & ~n6205;
  assign n6208 = ~n2598 & ~n4575;
  assign n6209 = n2661 & n4567;
  assign n6210 = ~n6208 & ~n6209;
  assign n6211 = ~n2598 & n4567;
  assign n6212 = n2661 & ~n4585;
  assign n6213 = ~n6211 & ~n6212;
  assign n6214 = ~n4565 & ~n6213;
  assign n6215 = n4565 & n6213;
  assign n6216 = ~n6214 & ~n6215;
  assign n6217 = ~n6210 & ~n6216;
  assign n6218 = ~n6207 & ~n6217;
  assign n6219 = ~n2529 & ~n4575;
  assign n6220 = ~n2604 & n4567;
  assign n6221 = ~n6219 & ~n6220;
  assign n6222 = ~n2529 & n4567;
  assign n6223 = ~n2604 & ~n4585;
  assign n6224 = ~n6222 & ~n6223;
  assign n6225 = ~n4565 & ~n6224;
  assign n6226 = n4565 & n6224;
  assign n6227 = ~n6225 & ~n6226;
  assign n6228 = ~n6221 & ~n6227;
  assign n6229 = n6210 & n6216;
  assign n6230 = ~n6206 & ~n6229;
  assign n6231 = n6228 & n6230;
  assign n6232 = n6218 & ~n6231;
  assign n6233 = ~n6206 & ~n6232;
  assign n6234 = n6221 & n6227;
  assign n6235 = n6230 & ~n6234;
  assign n6236 = ~n2458 & ~n4575;
  assign n6237 = ~n2536 & n4567;
  assign n6238 = ~n6236 & ~n6237;
  assign n6239 = ~n2458 & n4567;
  assign n6240 = ~n2536 & ~n4585;
  assign n6241 = ~n6239 & ~n6240;
  assign n6242 = ~n4565 & ~n6241;
  assign n6243 = n4565 & n6241;
  assign n6244 = ~n6242 & ~n6243;
  assign n6245 = ~n6238 & ~n6244;
  assign n6246 = n6238 & n6244;
  assign n6247 = ~n2387 & ~n4575;
  assign n6248 = ~n2467 & n4567;
  assign n6249 = ~n6247 & ~n6248;
  assign n6250 = ~n2321 & ~n4575;
  assign n6251 = ~n2394 & n4567;
  assign n6252 = ~n6250 & ~n6251;
  assign n6253 = ~n2321 & n4567;
  assign n6254 = ~n2394 & ~n4585;
  assign n6255 = ~n6253 & ~n6254;
  assign n6256 = ~n4565 & ~n6255;
  assign n6257 = n4565 & n6255;
  assign n6258 = ~n6256 & ~n6257;
  assign n6259 = ~n6252 & ~n6258;
  assign n6260 = ~n6249 & n6259;
  assign n6261 = ~n2387 & n4567;
  assign n6262 = ~n2467 & ~n4585;
  assign n6263 = ~n6261 & ~n6262;
  assign n6264 = ~n4565 & ~n6263;
  assign n6265 = n4565 & n6263;
  assign n6266 = ~n6264 & ~n6265;
  assign n6267 = n6249 & ~n6259;
  assign n6268 = ~n6266 & ~n6267;
  assign n6269 = ~n6260 & ~n6268;
  assign n6270 = n6252 & n6258;
  assign n6271 = n6249 & n6266;
  assign n6272 = ~n6270 & ~n6271;
  assign n6273 = ~n6107 & ~n6110;
  assign n6274 = n6107 & n6110;
  assign n6275 = ~n6101 & ~n6274;
  assign n6276 = ~n6273 & ~n6275;
  assign n6277 = n6272 & ~n6276;
  assign n6278 = n6269 & ~n6277;
  assign n6279 = ~n6246 & ~n6278;
  assign n6280 = ~n6245 & ~n6279;
  assign n6281 = n6235 & ~n6280;
  assign n6282 = ~n6233 & ~n6281;
  assign n6283 = ~n6196 & ~n6282;
  assign n6284 = ~n6195 & ~n6283;
  assign n6285 = ~n6185 & ~n6284;
  assign n6286 = ~n6184 & ~n6285;
  assign n6287 = ~n6174 & ~n6286;
  assign n6288 = n6173 & ~n6287;
  assign n6289 = n6161 & ~n6288;
  assign n6290 = n6141 & ~n6147;
  assign n6291 = ~n6141 & n6147;
  assign n6292 = ~n6290 & ~n6291;
  assign n6293 = ~n6172 & n6292;
  assign n6294 = ~n6171 & ~n6287;
  assign n6295 = ~n6158 & ~n6294;
  assign n6296 = n6293 & ~n6295;
  assign n6297 = ~n6289 & ~n6296;
  assign n6298 = n6118 & n6297;
  assign n6299 = ~n6127 & ~n6131;
  assign n6300 = ~n6132 & n6299;
  assign n6301 = ~n6138 & n6300;
  assign n1192 = n6298 | ~n6301;
  assign n6303 = ~n1611 & ~n5890;
  assign n6304 = ~n1691 & ~n5894;
  assign n6305 = ~n1684 & n5897;
  assign n6306 = ~n1546 & n5899;
  assign n6307 = ~n1611 & ~n5874;
  assign n6308 = ~n6305 & ~n6306;
  assign n6309 = ~n6307 & n6308;
  assign n6310 = n5896 & ~n6309;
  assign n6311 = n5977 & ~n5983;
  assign n6312 = ~n5977 & n5983;
  assign n6313 = ~n6311 & ~n6312;
  assign n6314 = ~n6023 & ~n6084;
  assign n6315 = ~n6003 & ~n6314;
  assign n6316 = ~n6313 & n6315;
  assign n6317 = ~n5984 & ~n6004;
  assign n6318 = ~n6315 & ~n6317;
  assign n6319 = ~n6316 & ~n6318;
  assign n6320 = n6118 & ~n6319;
  assign n6321 = ~n6303 & ~n6304;
  assign n6322 = ~n4493 & n6321;
  assign n6323 = ~n6310 & n6322;
  assign n1197 = n6320 | ~n6323;
  assign n6325 = ~n2451 & ~n5890;
  assign n6326 = ~n2536 & ~n5894;
  assign n6327 = ~n2529 & n5897;
  assign n6328 = ~n2387 & n5899;
  assign n6329 = ~n2451 & ~n5874;
  assign n6330 = ~n6327 & ~n6328;
  assign n6331 = ~n6329 & n6330;
  assign n6332 = n5896 & ~n6331;
  assign n6333 = n6238 & ~n6244;
  assign n6334 = ~n6238 & n6244;
  assign n6335 = ~n6333 & ~n6334;
  assign n6336 = n6278 & ~n6335;
  assign n6337 = ~n6278 & n6335;
  assign n6338 = ~n6336 & ~n6337;
  assign n6339 = n6118 & ~n6338;
  assign n6340 = ~n6325 & ~n6326;
  assign n6341 = ~n4151 & n6340;
  assign n6342 = ~n6332 & n6341;
  assign n1202 = n6339 | ~n6342;
  assign n6344 = n6041 & ~n6047;
  assign n6345 = ~n6041 & n6047;
  assign n6346 = ~n6344 & ~n6345;
  assign n6347 = n6079 & ~n6346;
  assign n6348 = ~n6048 & ~n6059;
  assign n6349 = ~n6079 & ~n6348;
  assign n6350 = ~n6347 & ~n6349;
  assign n6351 = n6118 & ~n6350;
  assign n6352 = ~n4640 & ~n6351;
  assign n6353 = ~n1422 & ~n5894;
  assign n6354 = n6352 & ~n6353;
  assign n6355 = REG3_REG_2_ & ~n5890;
  assign n6356 = ~n1415 & n5897;
  assign n6357 = ~n1302_1 & n5899;
  assign n6358 = REG3_REG_2_ & ~n5874;
  assign n6359 = ~n6356 & ~n6357;
  assign n6360 = ~n6358 & n6359;
  assign n6361 = n5896 & ~n6360;
  assign n6362 = n6354 & ~n6355;
  assign n1207 = n6361 | ~n6362;
  assign n6364 = ~n1969 & ~n5890;
  assign n6365 = ~n2050 & ~n5894;
  assign n6366 = ~n2041 & n5897;
  assign n6367 = ~n1904 & n5899;
  assign n6368 = ~n1969 & ~n5874;
  assign n6369 = ~n6366 & ~n6367;
  assign n6370 = ~n6368 & n6369;
  assign n6371 = n5896 & ~n6370;
  assign n6372 = ~n5967 & ~n6097;
  assign n6373 = ~n5925 & ~n6372;
  assign n6374 = ~n5952 & n5955;
  assign n6375 = n5952 & ~n5955;
  assign n6376 = ~n6374 & ~n6375;
  assign n6377 = n6373 & ~n6376;
  assign n6378 = ~n5956 & ~n5962;
  assign n6379 = ~n6373 & ~n6378;
  assign n6380 = ~n6377 & ~n6379;
  assign n6381 = n6118 & ~n6380;
  assign n6382 = ~n6364 & ~n6365;
  assign n6383 = ~n4349 & n6382;
  assign n6384 = ~n6371 & n6383;
  assign n1212 = n6381 | ~n6384;
  assign n6386 = ~n2714 & n6126;
  assign n6387 = n2784 & n6130;
  assign n6388 = REG3_REG_22_ & ~STATE_REG;
  assign n6389 = ~n2782 & n5897;
  assign n6390 = ~n2659 & n5899;
  assign n6391 = ~n2714 & ~n5874;
  assign n6392 = ~n6389 & ~n6390;
  assign n6393 = ~n6391 & n6392;
  assign n6394 = n5896 & ~n6393;
  assign n6395 = n6188 & ~n6194;
  assign n6396 = ~n6188 & n6194;
  assign n6397 = ~n6395 & ~n6396;
  assign n6398 = n6282 & ~n6397;
  assign n6399 = ~n6282 & n6397;
  assign n6400 = ~n6398 & ~n6399;
  assign n6401 = n6118 & ~n6400;
  assign n6402 = ~n6386 & ~n6387;
  assign n6403 = ~n6388 & n6402;
  assign n6404 = ~n6394 & n6403;
  assign n1217 = n6401 | ~n6404;
  assign n6406 = ~n2109 & ~n5890;
  assign n6407 = ~n2193 & ~n5894;
  assign n6408 = ~n2184 & n5897;
  assign n6409 = ~n2041 & n5899;
  assign n6410 = ~n2109 & ~n5874;
  assign n6411 = ~n6408 & ~n6409;
  assign n6412 = ~n6410 & n6411;
  assign n6413 = n5896 & ~n6412;
  assign n6414 = n5946 & ~n5959;
  assign n6415 = ~n5956 & ~n6373;
  assign n6416 = ~n5962 & ~n6415;
  assign n6417 = ~n5960 & n6416;
  assign n6418 = n6414 & ~n6417;
  assign n6419 = ~n5941 & n5944;
  assign n6420 = n5941 & ~n5944;
  assign n6421 = ~n6419 & ~n6420;
  assign n6422 = ~n5960 & n6421;
  assign n6423 = ~n5935 & ~n6416;
  assign n6424 = n6422 & ~n6423;
  assign n6425 = ~n6418 & ~n6424;
  assign n6426 = n6118 & n6425;
  assign n6427 = ~n6406 & ~n6407;
  assign n6428 = ~n4295 & n6427;
  assign n6429 = ~n6413 & n6428;
  assign n1222 = n6426 | ~n6429;
  assign n6431 = ~n2591 & n6126;
  assign n6432 = n2661 & n6130;
  assign n6433 = REG3_REG_20_ & ~STATE_REG;
  assign n6434 = ~n2659 & n5897;
  assign n6435 = ~n2529 & n5899;
  assign n6436 = ~n2591 & ~n5874;
  assign n6437 = ~n6434 & ~n6435;
  assign n6438 = ~n6436 & n6437;
  assign n6439 = n5896 & ~n6438;
  assign n6440 = n6210 & ~n6216;
  assign n6441 = ~n6210 & n6216;
  assign n6442 = ~n6440 & ~n6441;
  assign n6443 = ~n6234 & ~n6280;
  assign n6444 = ~n6228 & ~n6443;
  assign n6445 = ~n6442 & n6444;
  assign n6446 = ~n6217 & ~n6229;
  assign n6447 = ~n6444 & ~n6446;
  assign n6448 = ~n6445 & ~n6447;
  assign n6449 = n6118 & ~n6448;
  assign n6450 = ~n6431 & ~n6432;
  assign n6451 = ~n6433 & n6450;
  assign n6452 = ~n6439 & n6451;
  assign n1227 = n6449 | ~n6452;
  assign n6454 = ~n4593 & n6118;
  assign n6455 = ~n4704 & ~n6454;
  assign n6456 = ~n5872 & ~n5896;
  assign n6457 = ~n5874 & ~n6456;
  assign n6458 = ~n5889 & ~n6457;
  assign n6459 = REG3_REG_0_ & ~n6458;
  assign n6460 = ~n1281 & ~n5894;
  assign n6461 = ~n1302_1 & n5896;
  assign n6462 = n5897 & n6461;
  assign n6463 = ~n6460 & ~n6462;
  assign n6464 = n6455 & ~n6459;
  assign n1232 = ~n6463 | ~n6464;
  assign n6466 = ~n1828 & ~n5890;
  assign n6467 = ~n1913 & ~n5894;
  assign n6468 = ~n1904 & n5897;
  assign n6469 = ~n1766 & n5899;
  assign n6470 = ~n1828 & ~n5874;
  assign n6471 = ~n6468 & ~n6469;
  assign n6472 = ~n6470 & n6471;
  assign n6473 = n5896 & ~n6472;
  assign n6474 = n5971 & ~n6093;
  assign n6475 = ~n5971 & n6093;
  assign n6476 = ~n6474 & ~n6475;
  assign n6477 = n6086 & ~n6476;
  assign n6478 = ~n6086 & n6476;
  assign n6479 = ~n6477 & ~n6478;
  assign n6480 = n6118 & ~n6479;
  assign n6481 = ~n6466 & ~n6467;
  assign n6482 = ~n4403 & n6481;
  assign n6483 = ~n6473 & n6482;
  assign n1237 = n6480 | ~n6483;
  assign n6485 = ~n1473 & ~n5890;
  assign n6486 = ~n1553 & ~n5894;
  assign n6487 = ~n6031 & n6034;
  assign n6488 = n6031 & ~n6034;
  assign n6489 = ~n6487 & ~n6488;
  assign n6490 = n6081 & ~n6489;
  assign n6491 = ~n6081 & n6489;
  assign n6492 = ~n6490 & ~n6491;
  assign n6493 = n6118 & ~n6492;
  assign n6494 = ~n4540 & ~n6493;
  assign n6495 = ~n1546 & n5897;
  assign n6496 = ~n1415 & n5899;
  assign n6497 = ~n1473 & ~n5874;
  assign n6498 = ~n6495 & ~n6496;
  assign n6499 = ~n6497 & n6498;
  assign n6500 = n5896 & ~n6499;
  assign n6501 = ~n6485 & ~n6486;
  assign n6502 = n6494 & n6501;
  assign n1242 = n6500 | ~n6502;
  assign n6504 = ~n2851 & n6126;
  assign n6505 = n2947 & n6130;
  assign n6506 = REG3_REG_24_ & ~STATE_REG;
  assign n6507 = ~n2945 & n5897;
  assign n6508 = ~n2782 & n5899;
  assign n6509 = ~n2851 & ~n5874;
  assign n6510 = ~n6507 & ~n6508;
  assign n6511 = ~n6509 & n6510;
  assign n6512 = n5896 & ~n6511;
  assign n6513 = n6164 & ~n6170;
  assign n6514 = ~n6164 & n6170;
  assign n6515 = ~n6513 & ~n6514;
  assign n6516 = n6286 & ~n6515;
  assign n6517 = ~n6171 & ~n6174;
  assign n6518 = ~n6286 & ~n6517;
  assign n6519 = ~n6516 & ~n6518;
  assign n6520 = n6118 & ~n6519;
  assign n6521 = ~n6504 & ~n6505;
  assign n6522 = ~n6506 & n6521;
  assign n6523 = ~n6512 & n6522;
  assign n1247 = n6520 | ~n6523;
  assign n6525 = ~n2380 & ~n5890;
  assign n6526 = ~n2467 & ~n5894;
  assign n6527 = ~n2458 & n5897;
  assign n6528 = ~n2321 & n5899;
  assign n6529 = ~n2380 & ~n5874;
  assign n6530 = ~n6527 & ~n6528;
  assign n6531 = ~n6529 & n6530;
  assign n6532 = n5896 & ~n6531;
  assign n6533 = ~n6249 & ~n6266;
  assign n6534 = n6272 & ~n6533;
  assign n6535 = ~n6259 & n6276;
  assign n6536 = n6534 & ~n6535;
  assign n6537 = n6249 & ~n6266;
  assign n6538 = ~n6249 & n6266;
  assign n6539 = ~n6537 & ~n6538;
  assign n6540 = ~n6259 & n6539;
  assign n6541 = ~n6270 & ~n6276;
  assign n6542 = n6540 & ~n6541;
  assign n6543 = ~n6536 & ~n6542;
  assign n6544 = n6118 & n6543;
  assign n6545 = ~n6525 & ~n6526;
  assign n6546 = ~n4187 & n6545;
  assign n6547 = ~n6532 & n6546;
  assign n1252 = n6544 | ~n6547;
  assign n6549 = ~n1539 & ~n5890;
  assign n6550 = ~n1625 & ~n5894;
  assign n6551 = ~n1618 & n5897;
  assign n6552 = ~n1480 & n5899;
  assign n6553 = ~n1539 & ~n5874;
  assign n6554 = ~n6551 & ~n6552;
  assign n6555 = ~n6553 & n6554;
  assign n6556 = n5896 & ~n6555;
  assign n6557 = n5996 & ~n6002;
  assign n6558 = ~n5996 & n6002;
  assign n6559 = ~n6557 & ~n6558;
  assign n6560 = n6084 & ~n6559;
  assign n6561 = ~n6084 & n6559;
  assign n6562 = ~n6560 & ~n6561;
  assign n6563 = n6118 & ~n6562;
  assign n6564 = ~n4519 & ~n6563;
  assign n6565 = ~n6549 & ~n6550;
  assign n6566 = ~n6556 & n6565;
  assign n1257 = ~n6564 | ~n6566;
  assign n6568 = ~n2314 & ~n5890;
  assign n6569 = ~n2394 & ~n5894;
  assign n6570 = ~n2387 & n5897;
  assign n6571 = ~n2253 & n5899;
  assign n6572 = ~n2314 & ~n5874;
  assign n6573 = ~n6570 & ~n6571;
  assign n6574 = ~n6572 & n6573;
  assign n6575 = n5896 & ~n6574;
  assign n6576 = n6252 & ~n6258;
  assign n6577 = ~n6252 & n6258;
  assign n6578 = ~n6576 & ~n6577;
  assign n6579 = n6276 & ~n6578;
  assign n6580 = ~n6259 & ~n6270;
  assign n6581 = ~n6276 & ~n6580;
  assign n6582 = ~n6579 & ~n6581;
  assign n6583 = n6118 & ~n6582;
  assign n6584 = ~n6568 & ~n6569;
  assign n6585 = ~n4215 & n6584;
  assign n6586 = ~n6575 & n6585;
  assign n1262 = n6583 | ~n6586;
  assign n6588 = ~n2941 & n6126;
  assign n6589 = n3021 & n6130;
  assign n6590 = REG3_REG_25_ & ~STATE_REG;
  assign n6591 = ~n3017 & n5897;
  assign n6592 = ~n2855 & n5899;
  assign n6593 = ~n2941 & ~n5874;
  assign n6594 = ~n6591 & ~n6592;
  assign n6595 = ~n6593 & n6594;
  assign n6596 = n5896 & ~n6595;
  assign n6597 = ~n6154 & n6157;
  assign n6598 = n6154 & ~n6157;
  assign n6599 = ~n6597 & ~n6598;
  assign n6600 = n6294 & ~n6599;
  assign n6601 = ~n6158 & ~n6172;
  assign n6602 = ~n6294 & ~n6601;
  assign n6603 = ~n6600 & ~n6602;
  assign n6604 = n6118 & ~n6603;
  assign n6605 = ~n6588 & ~n6589;
  assign n6606 = ~n6590 & n6605;
  assign n6607 = ~n6596 & n6606;
  assign n1267 = n6604 | ~n6607;
  assign n6609 = ~n2034 & ~n5890;
  assign n6610 = ~n2123 & ~n5894;
  assign n6611 = ~n2116 & n5897;
  assign n6612 = ~n1976 & n5899;
  assign n6613 = ~n2034 & ~n5874;
  assign n6614 = ~n6611 & ~n6612;
  assign n6615 = ~n6613 & n6614;
  assign n6616 = n5896 & ~n6615;
  assign n6617 = ~n5931 & n5934;
  assign n6618 = n5931 & ~n5934;
  assign n6619 = ~n6617 & ~n6618;
  assign n6620 = n6416 & ~n6619;
  assign n6621 = ~n5935 & ~n5960;
  assign n6622 = ~n6416 & ~n6621;
  assign n6623 = ~n6620 & ~n6622;
  assign n6624 = n6118 & ~n6623;
  assign n6625 = ~n6609 & ~n6610;
  assign n6626 = ~n4321 & n6625;
  assign n6627 = ~n6616 & n6626;
  assign n1272 = n6624 | ~n6627;
  assign n6629 = ~n2655 & n6126;
  assign n6630 = n2722 & n6130;
  assign n6631 = REG3_REG_21_ & ~STATE_REG;
  assign n6632 = ~n2718 & n5897;
  assign n6633 = ~n2598 & n5899;
  assign n6634 = ~n2655 & ~n5874;
  assign n6635 = ~n6632 & ~n6633;
  assign n6636 = ~n6634 & n6635;
  assign n6637 = n5896 & ~n6636;
  assign n6638 = ~n6207 & n6230;
  assign n6639 = ~n6217 & n6444;
  assign n6640 = n6638 & ~n6639;
  assign n6641 = ~n6202 & n6205;
  assign n6642 = n6202 & ~n6205;
  assign n6643 = ~n6641 & ~n6642;
  assign n6644 = ~n6217 & n6643;
  assign n6645 = ~n6229 & ~n6444;
  assign n6646 = n6644 & ~n6645;
  assign n6647 = ~n6640 & ~n6646;
  assign n6648 = n6118 & n6647;
  assign n6649 = ~n6629 & ~n6630;
  assign n6650 = ~n6631 & n6649;
  assign n6651 = ~n6637 & n6650;
  assign n1277 = n6648 | ~n6651;
  assign n6653 = ~n6062 & ~n6076;
  assign n6654 = ~n6068 & n6071;
  assign n6655 = n6068 & ~n6071;
  assign n6656 = ~n6654 & ~n6655;
  assign n6657 = n6653 & ~n6656;
  assign n6658 = ~n6653 & n6656;
  assign n6659 = ~n6657 & ~n6658;
  assign n6660 = n6118 & ~n6659;
  assign n6661 = ~n4682 & ~n6660;
  assign n6662 = ~n1366 & ~n5894;
  assign n6663 = n6661 & ~n6662;
  assign n6664 = REG3_REG_1_ & ~n5890;
  assign n6665 = ~n1359 & n5897;
  assign n6666 = ~n1313 & n5899;
  assign n6667 = REG3_REG_1_ & ~n5874;
  assign n6668 = ~n6665 & ~n6666;
  assign n6669 = ~n6667 & n6668;
  assign n6670 = n5896 & ~n6669;
  assign n6671 = n6663 & ~n6664;
  assign n1282 = n6670 | ~n6671;
  assign n6673 = ~n1759 & ~n5890;
  assign n6674 = ~n1842 & ~n5894;
  assign n6675 = ~n1835 & n5897;
  assign n6676 = ~n1684 & n5899;
  assign n6677 = ~n1759 & ~n5874;
  assign n6678 = ~n6675 & ~n6676;
  assign n6679 = ~n6677 & n6678;
  assign n6680 = n5896 & ~n6679;
  assign n6681 = n6024 & ~n6084;
  assign n6682 = n6009 & ~n6681;
  assign n6683 = ~n6015 & n6018;
  assign n6684 = n6015 & ~n6018;
  assign n6685 = ~n6683 & ~n6684;
  assign n6686 = n6682 & ~n6685;
  assign n6687 = ~n6682 & n6685;
  assign n6688 = ~n6686 & ~n6687;
  assign n6689 = n6118 & ~n6688;
  assign n6690 = ~n6673 & ~n6674;
  assign n6691 = ~n4431 & n6690;
  assign n6692 = ~n6680 & n6691;
  assign n1287 = n6689 | ~n6692;
  assign n6694 = ~n3156 & n6126;
  assign n6695 = n3248 & n6130;
  assign n6696 = REG3_REG_28_ & ~STATE_REG;
  assign n6697 = ~n3246 & n5897;
  assign n6698 = ~n3084 & n5899;
  assign n6699 = ~n3156 & ~n5874;
  assign n6700 = ~n6697 & ~n6698;
  assign n6701 = ~n6699 & n6700;
  assign n6702 = n5896 & ~n6701;
  assign n6703 = ~n3084 & ~n4575;
  assign n6704 = n3164 & n4567;
  assign n6705 = ~n6703 & ~n6704;
  assign n6706 = ~n3084 & n4567;
  assign n6707 = n3164 & ~n4585;
  assign n6708 = ~n6706 & ~n6707;
  assign n6709 = ~n4565 & ~n6708;
  assign n6710 = n4565 & n6708;
  assign n6711 = ~n6709 & ~n6710;
  assign n6712 = ~n6705 & ~n6711;
  assign n6713 = n6705 & n6711;
  assign n6714 = ~n6148 & ~n6172;
  assign n6715 = n6160 & n6171;
  assign n6716 = n6714 & ~n6715;
  assign n6717 = ~n6159 & ~n6716;
  assign n6718 = n6160 & ~n6174;
  assign n6719 = ~n6286 & n6718;
  assign n6720 = ~n6717 & ~n6719;
  assign n6721 = ~n6713 & ~n6720;
  assign n6722 = ~n3160 & ~n4575;
  assign n6723 = n3248 & n4567;
  assign n6724 = ~n6722 & ~n6723;
  assign n6725 = ~n4565 & ~n6724;
  assign n6726 = n4565 & n6724;
  assign n6727 = ~n6725 & ~n6726;
  assign n6728 = ~n3160 & n4567;
  assign n6729 = n3248 & ~n4585;
  assign n6730 = ~n6728 & ~n6729;
  assign n6731 = ~n6727 & n6730;
  assign n6732 = n6727 & ~n6730;
  assign n6733 = ~n6731 & ~n6732;
  assign n6734 = ~n6712 & ~n6721;
  assign n6735 = ~n6733 & n6734;
  assign n6736 = ~n6712 & ~n6717;
  assign n6737 = ~n6719 & n6736;
  assign n6738 = ~n6713 & ~n6737;
  assign n6739 = n6733 & n6738;
  assign n6740 = ~n6735 & ~n6739;
  assign n6741 = n6118 & ~n6740;
  assign n6742 = ~n6694 & ~n6695;
  assign n6743 = ~n6696 & n6742;
  assign n6744 = ~n6702 & n6743;
  assign n1292 = n6741 | ~n6744;
  assign n6746 = ~n2522 & ~n5890;
  assign n6747 = ~n2604 & ~n5894;
  assign n6748 = ~n2598 & n5897;
  assign n6749 = ~n2458 & n5899;
  assign n6750 = ~n2522 & ~n5874;
  assign n6751 = ~n6748 & ~n6749;
  assign n6752 = ~n6750 & n6751;
  assign n6753 = n5896 & ~n6752;
  assign n6754 = n6221 & ~n6227;
  assign n6755 = ~n6221 & n6227;
  assign n6756 = ~n6754 & ~n6755;
  assign n6757 = n6280 & ~n6756;
  assign n6758 = ~n6228 & ~n6234;
  assign n6759 = ~n6280 & ~n6758;
  assign n6760 = ~n6757 & ~n6759;
  assign n6761 = n6118 & ~n6760;
  assign n6762 = ~n6746 & ~n6747;
  assign n6763 = ~n3954 & n6762;
  assign n6764 = ~n6753 & n6763;
  assign n1297 = n6761 | ~n6764;
  assign n6766 = ~n6038 & ~n6055;
  assign n6767 = n6061 & ~n6766;
  assign n6768 = ~n6048 & n6079;
  assign n6769 = n6767 & ~n6768;
  assign n6770 = n6038 & ~n6055;
  assign n6771 = ~n6038 & n6055;
  assign n6772 = ~n6770 & ~n6771;
  assign n6773 = ~n6048 & n6772;
  assign n6774 = ~n6059 & ~n6079;
  assign n6775 = n6773 & ~n6774;
  assign n6776 = ~n6769 & ~n6775;
  assign n6777 = n6118 & n6776;
  assign n6778 = ~n4619 & ~n6777;
  assign n6779 = ~n1487 & ~n5894;
  assign n6780 = n6778 & ~n6779;
  assign n6781 = ~REG3_REG_3_ & ~n5890;
  assign n6782 = ~n1480 & n5897;
  assign n6783 = ~n1359 & n5899;
  assign n6784 = ~REG3_REG_3_ & ~n5874;
  assign n6785 = ~n6782 & ~n6783;
  assign n6786 = ~n6784 & n6785;
  assign n6787 = n5896 & ~n6786;
  assign n6788 = n6780 & ~n6781;
  assign n1302 = n6787 | ~n6788;
  assign n6790 = ~n1897 & ~n5890;
  assign n6791 = ~n1983 & ~n5894;
  assign n6792 = ~n1976 & n5897;
  assign n6793 = ~n1835 & n5899;
  assign n6794 = ~n1897 & ~n5874;
  assign n6795 = ~n6792 & ~n6793;
  assign n6796 = ~n6794 & n6795;
  assign n6797 = n5896 & ~n6796;
  assign n6798 = n5918 & ~n5924;
  assign n6799 = ~n5918 & n5924;
  assign n6800 = ~n6798 & ~n6799;
  assign n6801 = n6097 & ~n6800;
  assign n6802 = ~n6097 & n6800;
  assign n6803 = ~n6801 & ~n6802;
  assign n6804 = n6118 & ~n6803;
  assign n6805 = ~n6790 & ~n6791;
  assign n6806 = ~n4377 & n6805;
  assign n6807 = ~n6797 & n6806;
  assign n1307 = n6804 | ~n6807;
  assign n6809 = ~n2778 & n6126;
  assign n6810 = n2859 & n6130;
  assign n6811 = REG3_REG_23_ & ~STATE_REG;
  assign n6812 = ~n2855 & n5897;
  assign n6813 = ~n2718 & n5899;
  assign n6814 = ~n2778 & ~n5874;
  assign n6815 = ~n6812 & ~n6813;
  assign n6816 = ~n6814 & n6815;
  assign n6817 = n5896 & ~n6816;
  assign n6818 = n6177 & ~n6183;
  assign n6819 = ~n6177 & n6183;
  assign n6820 = ~n6818 & ~n6819;
  assign n6821 = n6284 & ~n6820;
  assign n6822 = ~n6284 & n6820;
  assign n6823 = ~n6821 & ~n6822;
  assign n6824 = n6118 & ~n6823;
  assign n6825 = ~n6809 & ~n6810;
  assign n6826 = ~n6811 & n6825;
  assign n6827 = ~n6817 & n6826;
  assign n1312 = n6824 | ~n6827;
  assign n6829 = ~n2177 & ~n5890;
  assign n6830 = ~n2260 & ~n5894;
  assign n6831 = ~n2253 & n5897;
  assign n6832 = ~n2116 & n5899;
  assign n6833 = ~n2177 & ~n5874;
  assign n6834 = ~n6831 & ~n6832;
  assign n6835 = ~n6833 & n6834;
  assign n6836 = n5896 & ~n6835;
  assign n6837 = n5907 & ~n5913;
  assign n6838 = ~n5907 & n5913;
  assign n6839 = ~n6837 & ~n6838;
  assign n6840 = n6099 & ~n6839;
  assign n6841 = ~n6099 & n6839;
  assign n6842 = ~n6840 & ~n6841;
  assign n6843 = n6118 & ~n6842;
  assign n6844 = ~n6829 & ~n6830;
  assign n6845 = ~n4269 & n6844;
  assign n6846 = ~n6836 & n6845;
  assign n1317 = n6843 | ~n6846;
  assign n6848 = ~n3080 & n6126;
  assign n6849 = n3164 & n6130;
  assign n6850 = REG3_REG_27_ & ~STATE_REG;
  assign n6851 = ~n3160 & n5897;
  assign n6852 = ~n3017 & n5899;
  assign n6853 = ~n3080 & ~n5874;
  assign n6854 = ~n6851 & ~n6852;
  assign n6855 = ~n6853 & n6854;
  assign n6856 = n5896 & ~n6855;
  assign n6857 = n6705 & ~n6711;
  assign n6858 = ~n6705 & n6711;
  assign n6859 = ~n6857 & ~n6858;
  assign n6860 = n6720 & ~n6859;
  assign n6861 = ~n6720 & n6859;
  assign n6862 = ~n6860 & ~n6861;
  assign n6863 = n6118 & ~n6862;
  assign n6864 = ~n6848 & ~n6849;
  assign n6865 = ~n6850 & n6864;
  assign n6866 = ~n6856 & n6865;
  assign n1322 = n6863 | ~n6866;
  assign n6868 = ~n1677 & ~n5890;
  assign n6869 = ~n1773 & ~n5894;
  assign n6870 = ~n1766 & n5897;
  assign n6871 = ~n1618 & n5899;
  assign n6872 = ~n1677 & ~n5874;
  assign n6873 = ~n6870 & ~n6871;
  assign n6874 = ~n6872 & n6873;
  assign n6875 = n5896 & ~n6874;
  assign n6876 = ~n5974 & ~n5991;
  assign n6877 = n6006 & ~n6876;
  assign n6878 = ~n5984 & n6315;
  assign n6879 = n6877 & ~n6878;
  assign n6880 = n5974 & ~n5991;
  assign n6881 = ~n5974 & n5991;
  assign n6882 = ~n6880 & ~n6881;
  assign n6883 = ~n5984 & n6882;
  assign n6884 = ~n6004 & ~n6315;
  assign n6885 = n6883 & ~n6884;
  assign n6886 = ~n6879 & ~n6885;
  assign n6887 = n6118 & n6886;
  assign n6888 = ~n6868 & ~n6869;
  assign n6889 = ~n4465 & n6888;
  assign n6890 = ~n6875 & n6889;
  assign n1327 = n6887 | ~n6890;
  assign n1332 = ~STATE_REG;
  always @ (posedge clock) begin
    IR_REG_0_ <= n174;
    IR_REG_1_ <= n179;
    IR_REG_2_ <= n184;
    IR_REG_3_ <= n189;
    IR_REG_4_ <= n194;
    IR_REG_5_ <= n199;
    IR_REG_6_ <= n204;
    IR_REG_7_ <= n209;
    IR_REG_8_ <= n214;
    IR_REG_9_ <= n219;
    IR_REG_10_ <= n224;
    IR_REG_11_ <= n229;
    IR_REG_12_ <= n234;
    IR_REG_13_ <= n239;
    IR_REG_14_ <= n244;
    IR_REG_15_ <= n249;
    IR_REG_16_ <= n254;
    IR_REG_17_ <= n259;
    IR_REG_18_ <= n264;
    IR_REG_19_ <= n269;
    IR_REG_20_ <= n274;
    IR_REG_21_ <= n279;
    IR_REG_22_ <= n284;
    IR_REG_23_ <= n289;
    IR_REG_24_ <= n294;
    IR_REG_25_ <= n299;
    IR_REG_26_ <= n304;
    IR_REG_27_ <= n309;
    IR_REG_28_ <= n314;
    IR_REG_29_ <= n319;
    IR_REG_30_ <= n324;
    IR_REG_31_ <= n329;
    D_REG_0_ <= n334;
    D_REG_1_ <= n339;
    D_REG_2_ <= n344;
    D_REG_3_ <= n349;
    D_REG_4_ <= n354;
    D_REG_5_ <= n359;
    D_REG_6_ <= n364;
    D_REG_7_ <= n369;
    D_REG_8_ <= n374;
    D_REG_9_ <= n379;
    D_REG_10_ <= n384;
    D_REG_11_ <= n389;
    D_REG_12_ <= n394;
    D_REG_13_ <= n399;
    D_REG_14_ <= n404;
    D_REG_15_ <= n409;
    D_REG_16_ <= n414;
    D_REG_17_ <= n419;
    D_REG_18_ <= n424;
    D_REG_19_ <= n429;
    D_REG_20_ <= n434;
    D_REG_21_ <= n439;
    D_REG_22_ <= n444;
    D_REG_23_ <= n449;
    D_REG_24_ <= n454;
    D_REG_25_ <= n459;
    D_REG_26_ <= n464;
    D_REG_27_ <= n469;
    D_REG_28_ <= n474;
    D_REG_29_ <= n479;
    D_REG_30_ <= n484;
    D_REG_31_ <= n489;
    REG0_REG_0_ <= n494;
    REG0_REG_1_ <= n499;
    REG0_REG_2_ <= n504;
    REG0_REG_3_ <= n509;
    REG0_REG_4_ <= n514;
    REG0_REG_5_ <= n519;
    REG0_REG_6_ <= n524;
    REG0_REG_7_ <= n529;
    REG0_REG_8_ <= n534;
    REG0_REG_9_ <= n539;
    REG0_REG_10_ <= n544;
    REG0_REG_11_ <= n549;
    REG0_REG_12_ <= n554;
    REG0_REG_13_ <= n559;
    REG0_REG_14_ <= n564;
    REG0_REG_15_ <= n569;
    REG0_REG_16_ <= n574;
    REG0_REG_17_ <= n579;
    REG0_REG_18_ <= n584;
    REG0_REG_19_ <= n589;
    REG0_REG_20_ <= n594;
    REG0_REG_21_ <= n599;
    REG0_REG_22_ <= n604;
    REG0_REG_23_ <= n609;
    REG0_REG_24_ <= n614;
    REG0_REG_25_ <= n619;
    REG0_REG_26_ <= n624;
    REG0_REG_27_ <= n629;
    REG0_REG_28_ <= n634;
    REG0_REG_29_ <= n639;
    REG0_REG_30_ <= n644;
    REG0_REG_31_ <= n649;
    REG1_REG_0_ <= n654;
    REG1_REG_1_ <= n659;
    REG1_REG_2_ <= n664;
    REG1_REG_3_ <= n669;
    REG1_REG_4_ <= n674;
    REG1_REG_5_ <= n679;
    REG1_REG_6_ <= n684;
    REG1_REG_7_ <= n689;
    REG1_REG_8_ <= n694;
    REG1_REG_9_ <= n699;
    REG1_REG_10_ <= n704;
    REG1_REG_11_ <= n709;
    REG1_REG_12_ <= n714;
    REG1_REG_13_ <= n719;
    REG1_REG_14_ <= n724;
    REG1_REG_15_ <= n729;
    REG1_REG_16_ <= n734;
    REG1_REG_17_ <= n739;
    REG1_REG_18_ <= n744;
    REG1_REG_19_ <= n749;
    REG1_REG_20_ <= n754;
    REG1_REG_21_ <= n759;
    REG1_REG_22_ <= n764;
    REG1_REG_23_ <= n769;
    REG1_REG_24_ <= n774;
    REG1_REG_25_ <= n779;
    REG1_REG_26_ <= n784;
    REG1_REG_27_ <= n789;
    REG1_REG_28_ <= n794;
    REG1_REG_29_ <= n799;
    REG1_REG_30_ <= n804;
    REG1_REG_31_ <= n809;
    REG2_REG_0_ <= n814;
    REG2_REG_1_ <= n819;
    REG2_REG_2_ <= n824;
    REG2_REG_3_ <= n829;
    REG2_REG_4_ <= n834;
    REG2_REG_5_ <= n839;
    REG2_REG_6_ <= n844;
    REG2_REG_7_ <= n849;
    REG2_REG_8_ <= n854;
    REG2_REG_9_ <= n859;
    REG2_REG_10_ <= n864;
    REG2_REG_11_ <= n869;
    REG2_REG_12_ <= n874;
    REG2_REG_13_ <= n879;
    REG2_REG_14_ <= n884;
    REG2_REG_15_ <= n889;
    REG2_REG_16_ <= n894;
    REG2_REG_17_ <= n899;
    REG2_REG_18_ <= n904;
    REG2_REG_19_ <= n909;
    REG2_REG_20_ <= n914;
    REG2_REG_21_ <= n919;
    REG2_REG_22_ <= n924;
    REG2_REG_23_ <= n929;
    REG2_REG_24_ <= n934;
    REG2_REG_25_ <= n939;
    REG2_REG_26_ <= n944;
    REG2_REG_27_ <= n949;
    REG2_REG_28_ <= n954;
    REG2_REG_29_ <= n959;
    REG2_REG_30_ <= n964;
    REG2_REG_31_ <= n969;
    ADDR_REG_19_ <= n974;
    ADDR_REG_18_ <= n978;
    ADDR_REG_17_ <= n982;
    ADDR_REG_16_ <= n986;
    ADDR_REG_15_ <= n990;
    ADDR_REG_14_ <= n994;
    ADDR_REG_13_ <= n998;
    ADDR_REG_12_ <= n1002;
    ADDR_REG_11_ <= n1006;
    ADDR_REG_10_ <= n1010;
    ADDR_REG_9_ <= n1014;
    ADDR_REG_8_ <= n1018;
    ADDR_REG_7_ <= n1022;
    ADDR_REG_6_ <= n1026;
    ADDR_REG_5_ <= n1030;
    ADDR_REG_4_ <= n1034;
    ADDR_REG_3_ <= n1038;
    ADDR_REG_2_ <= n1042;
    ADDR_REG_1_ <= n1046;
    ADDR_REG_0_ <= n1050;
    DATAO_REG_0_ <= n1054;
    DATAO_REG_1_ <= n1058;
    DATAO_REG_2_ <= n1062;
    DATAO_REG_3_ <= n1066;
    DATAO_REG_4_ <= n1070;
    DATAO_REG_5_ <= n1074;
    DATAO_REG_6_ <= n1078;
    DATAO_REG_7_ <= n1082;
    DATAO_REG_8_ <= n1086;
    DATAO_REG_9_ <= n1090;
    DATAO_REG_10_ <= n1094;
    DATAO_REG_11_ <= n1098;
    DATAO_REG_12_ <= n1102;
    DATAO_REG_13_ <= n1106;
    DATAO_REG_14_ <= n1110;
    DATAO_REG_15_ <= n1114;
    DATAO_REG_16_ <= n1118;
    DATAO_REG_17_ <= n1122;
    DATAO_REG_18_ <= n1126;
    DATAO_REG_19_ <= n1130;
    DATAO_REG_20_ <= n1134;
    DATAO_REG_21_ <= n1138;
    DATAO_REG_22_ <= n1142;
    DATAO_REG_23_ <= n1146;
    DATAO_REG_24_ <= n1150;
    DATAO_REG_25_ <= n1154;
    DATAO_REG_26_ <= n1158;
    DATAO_REG_27_ <= n1162;
    DATAO_REG_28_ <= n1166;
    DATAO_REG_29_ <= n1170;
    DATAO_REG_30_ <= n1174;
    DATAO_REG_31_ <= n1178;
    B_REG <= n1182;
    REG3_REG_15_ <= n1187;
    REG3_REG_26_ <= n1192;
    REG3_REG_6_ <= n1197;
    REG3_REG_18_ <= n1202;
    REG3_REG_2_ <= n1207;
    REG3_REG_11_ <= n1212;
    REG3_REG_22_ <= n1217;
    REG3_REG_13_ <= n1222;
    REG3_REG_20_ <= n1227;
    REG3_REG_0_ <= n1232;
    REG3_REG_9_ <= n1237;
    REG3_REG_4_ <= n1242;
    REG3_REG_24_ <= n1247;
    REG3_REG_17_ <= n1252;
    REG3_REG_5_ <= n1257;
    REG3_REG_16_ <= n1262;
    REG3_REG_25_ <= n1267;
    REG3_REG_12_ <= n1272;
    REG3_REG_21_ <= n1277;
    REG3_REG_1_ <= n1282;
    REG3_REG_8_ <= n1287;
    REG3_REG_28_ <= n1292;
    REG3_REG_19_ <= n1297;
    REG3_REG_3_ <= n1302;
    REG3_REG_10_ <= n1307;
    REG3_REG_23_ <= n1312;
    REG3_REG_14_ <= n1317;
    REG3_REG_27_ <= n1322;
    REG3_REG_7_ <= n1327;
    STATE_REG <= n1332;
    RD_REG <= n1337;
    WR_REG <= n1341;
  end
endmodule


