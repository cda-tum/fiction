// Benchmark "top" written by ABC on Mon Feb 19 11:52:42 2024

module top ( 
    _77_9_, _87_10_, _169_22_, _238_31_, _2897_49_, _68_8_, _128_16_,
    _226_29_, _294_39_, _326_44_, _58_7_, _190_24_, _264_35_, _283_38_,
    _250_33_, _329_45_, _213_26_, _257_34_, _20_2_, _223_28_, _159_21_,
    _232_30_, _41_4_, _124_14_, _13_1_, _50_6_, _222_27_, _97_11_,
    _125_15_, _322_43_, _244_32_, _274_37_, _317_42_, _1_0_, _33_3_,
    _270_36_, _200_25_, _343_47_, _330_46_, _1698_48_, _132_17_, _45_5_,
    _116_13_, _143_19_, _303_40_, _311_41_, _107_12_, _137_18_, _150_20_,
    _179_23_,
    _381_1626_, _351_1247_, _353_405_, _375_1624_, _393_1605_, _364_1484_,
    _369_1321_, _384_1553_, _387_1616_, _358_1161_, _355_399_, _399_1428_,
    _402_1718_, _372_1243_, _396_1504_, _405_1717_, _409_1670_, _378_1597_,
    _390_1603_, _361_940_, _367_1585_, _407_1657_  );
  input  _77_9_, _87_10_, _169_22_, _238_31_, _2897_49_, _68_8_,
    _128_16_, _226_29_, _294_39_, _326_44_, _58_7_, _190_24_, _264_35_,
    _283_38_, _250_33_, _329_45_, _213_26_, _257_34_, _20_2_, _223_28_,
    _159_21_, _232_30_, _41_4_, _124_14_, _13_1_, _50_6_, _222_27_,
    _97_11_, _125_15_, _322_43_, _244_32_, _274_37_, _317_42_, _1_0_,
    _33_3_, _270_36_, _200_25_, _343_47_, _330_46_, _1698_48_, _132_17_,
    _45_5_, _116_13_, _143_19_, _303_40_, _311_41_, _107_12_, _137_18_,
    _150_20_, _179_23_;
  output _381_1626_, _351_1247_, _353_405_, _375_1624_, _393_1605_,
    _364_1484_, _369_1321_, _384_1553_, _387_1616_, _358_1161_, _355_399_,
    _399_1428_, _402_1718_, _372_1243_, _396_1504_, _405_1717_, _409_1670_,
    _378_1597_, _390_1603_, _361_940_, _367_1585_, _407_1657_;
  wire new_n73, new_n74, new_n75, new_n76, new_n77, new_n78, new_n79,
    new_n80, new_n81, new_n82, new_n83, new_n84, new_n85, new_n86, new_n87,
    new_n88, new_n89, new_n90, new_n91, new_n92, new_n93, new_n94, new_n95,
    new_n96, new_n97, new_n98, new_n99, new_n100, new_n101, new_n102,
    new_n103, new_n104, new_n105, new_n106, new_n107, new_n108, new_n109,
    new_n110, new_n111, new_n112, new_n113, new_n114, new_n115, new_n116,
    new_n117, new_n118, new_n119, new_n120, new_n121, new_n122, new_n123,
    new_n124, new_n125, new_n126, new_n127, new_n128, new_n129, new_n130,
    new_n131, new_n132, new_n133, new_n134, new_n135, new_n136, new_n137,
    new_n138, new_n139, new_n140, new_n141, new_n142, new_n143, new_n144,
    new_n145, new_n146, new_n147, new_n148, new_n149, new_n150, new_n151,
    new_n152, new_n153, new_n154, new_n155, new_n156, new_n157, new_n158,
    new_n159, new_n160, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115;
  assign new_n73 = ~_41_4_ & ~_13_1_;
  assign new_n74 = _20_2_ & new_n73;
  assign new_n75 = _1_0_ & new_n74;
  assign new_n76 = _20_2_ & _13_1_;
  assign new_n77 = ~_1_0_ & new_n76;
  assign new_n78 = ~_77_9_ & new_n77;
  assign new_n79 = _20_2_ & ~_1_0_;
  assign new_n80 = _20_2_ & _33_3_;
  assign new_n81 = _1_0_ & new_n80;
  assign new_n82 = _13_1_ & _1_0_;
  assign new_n83 = ~new_n81 & ~new_n82;
  assign new_n84 = ~new_n77 & new_n83;
  assign new_n85 = ~new_n79 & new_n84;
  assign new_n86 = _77_9_ & new_n85;
  assign new_n87 = ~_20_2_ & _33_3_;
  assign new_n88 = _87_10_ & new_n87;
  assign new_n89 = ~_20_2_ & ~new_n87;
  assign new_n90 = _58_7_ & new_n89;
  assign new_n91 = _77_9_ & _20_2_;
  assign new_n92 = ~new_n88 & ~new_n90;
  assign new_n93 = ~new_n91 & new_n92;
  assign new_n94 = ~new_n83 & ~new_n93;
  assign new_n95 = ~new_n78 & ~new_n86;
  assign new_n96 = ~new_n94 & new_n95;
  assign new_n97 = ~_41_4_ & ~_45_5_;
  assign new_n98 = ~_1_0_ & ~new_n97;
  assign new_n99 = _41_4_ & _33_3_;
  assign new_n100 = _13_1_ & ~new_n99;
  assign new_n101 = _1_0_ & new_n100;
  assign new_n102 = _274_37_ & new_n98;
  assign new_n103 = ~new_n101 & new_n102;
  assign new_n104 = ~_33_3_ & ~_1698_48_;
  assign new_n105 = _232_30_ & new_n104;
  assign new_n106 = ~_33_3_ & ~new_n104;
  assign new_n107 = _238_31_ & new_n106;
  assign new_n108 = _33_3_ & _107_12_;
  assign new_n109 = ~new_n105 & ~new_n107;
  assign new_n110 = ~new_n108 & new_n109;
  assign new_n111 = new_n101 & ~new_n110;
  assign new_n112 = _244_32_ & ~new_n98;
  assign new_n113 = ~new_n101 & new_n112;
  assign new_n114 = ~new_n103 & ~new_n111;
  assign new_n115 = ~new_n113 & new_n114;
  assign new_n116 = new_n96 & ~new_n115;
  assign new_n117 = _200_25_ & new_n116;
  assign new_n118 = new_n96 & new_n115;
  assign new_n119 = _190_24_ & new_n118;
  assign new_n120 = new_n96 & ~new_n117;
  assign new_n121 = ~new_n119 & new_n120;
  assign new_n122 = ~new_n96 & new_n115;
  assign new_n123 = _179_23_ & new_n122;
  assign new_n124 = ~new_n96 & ~new_n115;
  assign new_n125 = _169_22_ & new_n124;
  assign new_n126 = ~new_n123 & ~new_n125;
  assign new_n127 = ~new_n121 & new_n126;
  assign new_n128 = ~_58_7_ & new_n77;
  assign new_n129 = _58_7_ & new_n85;
  assign new_n130 = _68_8_ & new_n87;
  assign new_n131 = _159_21_ & new_n89;
  assign new_n132 = ~_68_8_ & _58_7_;
  assign new_n133 = _68_8_ & ~_58_7_;
  assign new_n134 = ~new_n132 & ~new_n133;
  assign new_n135 = _20_2_ & new_n134;
  assign new_n136 = ~new_n130 & ~new_n131;
  assign new_n137 = ~new_n135 & new_n136;
  assign new_n138 = ~new_n83 & ~new_n137;
  assign new_n139 = ~new_n128 & ~new_n129;
  assign new_n140 = ~new_n138 & new_n139;
  assign new_n141 = _223_28_ & new_n104;
  assign new_n142 = _226_29_ & new_n106;
  assign new_n143 = _87_10_ & _33_3_;
  assign new_n144 = ~new_n141 & ~new_n142;
  assign new_n145 = ~new_n143 & new_n144;
  assign new_n146 = new_n101 & ~new_n145;
  assign new_n147 = _232_30_ & ~new_n98;
  assign new_n148 = ~new_n101 & new_n147;
  assign new_n149 = ~new_n103 & ~new_n146;
  assign new_n150 = ~new_n148 & new_n149;
  assign new_n151 = new_n140 & ~new_n150;
  assign new_n152 = _200_25_ & new_n151;
  assign new_n153 = new_n140 & new_n150;
  assign new_n154 = _190_24_ & new_n153;
  assign new_n155 = new_n140 & ~new_n152;
  assign new_n156 = ~new_n154 & new_n155;
  assign new_n157 = ~new_n140 & new_n150;
  assign new_n158 = _179_23_ & new_n157;
  assign new_n159 = ~new_n140 & ~new_n150;
  assign new_n160 = _169_22_ & new_n159;
  assign new_n161 = ~new_n158 & ~new_n160;
  assign new_n162 = ~new_n156 & new_n161;
  assign new_n163 = ~_68_8_ & new_n77;
  assign new_n164 = _68_8_ & new_n85;
  assign new_n165 = _77_9_ & new_n87;
  assign new_n166 = _50_6_ & new_n89;
  assign new_n167 = ~_68_8_ & _20_2_;
  assign new_n168 = ~new_n165 & ~new_n166;
  assign new_n169 = ~new_n167 & new_n168;
  assign new_n170 = ~new_n83 & ~new_n169;
  assign new_n171 = ~new_n163 & ~new_n164;
  assign new_n172 = ~new_n170 & new_n171;
  assign new_n173 = _226_29_ & new_n104;
  assign new_n174 = _232_30_ & new_n106;
  assign new_n175 = _97_11_ & _33_3_;
  assign new_n176 = ~new_n173 & ~new_n174;
  assign new_n177 = ~new_n175 & new_n176;
  assign new_n178 = new_n101 & ~new_n177;
  assign new_n179 = _238_31_ & ~new_n98;
  assign new_n180 = ~new_n101 & new_n179;
  assign new_n181 = ~new_n103 & ~new_n178;
  assign new_n182 = ~new_n180 & new_n181;
  assign new_n183 = new_n172 & ~new_n182;
  assign new_n184 = _200_25_ & new_n183;
  assign new_n185 = new_n172 & new_n182;
  assign new_n186 = _190_24_ & new_n185;
  assign new_n187 = new_n172 & ~new_n184;
  assign new_n188 = ~new_n186 & new_n187;
  assign new_n189 = ~new_n172 & new_n182;
  assign new_n190 = _179_23_ & new_n189;
  assign new_n191 = ~new_n172 & ~new_n182;
  assign new_n192 = _169_22_ & new_n191;
  assign new_n193 = ~new_n190 & ~new_n192;
  assign new_n194 = ~new_n188 & new_n193;
  assign new_n195 = ~_50_6_ & new_n77;
  assign new_n196 = _50_6_ & new_n85;
  assign new_n197 = _58_7_ & new_n87;
  assign new_n198 = _150_20_ & new_n89;
  assign new_n199 = ~_68_8_ & ~_58_7_;
  assign new_n200 = ~_50_6_ & new_n199;
  assign new_n201 = _20_2_ & ~new_n200;
  assign new_n202 = ~new_n197 & ~new_n198;
  assign new_n203 = ~new_n201 & new_n202;
  assign new_n204 = ~new_n83 & ~new_n203;
  assign new_n205 = ~new_n195 & ~new_n196;
  assign new_n206 = ~new_n204 & new_n205;
  assign new_n207 = _222_27_ & new_n104;
  assign new_n208 = _223_28_ & new_n106;
  assign new_n209 = _77_9_ & _33_3_;
  assign new_n210 = ~new_n207 & ~new_n208;
  assign new_n211 = ~new_n209 & new_n210;
  assign new_n212 = new_n101 & ~new_n211;
  assign new_n213 = _226_29_ & ~new_n98;
  assign new_n214 = ~new_n101 & new_n213;
  assign new_n215 = ~new_n103 & ~new_n212;
  assign new_n216 = ~new_n214 & new_n215;
  assign new_n217 = new_n206 & ~new_n216;
  assign new_n218 = _200_25_ & new_n217;
  assign new_n219 = new_n206 & new_n216;
  assign new_n220 = _190_24_ & new_n219;
  assign new_n221 = new_n206 & ~new_n218;
  assign new_n222 = ~new_n220 & new_n221;
  assign new_n223 = ~new_n206 & new_n216;
  assign new_n224 = _179_23_ & new_n223;
  assign new_n225 = ~new_n206 & ~new_n216;
  assign new_n226 = _169_22_ & new_n225;
  assign new_n227 = ~new_n224 & ~new_n226;
  assign new_n228 = ~new_n222 & new_n227;
  assign new_n229 = new_n127 & new_n162;
  assign new_n230 = new_n194 & new_n229;
  assign new_n231 = new_n228 & new_n230;
  assign new_n232 = ~_20_2_ & _13_1_;
  assign new_n233 = ~_1_0_ & new_n232;
  assign new_n234 = _213_26_ & _343_47_;
  assign new_n235 = new_n233 & new_n234;
  assign new_n236 = ~_87_10_ & new_n77;
  assign new_n237 = ~_1_0_ & _33_3_;
  assign new_n238 = new_n84 & ~new_n237;
  assign new_n239 = _87_10_ & new_n238;
  assign new_n240 = _97_11_ & new_n87;
  assign new_n241 = _68_8_ & new_n89;
  assign new_n242 = ~_97_11_ & ~_107_12_;
  assign new_n243 = ~_87_10_ & new_n242;
  assign new_n244 = _20_2_ & ~new_n243;
  assign new_n245 = ~new_n240 & ~new_n241;
  assign new_n246 = ~new_n244 & new_n245;
  assign new_n247 = ~new_n83 & ~new_n246;
  assign new_n248 = ~new_n236 & ~new_n239;
  assign new_n249 = ~new_n247 & new_n248;
  assign new_n250 = ~_1_0_ & _45_5_;
  assign new_n251 = _274_37_ & new_n250;
  assign new_n252 = ~new_n101 & new_n251;
  assign new_n253 = _238_31_ & new_n104;
  assign new_n254 = _244_32_ & new_n106;
  assign new_n255 = _33_3_ & _116_13_;
  assign new_n256 = ~new_n253 & ~new_n254;
  assign new_n257 = ~new_n255 & new_n256;
  assign new_n258 = new_n101 & ~new_n257;
  assign new_n259 = _250_33_ & ~new_n250;
  assign new_n260 = ~new_n101 & new_n259;
  assign new_n261 = ~new_n252 & ~new_n258;
  assign new_n262 = ~new_n260 & new_n261;
  assign new_n263 = new_n249 & ~new_n262;
  assign new_n264 = _200_25_ & new_n263;
  assign new_n265 = new_n249 & new_n262;
  assign new_n266 = _190_24_ & new_n265;
  assign new_n267 = new_n249 & ~new_n264;
  assign new_n268 = ~new_n266 & new_n267;
  assign new_n269 = ~new_n249 & new_n262;
  assign new_n270 = _179_23_ & new_n269;
  assign new_n271 = ~new_n249 & ~new_n262;
  assign new_n272 = _169_22_ & new_n271;
  assign new_n273 = ~new_n270 & ~new_n272;
  assign new_n274 = ~new_n268 & new_n273;
  assign new_n275 = ~_97_11_ & new_n77;
  assign new_n276 = _97_11_ & new_n238;
  assign new_n277 = _107_12_ & new_n87;
  assign new_n278 = _77_9_ & new_n89;
  assign new_n279 = _97_11_ & ~_107_12_;
  assign new_n280 = ~_97_11_ & _107_12_;
  assign new_n281 = ~new_n279 & ~new_n280;
  assign new_n282 = _20_2_ & new_n281;
  assign new_n283 = ~new_n277 & ~new_n278;
  assign new_n284 = ~new_n282 & new_n283;
  assign new_n285 = ~new_n83 & ~new_n284;
  assign new_n286 = ~new_n275 & ~new_n276;
  assign new_n287 = ~new_n285 & new_n286;
  assign new_n288 = ~_41_4_ & _45_5_;
  assign new_n289 = ~_1_0_ & new_n288;
  assign new_n290 = _274_37_ & new_n289;
  assign new_n291 = ~new_n101 & new_n290;
  assign new_n292 = _244_32_ & new_n104;
  assign new_n293 = _250_33_ & new_n106;
  assign new_n294 = _283_38_ & _33_3_;
  assign new_n295 = ~new_n292 & ~new_n293;
  assign new_n296 = ~new_n294 & new_n295;
  assign new_n297 = new_n101 & ~new_n296;
  assign new_n298 = _257_34_ & ~new_n289;
  assign new_n299 = ~new_n101 & new_n298;
  assign new_n300 = ~new_n291 & ~new_n297;
  assign new_n301 = ~new_n299 & new_n300;
  assign new_n302 = new_n287 & ~new_n301;
  assign new_n303 = _200_25_ & new_n302;
  assign new_n304 = new_n287 & new_n301;
  assign new_n305 = _190_24_ & new_n304;
  assign new_n306 = new_n287 & ~new_n303;
  assign new_n307 = ~new_n305 & new_n306;
  assign new_n308 = ~new_n287 & new_n301;
  assign new_n309 = _179_23_ & new_n308;
  assign new_n310 = ~new_n287 & ~new_n301;
  assign new_n311 = _169_22_ & new_n310;
  assign new_n312 = ~new_n309 & ~new_n311;
  assign new_n313 = ~new_n307 & new_n312;
  assign new_n314 = ~_107_12_ & new_n77;
  assign new_n315 = _107_12_ & new_n238;
  assign new_n316 = _116_13_ & new_n87;
  assign new_n317 = _87_10_ & new_n89;
  assign new_n318 = _20_2_ & ~_107_12_;
  assign new_n319 = ~new_n316 & ~new_n317;
  assign new_n320 = ~new_n318 & new_n319;
  assign new_n321 = ~new_n83 & ~new_n320;
  assign new_n322 = ~new_n314 & ~new_n315;
  assign new_n323 = ~new_n321 & new_n322;
  assign new_n324 = _250_33_ & new_n104;
  assign new_n325 = _257_34_ & new_n106;
  assign new_n326 = _294_39_ & _33_3_;
  assign new_n327 = ~new_n324 & ~new_n325;
  assign new_n328 = ~new_n326 & new_n327;
  assign new_n329 = new_n101 & ~new_n328;
  assign new_n330 = _264_35_ & ~new_n289;
  assign new_n331 = ~new_n101 & new_n330;
  assign new_n332 = ~new_n291 & ~new_n329;
  assign new_n333 = ~new_n331 & new_n332;
  assign new_n334 = new_n323 & ~new_n333;
  assign new_n335 = _200_25_ & new_n334;
  assign new_n336 = new_n323 & new_n333;
  assign new_n337 = _190_24_ & new_n336;
  assign new_n338 = new_n323 & ~new_n335;
  assign new_n339 = ~new_n337 & new_n338;
  assign new_n340 = ~new_n323 & new_n333;
  assign new_n341 = _179_23_ & new_n340;
  assign new_n342 = ~new_n323 & ~new_n333;
  assign new_n343 = _169_22_ & new_n342;
  assign new_n344 = ~new_n341 & ~new_n343;
  assign new_n345 = ~new_n339 & new_n344;
  assign new_n346 = ~_116_13_ & new_n77;
  assign new_n347 = _116_13_ & new_n238;
  assign new_n348 = _283_38_ & new_n87;
  assign new_n349 = _97_11_ & new_n89;
  assign new_n350 = _20_2_ & _116_13_;
  assign new_n351 = ~new_n348 & ~new_n349;
  assign new_n352 = ~new_n350 & new_n351;
  assign new_n353 = ~new_n83 & ~new_n352;
  assign new_n354 = ~new_n346 & ~new_n347;
  assign new_n355 = ~new_n353 & new_n354;
  assign new_n356 = _257_34_ & new_n104;
  assign new_n357 = _264_35_ & new_n106;
  assign new_n358 = _33_3_ & _303_40_;
  assign new_n359 = ~new_n356 & ~new_n357;
  assign new_n360 = ~new_n358 & new_n359;
  assign new_n361 = new_n101 & ~new_n360;
  assign new_n362 = _270_36_ & ~new_n289;
  assign new_n363 = ~new_n101 & new_n362;
  assign new_n364 = ~new_n291 & ~new_n361;
  assign new_n365 = ~new_n363 & new_n364;
  assign new_n366 = ~new_n355 & new_n365;
  assign new_n367 = _179_23_ & new_n366;
  assign new_n368 = ~new_n355 & ~new_n365;
  assign new_n369 = _169_22_ & new_n368;
  assign new_n370 = ~new_n367 & ~new_n369;
  assign new_n371 = new_n274 & new_n313;
  assign new_n372 = new_n345 & new_n371;
  assign new_n373 = ~new_n370 & new_n372;
  assign new_n374 = new_n274 & ~new_n312;
  assign new_n375 = new_n313 & ~new_n344;
  assign new_n376 = new_n274 & new_n375;
  assign new_n377 = ~new_n373 & ~new_n374;
  assign new_n378 = ~new_n376 & new_n377;
  assign new_n379 = new_n273 & new_n378;
  assign new_n380 = ~new_n235 & ~new_n379;
  assign new_n381 = new_n231 & new_n380;
  assign new_n382 = new_n162 & new_n228;
  assign new_n383 = new_n194 & new_n382;
  assign new_n384 = ~new_n126 & new_n383;
  assign new_n385 = ~new_n161 & new_n228;
  assign new_n386 = new_n162 & ~new_n193;
  assign new_n387 = new_n228 & new_n386;
  assign new_n388 = ~new_n384 & ~new_n385;
  assign new_n389 = ~new_n387 & new_n388;
  assign new_n390 = new_n227 & new_n389;
  assign new_n391 = ~new_n381 & new_n390;
  assign new_n392 = new_n355 & ~new_n365;
  assign new_n393 = _200_25_ & new_n392;
  assign new_n394 = new_n355 & new_n365;
  assign new_n395 = _190_24_ & new_n394;
  assign new_n396 = new_n355 & ~new_n393;
  assign new_n397 = ~new_n395 & new_n396;
  assign new_n398 = new_n370 & ~new_n397;
  assign new_n399 = new_n313 & new_n398;
  assign new_n400 = new_n345 & new_n399;
  assign new_n401 = new_n274 & new_n400;
  assign new_n402 = ~new_n235 & new_n401;
  assign new_n403 = _179_23_ & new_n365;
  assign new_n404 = new_n301 & new_n403;
  assign new_n405 = new_n333 & new_n404;
  assign new_n406 = new_n262 & new_n405;
  assign new_n407 = ~_179_23_ & ~new_n365;
  assign new_n408 = ~new_n301 & new_n407;
  assign new_n409 = ~new_n333 & new_n408;
  assign new_n410 = ~new_n262 & new_n409;
  assign new_n411 = ~new_n406 & ~new_n410;
  assign new_n412 = new_n235 & ~new_n411;
  assign new_n413 = ~new_n402 & ~new_n412;
  assign new_n414 = new_n231 & ~new_n413;
  assign new_n415 = new_n391 & new_n414;
  assign new_n416 = _330_46_ & new_n415;
  assign new_n417 = new_n391 & ~new_n416;
  assign new_n418 = ~new_n96 & new_n235;
  assign new_n419 = new_n127 & ~new_n418;
  assign new_n420 = ~new_n127 & new_n418;
  assign new_n421 = ~new_n419 & ~new_n420;
  assign new_n422 = ~new_n413 & ~new_n421;
  assign new_n423 = _330_46_ & new_n422;
  assign new_n424 = ~new_n172 & new_n235;
  assign new_n425 = new_n194 & ~new_n424;
  assign new_n426 = ~new_n194 & new_n424;
  assign new_n427 = ~new_n425 & ~new_n426;
  assign new_n428 = new_n380 & ~new_n421;
  assign new_n429 = ~new_n126 & ~new_n235;
  assign new_n430 = ~new_n428 & ~new_n429;
  assign new_n431 = new_n427 & ~new_n430;
  assign new_n432 = ~new_n427 & new_n430;
  assign new_n433 = ~new_n431 & ~new_n432;
  assign new_n434 = ~new_n423 & ~new_n433;
  assign new_n435 = new_n423 & new_n433;
  assign new_n436 = ~new_n434 & ~new_n435;
  assign new_n437 = ~new_n417 & new_n436;
  assign new_n438 = new_n417 & ~new_n436;
  assign new_n439 = ~new_n437 & ~new_n438;
  assign new_n440 = new_n75 & new_n439;
  assign new_n441 = ~_20_2_ & _45_5_;
  assign new_n442 = _13_1_ & new_n441;
  assign new_n443 = _1_0_ & ~new_n442;
  assign new_n444 = ~new_n75 & new_n443;
  assign new_n445 = ~_13_1_ & ~_33_3_;
  assign new_n446 = new_n427 & new_n445;
  assign new_n447 = ~_169_22_ & _20_2_;
  assign new_n448 = _13_1_ & ~new_n447;
  assign new_n449 = _1_0_ & new_n448;
  assign new_n450 = ~new_n445 & ~new_n449;
  assign new_n451 = ~_68_8_ & new_n450;
  assign new_n452 = _20_2_ & _179_23_;
  assign new_n453 = _20_2_ & _200_25_;
  assign new_n454 = ~new_n452 & new_n453;
  assign new_n455 = ~_190_24_ & _20_2_;
  assign new_n456 = new_n454 & ~new_n455;
  assign new_n457 = _97_11_ & new_n456;
  assign new_n458 = ~_200_25_ & new_n452;
  assign new_n459 = new_n455 & new_n458;
  assign new_n460 = _107_12_ & new_n459;
  assign new_n461 = new_n454 & new_n455;
  assign new_n462 = _77_9_ & new_n461;
  assign new_n463 = ~new_n452 & ~new_n453;
  assign new_n464 = ~new_n455 & new_n463;
  assign new_n465 = _87_10_ & new_n464;
  assign new_n466 = new_n455 & new_n463;
  assign new_n467 = _303_40_ & new_n466;
  assign new_n468 = _200_25_ & new_n452;
  assign new_n469 = ~new_n455 & new_n468;
  assign new_n470 = _294_39_ & new_n469;
  assign new_n471 = new_n455 & new_n468;
  assign new_n472 = _116_13_ & new_n471;
  assign new_n473 = ~new_n455 & new_n458;
  assign new_n474 = _283_38_ & new_n473;
  assign new_n475 = ~new_n457 & ~new_n460;
  assign new_n476 = ~new_n462 & new_n475;
  assign new_n477 = ~new_n465 & new_n476;
  assign new_n478 = ~new_n467 & new_n477;
  assign new_n479 = ~new_n470 & new_n478;
  assign new_n480 = ~new_n472 & new_n479;
  assign new_n481 = ~new_n474 & new_n480;
  assign new_n482 = _33_3_ & new_n481;
  assign new_n483 = _159_21_ & new_n456;
  assign new_n484 = _150_20_ & new_n459;
  assign new_n485 = _58_7_ & new_n461;
  assign new_n486 = _50_6_ & new_n464;
  assign new_n487 = _128_16_ & new_n466;
  assign new_n488 = _132_17_ & new_n469;
  assign new_n489 = _143_19_ & new_n471;
  assign new_n490 = _137_18_ & new_n473;
  assign new_n491 = ~new_n483 & ~new_n484;
  assign new_n492 = ~new_n485 & new_n491;
  assign new_n493 = ~new_n486 & new_n492;
  assign new_n494 = ~new_n487 & new_n493;
  assign new_n495 = ~new_n488 & new_n494;
  assign new_n496 = ~new_n489 & new_n495;
  assign new_n497 = ~new_n490 & new_n496;
  assign new_n498 = ~_33_3_ & new_n497;
  assign new_n499 = ~new_n482 & ~new_n498;
  assign new_n500 = new_n449 & ~new_n499;
  assign new_n501 = ~new_n446 & ~new_n451;
  assign new_n502 = ~new_n500 & new_n501;
  assign new_n503 = new_n444 & new_n502;
  assign new_n504 = ~new_n436 & ~new_n443;
  assign new_n505 = ~new_n440 & ~new_n503;
  assign _381_1626_ = new_n504 | ~new_n505;
  assign new_n507 = _116_13_ & ~_107_12_;
  assign new_n508 = ~_116_13_ & _107_12_;
  assign new_n509 = ~new_n507 & ~new_n508;
  assign new_n510 = ~_87_10_ & _97_11_;
  assign new_n511 = _87_10_ & ~_97_11_;
  assign new_n512 = ~new_n510 & ~new_n511;
  assign new_n513 = new_n509 & ~new_n512;
  assign new_n514 = ~new_n509 & new_n512;
  assign new_n515 = ~new_n513 & ~new_n514;
  assign new_n516 = _77_9_ & ~_68_8_;
  assign new_n517 = ~_77_9_ & _68_8_;
  assign new_n518 = ~new_n516 & ~new_n517;
  assign new_n519 = _58_7_ & _50_6_;
  assign new_n520 = ~_58_7_ & ~_50_6_;
  assign new_n521 = ~new_n519 & ~new_n520;
  assign new_n522 = new_n518 & ~new_n521;
  assign new_n523 = ~new_n518 & new_n521;
  assign new_n524 = ~new_n522 & ~new_n523;
  assign new_n525 = new_n515 & ~new_n524;
  assign new_n526 = ~new_n515 & new_n524;
  assign _351_1247_ = new_n525 | new_n526;
  assign _353_405_ = ~_77_9_ & new_n200;
  assign new_n529 = ~new_n421 & ~new_n427;
  assign new_n530 = ~new_n413 & new_n529;
  assign new_n531 = _330_46_ & new_n530;
  assign new_n532 = _213_26_ & new_n233;
  assign new_n533 = ~new_n140 & new_n532;
  assign new_n534 = new_n162 & ~new_n533;
  assign new_n535 = ~new_n162 & new_n533;
  assign new_n536 = ~new_n534 & ~new_n535;
  assign new_n537 = ~new_n427 & new_n429;
  assign new_n538 = ~new_n427 & new_n428;
  assign new_n539 = ~new_n193 & ~new_n235;
  assign new_n540 = ~new_n537 & ~new_n538;
  assign new_n541 = ~new_n539 & new_n540;
  assign new_n542 = new_n536 & ~new_n541;
  assign new_n543 = ~new_n536 & new_n541;
  assign new_n544 = ~new_n542 & ~new_n543;
  assign new_n545 = ~new_n531 & ~new_n544;
  assign new_n546 = new_n531 & new_n544;
  assign new_n547 = ~new_n545 & ~new_n546;
  assign new_n548 = ~new_n421 & ~new_n536;
  assign new_n549 = ~new_n427 & new_n548;
  assign new_n550 = ~new_n413 & new_n549;
  assign new_n551 = _330_46_ & new_n550;
  assign new_n552 = ~new_n206 & new_n532;
  assign new_n553 = new_n228 & ~new_n552;
  assign new_n554 = ~new_n228 & new_n552;
  assign new_n555 = ~new_n553 & ~new_n554;
  assign new_n556 = new_n380 & ~new_n427;
  assign new_n557 = ~new_n421 & new_n556;
  assign new_n558 = ~new_n536 & new_n557;
  assign new_n559 = ~new_n536 & new_n539;
  assign new_n560 = ~new_n536 & new_n537;
  assign new_n561 = ~new_n161 & ~new_n532;
  assign new_n562 = ~new_n558 & ~new_n559;
  assign new_n563 = ~new_n560 & new_n562;
  assign new_n564 = ~new_n561 & new_n563;
  assign new_n565 = new_n555 & ~new_n564;
  assign new_n566 = ~new_n555 & new_n564;
  assign new_n567 = ~new_n565 & ~new_n566;
  assign new_n568 = ~new_n551 & ~new_n567;
  assign new_n569 = new_n551 & new_n567;
  assign new_n570 = ~new_n568 & ~new_n569;
  assign new_n571 = new_n417 & ~new_n547;
  assign new_n572 = ~new_n570 & new_n571;
  assign new_n573 = ~new_n436 & new_n572;
  assign new_n574 = ~new_n417 & ~new_n570;
  assign new_n575 = ~new_n573 & ~new_n574;
  assign new_n576 = new_n75 & ~new_n575;
  assign new_n577 = new_n445 & new_n555;
  assign new_n578 = ~_50_6_ & new_n450;
  assign new_n579 = ~_41_4_ & _33_3_;
  assign new_n580 = _77_9_ & new_n456;
  assign new_n581 = _87_10_ & new_n459;
  assign new_n582 = _68_8_ & new_n464;
  assign new_n583 = _283_38_ & new_n466;
  assign new_n584 = _116_13_ & new_n469;
  assign new_n585 = _97_11_ & new_n471;
  assign new_n586 = _107_12_ & new_n473;
  assign new_n587 = ~new_n580 & ~new_n581;
  assign new_n588 = ~new_n485 & new_n587;
  assign new_n589 = ~new_n582 & new_n588;
  assign new_n590 = ~new_n583 & new_n589;
  assign new_n591 = ~new_n584 & new_n590;
  assign new_n592 = ~new_n585 & new_n591;
  assign new_n593 = ~new_n586 & new_n592;
  assign new_n594 = new_n579 & new_n593;
  assign new_n595 = ~_41_4_ & ~_33_3_;
  assign new_n596 = ~new_n579 & ~new_n595;
  assign new_n597 = ~_50_6_ & new_n596;
  assign new_n598 = _143_19_ & new_n456;
  assign new_n599 = _137_18_ & new_n459;
  assign new_n600 = _159_21_ & new_n461;
  assign new_n601 = _150_20_ & new_n464;
  assign new_n602 = _124_14_ & new_n466;
  assign new_n603 = _125_15_ & new_n469;
  assign new_n604 = _132_17_ & new_n471;
  assign new_n605 = _128_16_ & new_n473;
  assign new_n606 = ~new_n598 & ~new_n599;
  assign new_n607 = ~new_n600 & new_n606;
  assign new_n608 = ~new_n601 & new_n607;
  assign new_n609 = ~new_n602 & new_n608;
  assign new_n610 = ~new_n603 & new_n609;
  assign new_n611 = ~new_n604 & new_n610;
  assign new_n612 = ~new_n605 & new_n611;
  assign new_n613 = new_n595 & new_n612;
  assign new_n614 = ~new_n594 & ~new_n597;
  assign new_n615 = ~new_n613 & new_n614;
  assign new_n616 = new_n449 & ~new_n615;
  assign new_n617 = ~new_n577 & ~new_n578;
  assign new_n618 = ~new_n616 & new_n617;
  assign new_n619 = new_n444 & new_n618;
  assign new_n620 = ~new_n443 & ~new_n570;
  assign new_n621 = ~new_n576 & ~new_n619;
  assign _375_1624_ = new_n620 | ~new_n621;
  assign new_n623 = ~new_n380 & ~new_n413;
  assign new_n624 = _330_46_ & new_n623;
  assign new_n625 = ~new_n380 & ~new_n624;
  assign new_n626 = new_n235 & ~new_n355;
  assign new_n627 = new_n398 & ~new_n626;
  assign new_n628 = ~new_n398 & new_n626;
  assign new_n629 = ~new_n627 & ~new_n628;
  assign new_n630 = _330_46_ & ~new_n629;
  assign new_n631 = new_n235 & ~new_n323;
  assign new_n632 = new_n345 & ~new_n631;
  assign new_n633 = ~new_n345 & new_n631;
  assign new_n634 = ~new_n632 & ~new_n633;
  assign new_n635 = ~new_n235 & ~new_n370;
  assign new_n636 = new_n634 & new_n635;
  assign new_n637 = ~new_n634 & ~new_n635;
  assign new_n638 = ~new_n636 & ~new_n637;
  assign new_n639 = ~new_n630 & ~new_n638;
  assign new_n640 = new_n630 & new_n638;
  assign new_n641 = ~new_n639 & ~new_n640;
  assign new_n642 = ~new_n625 & new_n641;
  assign new_n643 = new_n625 & ~new_n641;
  assign new_n644 = ~new_n642 & ~new_n643;
  assign new_n645 = new_n75 & new_n644;
  assign new_n646 = ~_20_2_ & ~_33_3_;
  assign new_n647 = ~_13_1_ & new_n646;
  assign new_n648 = new_n634 & new_n647;
  assign new_n649 = ~new_n449 & ~new_n647;
  assign new_n650 = _20_2_ & ~_13_1_;
  assign new_n651 = _1_0_ & new_n650;
  assign new_n652 = ~_33_3_ & new_n651;
  assign new_n653 = ~_116_13_ & new_n243;
  assign new_n654 = new_n652 & ~new_n653;
  assign new_n655 = _33_3_ & new_n651;
  assign new_n656 = ~new_n652 & ~new_n655;
  assign new_n657 = ~_107_12_ & new_n656;
  assign new_n658 = _77_9_ & _68_8_;
  assign new_n659 = _58_7_ & ~new_n658;
  assign new_n660 = ~_50_6_ & new_n659;
  assign new_n661 = new_n653 & new_n660;
  assign new_n662 = ~_45_5_ & new_n661;
  assign new_n663 = _238_31_ & ~_244_32_;
  assign new_n664 = ~_238_31_ & _244_32_;
  assign new_n665 = ~new_n663 & ~new_n664;
  assign new_n666 = _226_29_ & ~_232_30_;
  assign new_n667 = ~_226_29_ & _232_30_;
  assign new_n668 = ~new_n666 & ~new_n667;
  assign new_n669 = new_n665 & ~new_n668;
  assign new_n670 = ~new_n665 & new_n668;
  assign new_n671 = ~new_n669 & ~new_n670;
  assign new_n672 = _45_5_ & new_n671;
  assign new_n673 = ~new_n662 & ~new_n672;
  assign new_n674 = new_n655 & new_n673;
  assign new_n675 = ~new_n654 & ~new_n657;
  assign new_n676 = ~new_n674 & new_n675;
  assign new_n677 = new_n649 & ~new_n676;
  assign new_n678 = _294_39_ & new_n456;
  assign new_n679 = _303_40_ & new_n459;
  assign new_n680 = _116_13_ & new_n461;
  assign new_n681 = _283_38_ & new_n464;
  assign new_n682 = _326_44_ & new_n466;
  assign new_n683 = _322_43_ & new_n469;
  assign new_n684 = _311_41_ & new_n471;
  assign new_n685 = _317_42_ & new_n473;
  assign new_n686 = ~new_n678 & ~new_n679;
  assign new_n687 = ~new_n680 & new_n686;
  assign new_n688 = ~new_n681 & new_n687;
  assign new_n689 = ~new_n682 & new_n688;
  assign new_n690 = ~new_n683 & new_n689;
  assign new_n691 = ~new_n684 & new_n690;
  assign new_n692 = ~new_n685 & new_n691;
  assign new_n693 = _33_3_ & new_n692;
  assign new_n694 = _68_8_ & new_n459;
  assign new_n695 = _97_11_ & new_n461;
  assign new_n696 = _150_20_ & new_n466;
  assign new_n697 = _159_21_ & new_n469;
  assign new_n698 = _58_7_ & new_n471;
  assign new_n699 = _50_6_ & new_n473;
  assign new_n700 = ~new_n580 & ~new_n694;
  assign new_n701 = ~new_n695 & new_n700;
  assign new_n702 = ~new_n465 & new_n701;
  assign new_n703 = ~new_n696 & new_n702;
  assign new_n704 = ~new_n697 & new_n703;
  assign new_n705 = ~new_n698 & new_n704;
  assign new_n706 = ~new_n699 & new_n705;
  assign new_n707 = ~_33_3_ & new_n706;
  assign new_n708 = ~new_n693 & ~new_n707;
  assign new_n709 = new_n449 & ~new_n708;
  assign new_n710 = ~new_n648 & ~new_n677;
  assign new_n711 = ~new_n709 & new_n710;
  assign new_n712 = new_n444 & new_n711;
  assign new_n713 = ~new_n443 & ~new_n641;
  assign new_n714 = ~new_n645 & ~new_n712;
  assign _393_1605_ = new_n713 | ~new_n714;
  assign new_n716 = ~_1_0_ & ~new_n625;
  assign new_n717 = _1_0_ & ~new_n75;
  assign new_n718 = new_n653 & new_n717;
  assign new_n719 = _50_6_ & ~new_n199;
  assign new_n720 = new_n75 & new_n719;
  assign new_n721 = ~new_n716 & ~new_n718;
  assign _364_1484_ = new_n720 | ~new_n721;
  assign new_n723 = new_n231 & ~new_n379;
  assign _369_1321_ = ~new_n390 | new_n723;
  assign new_n725 = _330_46_ & ~new_n413;
  assign new_n726 = new_n380 & new_n421;
  assign new_n727 = ~new_n380 & ~new_n421;
  assign new_n728 = ~new_n726 & ~new_n727;
  assign new_n729 = ~new_n725 & ~new_n728;
  assign new_n730 = new_n725 & new_n728;
  assign new_n731 = ~new_n729 & ~new_n730;
  assign new_n732 = new_n75 & ~new_n731;
  assign new_n733 = new_n421 & new_n445;
  assign new_n734 = ~_77_9_ & new_n450;
  assign new_n735 = _107_12_ & new_n456;
  assign new_n736 = _116_13_ & new_n459;
  assign new_n737 = _87_10_ & new_n461;
  assign new_n738 = _97_11_ & new_n464;
  assign new_n739 = _311_41_ & new_n466;
  assign new_n740 = _303_40_ & new_n469;
  assign new_n741 = _283_38_ & new_n471;
  assign new_n742 = _294_39_ & new_n473;
  assign new_n743 = ~new_n735 & ~new_n736;
  assign new_n744 = ~new_n737 & new_n743;
  assign new_n745 = ~new_n738 & new_n744;
  assign new_n746 = ~new_n739 & new_n745;
  assign new_n747 = ~new_n740 & new_n746;
  assign new_n748 = ~new_n741 & new_n747;
  assign new_n749 = ~new_n742 & new_n748;
  assign new_n750 = _33_3_ & new_n749;
  assign new_n751 = _50_6_ & new_n456;
  assign new_n752 = _159_21_ & new_n459;
  assign new_n753 = _68_8_ & new_n461;
  assign new_n754 = _58_7_ & new_n464;
  assign new_n755 = _132_17_ & new_n466;
  assign new_n756 = _137_18_ & new_n469;
  assign new_n757 = _150_20_ & new_n471;
  assign new_n758 = _143_19_ & new_n473;
  assign new_n759 = ~new_n751 & ~new_n752;
  assign new_n760 = ~new_n753 & new_n759;
  assign new_n761 = ~new_n754 & new_n760;
  assign new_n762 = ~new_n755 & new_n761;
  assign new_n763 = ~new_n756 & new_n762;
  assign new_n764 = ~new_n757 & new_n763;
  assign new_n765 = ~new_n758 & new_n764;
  assign new_n766 = ~_33_3_ & new_n765;
  assign new_n767 = ~new_n750 & ~new_n766;
  assign new_n768 = new_n449 & ~new_n767;
  assign new_n769 = ~new_n733 & ~new_n734;
  assign new_n770 = ~new_n768 & new_n769;
  assign new_n771 = new_n444 & new_n770;
  assign new_n772 = ~new_n443 & ~new_n731;
  assign new_n773 = ~new_n732 & ~new_n771;
  assign _384_1553_ = new_n772 | ~new_n773;
  assign new_n775 = ~new_n629 & ~new_n634;
  assign new_n776 = _330_46_ & new_n775;
  assign new_n777 = new_n235 & ~new_n287;
  assign new_n778 = new_n313 & ~new_n777;
  assign new_n779 = ~new_n313 & new_n777;
  assign new_n780 = ~new_n778 & ~new_n779;
  assign new_n781 = ~new_n634 & new_n635;
  assign new_n782 = ~new_n235 & ~new_n344;
  assign new_n783 = ~new_n781 & ~new_n782;
  assign new_n784 = new_n780 & ~new_n783;
  assign new_n785 = ~new_n780 & new_n783;
  assign new_n786 = ~new_n784 & ~new_n785;
  assign new_n787 = ~new_n776 & ~new_n786;
  assign new_n788 = new_n776 & new_n786;
  assign new_n789 = ~new_n787 & ~new_n788;
  assign new_n790 = ~new_n634 & ~new_n780;
  assign new_n791 = ~new_n629 & new_n790;
  assign new_n792 = _330_46_ & new_n791;
  assign new_n793 = new_n235 & ~new_n249;
  assign new_n794 = new_n274 & ~new_n793;
  assign new_n795 = ~new_n274 & new_n793;
  assign new_n796 = ~new_n794 & ~new_n795;
  assign new_n797 = ~new_n780 & new_n782;
  assign new_n798 = ~new_n780 & new_n781;
  assign new_n799 = ~new_n235 & ~new_n312;
  assign new_n800 = ~new_n797 & ~new_n798;
  assign new_n801 = ~new_n799 & new_n800;
  assign new_n802 = new_n796 & ~new_n801;
  assign new_n803 = ~new_n796 & new_n801;
  assign new_n804 = ~new_n802 & ~new_n803;
  assign new_n805 = ~new_n792 & ~new_n804;
  assign new_n806 = new_n792 & new_n804;
  assign new_n807 = ~new_n805 & ~new_n806;
  assign new_n808 = new_n625 & ~new_n789;
  assign new_n809 = ~new_n807 & new_n808;
  assign new_n810 = ~new_n641 & new_n809;
  assign new_n811 = ~new_n625 & ~new_n807;
  assign new_n812 = ~new_n810 & ~new_n811;
  assign new_n813 = new_n75 & ~new_n812;
  assign new_n814 = new_n647 & new_n796;
  assign new_n815 = ~_87_10_ & new_n656;
  assign new_n816 = _264_35_ & ~_270_36_;
  assign new_n817 = ~_264_35_ & _270_36_;
  assign new_n818 = ~new_n816 & ~new_n817;
  assign new_n819 = _250_33_ & ~_257_34_;
  assign new_n820 = ~_250_33_ & _257_34_;
  assign new_n821 = ~new_n819 & ~new_n820;
  assign new_n822 = new_n818 & ~new_n821;
  assign new_n823 = ~new_n818 & new_n821;
  assign new_n824 = ~new_n822 & ~new_n823;
  assign new_n825 = new_n655 & ~new_n824;
  assign new_n826 = ~new_n652 & ~new_n815;
  assign new_n827 = ~new_n825 & new_n826;
  assign new_n828 = new_n649 & ~new_n827;
  assign new_n829 = _116_13_ & new_n456;
  assign new_n830 = _283_38_ & new_n459;
  assign new_n831 = _107_12_ & new_n464;
  assign new_n832 = _317_42_ & new_n466;
  assign new_n833 = _311_41_ & new_n469;
  assign new_n834 = _294_39_ & new_n471;
  assign new_n835 = _303_40_ & new_n473;
  assign new_n836 = ~new_n829 & ~new_n830;
  assign new_n837 = ~new_n695 & new_n836;
  assign new_n838 = ~new_n831 & new_n837;
  assign new_n839 = ~new_n832 & new_n838;
  assign new_n840 = ~new_n833 & new_n839;
  assign new_n841 = ~new_n834 & new_n840;
  assign new_n842 = ~new_n835 & new_n841;
  assign new_n843 = _33_3_ & new_n842;
  assign new_n844 = _58_7_ & new_n456;
  assign new_n845 = _50_6_ & new_n459;
  assign new_n846 = _137_18_ & new_n466;
  assign new_n847 = _143_19_ & new_n469;
  assign new_n848 = _159_21_ & new_n471;
  assign new_n849 = _150_20_ & new_n473;
  assign new_n850 = ~new_n844 & ~new_n845;
  assign new_n851 = ~new_n462 & new_n850;
  assign new_n852 = ~new_n582 & new_n851;
  assign new_n853 = ~new_n846 & new_n852;
  assign new_n854 = ~new_n847 & new_n853;
  assign new_n855 = ~new_n848 & new_n854;
  assign new_n856 = ~new_n849 & new_n855;
  assign new_n857 = ~_33_3_ & new_n856;
  assign new_n858 = ~new_n843 & ~new_n857;
  assign new_n859 = new_n449 & ~new_n858;
  assign new_n860 = ~new_n814 & ~new_n828;
  assign new_n861 = ~new_n859 & new_n860;
  assign new_n862 = new_n444 & new_n861;
  assign new_n863 = ~new_n443 & ~new_n807;
  assign new_n864 = ~new_n813 & ~new_n862;
  assign _387_1616_ = new_n863 | ~new_n864;
  assign new_n866 = ~new_n671 & new_n824;
  assign new_n867 = new_n671 & ~new_n824;
  assign _358_1161_ = ~new_n866 & ~new_n867;
  assign _355_399_ = ~_87_10_ | new_n242;
  assign new_n870 = new_n775 & new_n783;
  assign new_n871 = _330_46_ & new_n870;
  assign _399_1428_ = ~new_n783 | new_n871;
  assign new_n873 = ~new_n438 & ~new_n547;
  assign new_n874 = new_n438 & new_n547;
  assign new_n875 = ~new_n873 & ~new_n874;
  assign new_n876 = new_n75 & ~new_n875;
  assign new_n877 = new_n445 & new_n536;
  assign new_n878 = ~_58_7_ & new_n450;
  assign new_n879 = _87_10_ & new_n456;
  assign new_n880 = _97_11_ & new_n459;
  assign new_n881 = _77_9_ & new_n464;
  assign new_n882 = _294_39_ & new_n466;
  assign new_n883 = _283_38_ & new_n469;
  assign new_n884 = _107_12_ & new_n471;
  assign new_n885 = _116_13_ & new_n473;
  assign new_n886 = ~new_n879 & ~new_n880;
  assign new_n887 = ~new_n753 & new_n886;
  assign new_n888 = ~new_n881 & new_n887;
  assign new_n889 = ~new_n882 & new_n888;
  assign new_n890 = ~new_n883 & new_n889;
  assign new_n891 = ~new_n884 & new_n890;
  assign new_n892 = ~new_n885 & new_n891;
  assign new_n893 = _33_3_ & new_n892;
  assign new_n894 = _150_20_ & new_n456;
  assign new_n895 = _143_19_ & new_n459;
  assign new_n896 = _50_6_ & new_n461;
  assign new_n897 = _159_21_ & new_n464;
  assign new_n898 = _125_15_ & new_n466;
  assign new_n899 = _128_16_ & new_n469;
  assign new_n900 = _137_18_ & new_n471;
  assign new_n901 = _132_17_ & new_n473;
  assign new_n902 = ~new_n894 & ~new_n895;
  assign new_n903 = ~new_n896 & new_n902;
  assign new_n904 = ~new_n897 & new_n903;
  assign new_n905 = ~new_n898 & new_n904;
  assign new_n906 = ~new_n899 & new_n905;
  assign new_n907 = ~new_n900 & new_n906;
  assign new_n908 = ~new_n901 & new_n907;
  assign new_n909 = ~_33_3_ & new_n908;
  assign new_n910 = ~new_n893 & ~new_n909;
  assign new_n911 = new_n449 & ~new_n910;
  assign new_n912 = ~new_n877 & ~new_n878;
  assign new_n913 = ~new_n911 & new_n912;
  assign new_n914 = new_n444 & new_n913;
  assign new_n915 = ~new_n443 & ~new_n547;
  assign new_n916 = ~new_n876 & ~new_n914;
  assign _378_1597_ = new_n915 | ~new_n916;
  assign new_n918 = ~_375_1624_ & _378_1597_;
  assign new_n919 = _375_1624_ & ~_378_1597_;
  assign new_n920 = ~new_n918 & ~new_n919;
  assign new_n921 = ~_381_1626_ & _384_1553_;
  assign new_n922 = _381_1626_ & ~_384_1553_;
  assign new_n923 = ~new_n921 & ~new_n922;
  assign new_n924 = new_n920 & ~new_n923;
  assign new_n925 = ~new_n920 & new_n923;
  assign new_n926 = ~new_n924 & ~new_n925;
  assign new_n927 = ~new_n643 & ~new_n789;
  assign new_n928 = new_n643 & new_n789;
  assign new_n929 = ~new_n927 & ~new_n928;
  assign new_n930 = new_n75 & ~new_n929;
  assign new_n931 = new_n647 & new_n780;
  assign new_n932 = ~_97_11_ & new_n656;
  assign new_n933 = ~new_n515 & new_n655;
  assign new_n934 = ~new_n652 & ~new_n932;
  assign new_n935 = ~new_n933 & new_n934;
  assign new_n936 = new_n649 & ~new_n935;
  assign new_n937 = _283_38_ & new_n456;
  assign new_n938 = _294_39_ & new_n459;
  assign new_n939 = _107_12_ & new_n461;
  assign new_n940 = _116_13_ & new_n464;
  assign new_n941 = _322_43_ & new_n466;
  assign new_n942 = _317_42_ & new_n469;
  assign new_n943 = _303_40_ & new_n471;
  assign new_n944 = _311_41_ & new_n473;
  assign new_n945 = ~new_n937 & ~new_n938;
  assign new_n946 = ~new_n939 & new_n945;
  assign new_n947 = ~new_n940 & new_n946;
  assign new_n948 = ~new_n941 & new_n947;
  assign new_n949 = ~new_n942 & new_n948;
  assign new_n950 = ~new_n943 & new_n949;
  assign new_n951 = ~new_n944 & new_n950;
  assign new_n952 = _33_3_ & new_n951;
  assign new_n953 = _68_8_ & new_n456;
  assign new_n954 = _58_7_ & new_n459;
  assign new_n955 = _143_19_ & new_n466;
  assign new_n956 = _150_20_ & new_n469;
  assign new_n957 = _50_6_ & new_n471;
  assign new_n958 = _159_21_ & new_n473;
  assign new_n959 = ~new_n953 & ~new_n954;
  assign new_n960 = ~new_n737 & new_n959;
  assign new_n961 = ~new_n881 & new_n960;
  assign new_n962 = ~new_n955 & new_n961;
  assign new_n963 = ~new_n956 & new_n962;
  assign new_n964 = ~new_n957 & new_n963;
  assign new_n965 = ~new_n958 & new_n964;
  assign new_n966 = ~_33_3_ & new_n965;
  assign new_n967 = ~new_n952 & ~new_n966;
  assign new_n968 = new_n449 & ~new_n967;
  assign new_n969 = ~new_n931 & ~new_n936;
  assign new_n970 = ~new_n968 & new_n969;
  assign new_n971 = new_n444 & new_n970;
  assign new_n972 = ~new_n443 & ~new_n789;
  assign new_n973 = ~new_n930 & ~new_n971;
  assign _390_1603_ = new_n972 | ~new_n973;
  assign new_n975 = ~_387_1616_ & _390_1603_;
  assign new_n976 = _387_1616_ & ~_390_1603_;
  assign new_n977 = ~new_n975 & ~new_n976;
  assign new_n978 = _330_46_ & new_n629;
  assign new_n979 = ~_330_46_ & ~new_n629;
  assign new_n980 = ~new_n978 & ~new_n979;
  assign new_n981 = new_n75 & ~new_n980;
  assign new_n982 = new_n629 & new_n647;
  assign new_n983 = new_n652 & _355_399_;
  assign new_n984 = ~_116_13_ & new_n656;
  assign new_n985 = ~_45_5_ & new_n719;
  assign new_n986 = _45_5_ & ~new_n524;
  assign new_n987 = ~new_n985 & ~new_n986;
  assign new_n988 = new_n655 & new_n987;
  assign new_n989 = ~new_n983 & ~new_n984;
  assign new_n990 = ~new_n988 & new_n989;
  assign new_n991 = new_n649 & ~new_n990;
  assign new_n992 = _303_40_ & new_n456;
  assign new_n993 = _311_41_ & new_n459;
  assign new_n994 = _283_38_ & new_n461;
  assign new_n995 = _294_39_ & new_n464;
  assign new_n996 = _329_45_ & new_n466;
  assign new_n997 = _326_44_ & new_n469;
  assign new_n998 = _317_42_ & new_n471;
  assign new_n999 = _322_43_ & new_n473;
  assign new_n1000 = ~new_n992 & ~new_n993;
  assign new_n1001 = ~new_n994 & new_n1000;
  assign new_n1002 = ~new_n995 & new_n1001;
  assign new_n1003 = ~new_n996 & new_n1002;
  assign new_n1004 = ~new_n997 & new_n1003;
  assign new_n1005 = ~new_n998 & new_n1004;
  assign new_n1006 = ~new_n999 & new_n1005;
  assign new_n1007 = _33_3_ & new_n1006;
  assign new_n1008 = _77_9_ & new_n459;
  assign new_n1009 = _159_21_ & new_n466;
  assign new_n1010 = _50_6_ & new_n469;
  assign new_n1011 = _68_8_ & new_n471;
  assign new_n1012 = _58_7_ & new_n473;
  assign new_n1013 = ~new_n879 & ~new_n1008;
  assign new_n1014 = ~new_n939 & new_n1013;
  assign new_n1015 = ~new_n738 & new_n1014;
  assign new_n1016 = ~new_n1009 & new_n1015;
  assign new_n1017 = ~new_n1010 & new_n1016;
  assign new_n1018 = ~new_n1011 & new_n1017;
  assign new_n1019 = ~new_n1012 & new_n1018;
  assign new_n1020 = ~_33_3_ & new_n1019;
  assign new_n1021 = ~new_n1007 & ~new_n1020;
  assign new_n1022 = new_n449 & ~new_n1021;
  assign new_n1023 = ~new_n982 & ~new_n991;
  assign new_n1024 = ~new_n1022 & new_n1023;
  assign new_n1025 = new_n444 & new_n1024;
  assign new_n1026 = ~new_n443 & ~new_n980;
  assign new_n1027 = ~new_n981 & ~new_n1025;
  assign _396_1504_ = new_n1026 | ~new_n1027;
  assign new_n1029 = ~_393_1605_ & _396_1504_;
  assign new_n1030 = _393_1605_ & ~_396_1504_;
  assign new_n1031 = ~new_n1029 & ~new_n1030;
  assign new_n1032 = new_n977 & ~new_n1031;
  assign new_n1033 = ~new_n977 & new_n1031;
  assign new_n1034 = ~new_n1032 & ~new_n1033;
  assign new_n1035 = new_n926 & ~new_n1034;
  assign new_n1036 = ~new_n926 & new_n1034;
  assign _402_1718_ = ~new_n1035 & ~new_n1036;
  assign _372_1243_ = new_n231 & new_n401;
  assign new_n1039 = _213_26_ & ~_343_47_;
  assign new_n1040 = _378_1597_ & ~new_n1039;
  assign new_n1041 = _375_1624_ & ~new_n1039;
  assign new_n1042 = ~new_n1040 & new_n1041;
  assign new_n1043 = new_n1040 & ~new_n1041;
  assign new_n1044 = ~new_n1042 & ~new_n1043;
  assign new_n1045 = _2897_49_ & new_n1039;
  assign new_n1046 = new_n1044 & new_n1045;
  assign new_n1047 = new_n923 & new_n1046;
  assign new_n1048 = new_n1044 & ~new_n1045;
  assign new_n1049 = ~new_n923 & new_n1048;
  assign new_n1050 = ~new_n1044 & ~new_n1045;
  assign new_n1051 = new_n923 & new_n1050;
  assign new_n1052 = ~new_n1044 & new_n1045;
  assign new_n1053 = ~new_n923 & new_n1052;
  assign new_n1054 = ~new_n1047 & ~new_n1049;
  assign new_n1055 = ~new_n1051 & new_n1054;
  assign new_n1056 = ~new_n1053 & new_n1055;
  assign new_n1057 = ~new_n1034 & ~new_n1056;
  assign new_n1058 = new_n1034 & new_n1056;
  assign _405_1717_ = new_n1057 | new_n1058;
  assign new_n1060 = ~_381_1626_ & ~_375_1624_;
  assign new_n1061 = ~_378_1597_ & new_n1060;
  assign new_n1062 = ~_384_1553_ & new_n1061;
  assign new_n1063 = ~_393_1605_ & ~_387_1616_;
  assign new_n1064 = ~_390_1603_ & new_n1063;
  assign new_n1065 = ~_396_1504_ & new_n1064;
  assign _407_1657_ = ~new_n1062 | ~new_n1065;
  assign new_n1067 = ~_375_1624_ & new_n1039;
  assign new_n1068 = ~_378_1597_ & new_n1067;
  assign new_n1069 = _407_1657_ & ~new_n1068;
  assign _409_1670_ = ~_213_26_ | ~new_n1069;
  assign new_n1071 = ~_264_35_ & ~_257_34_;
  assign new_n1072 = _250_33_ & ~new_n1071;
  assign new_n1073 = new_n651 & new_n1072;
  assign new_n1074 = _1_0_ & new_n76;
  assign new_n1075 = ~new_n651 & ~new_n1074;
  assign new_n1076 = _270_36_ & _116_13_;
  assign new_n1077 = _257_34_ & _97_11_;
  assign new_n1078 = _264_35_ & _107_12_;
  assign new_n1079 = _87_10_ & _250_33_;
  assign new_n1080 = ~new_n1076 & ~new_n1077;
  assign new_n1081 = ~new_n1078 & new_n1080;
  assign new_n1082 = ~new_n1079 & new_n1081;
  assign new_n1083 = _77_9_ & _244_32_;
  assign new_n1084 = _58_7_ & _232_30_;
  assign new_n1085 = _238_31_ & _68_8_;
  assign new_n1086 = _226_29_ & _50_6_;
  assign new_n1087 = ~new_n1083 & ~new_n1084;
  assign new_n1088 = ~new_n1085 & new_n1087;
  assign new_n1089 = ~new_n1086 & new_n1088;
  assign new_n1090 = new_n1082 & new_n1089;
  assign new_n1091 = new_n1075 & ~new_n1090;
  assign new_n1092 = new_n719 & new_n1074;
  assign new_n1093 = ~new_n1073 & ~new_n1091;
  assign _361_940_ = ~new_n1092 & new_n1093;
  assign new_n1095 = _116_13_ & ~new_n281;
  assign new_n1096 = new_n1074 & new_n1095;
  assign new_n1097 = ~_13_1_ & _1_0_;
  assign new_n1098 = ~new_n1074 & ~new_n1097;
  assign new_n1099 = new_n414 & ~new_n550;
  assign new_n1100 = ~new_n414 & new_n550;
  assign new_n1101 = ~new_n1099 & ~new_n1100;
  assign new_n1102 = _330_46_ & ~new_n1101;
  assign new_n1103 = new_n391 & ~new_n564;
  assign new_n1104 = ~new_n391 & new_n564;
  assign new_n1105 = ~new_n1103 & ~new_n1104;
  assign new_n1106 = ~new_n1102 & ~new_n1105;
  assign new_n1107 = new_n1102 & new_n1105;
  assign new_n1108 = ~new_n1106 & ~new_n1107;
  assign new_n1109 = new_n1098 & ~new_n1108;
  assign new_n1110 = _68_8_ & ~_50_6_;
  assign new_n1111 = _77_9_ & _50_6_;
  assign new_n1112 = ~new_n134 & new_n1111;
  assign new_n1113 = ~new_n1110 & ~new_n1112;
  assign new_n1114 = new_n1097 & ~new_n1113;
  assign new_n1115 = ~new_n1096 & ~new_n1109;
  assign _367_1585_ = new_n1114 | ~new_n1115;
endmodule


