module dec ( 
    \count0 , \count1 , \count2 , \count3 , \count4 , \count5 ,
    \count6 , \count7 ,
    \selectp10 , \selectp11 , \selectp12 , \selectp13 ,
    \selectp14 , \selectp15 , \selectp16 , \selectp17 ,
    \selectp18 , \selectp19 , \selectp110 , \selectp111 ,
    \selectp112 , \selectp113 , \selectp114 , \selectp115 ,
    \selectp116 , \selectp117 , \selectp118 , \selectp119 ,
    \selectp120 , \selectp121 , \selectp122 , \selectp123 ,
    \selectp124 , \selectp125 , \selectp126 , \selectp127 ,
    \selectp128 , \selectp129 , \selectp130 , \selectp131 ,
    \selectp132 , \selectp133 , \selectp134 , \selectp135 ,
    \selectp136 , \selectp137 , \selectp138 , \selectp139 ,
    \selectp140 , \selectp141 , \selectp142 , \selectp143 ,
    \selectp144 , \selectp145 , \selectp146 , \selectp147 ,
    \selectp148 , \selectp149 , \selectp150 , \selectp151 ,
    \selectp152 , \selectp153 , \selectp154 , \selectp155 ,
    \selectp156 , \selectp157 , \selectp158 , \selectp159 ,
    \selectp160 , \selectp161 , \selectp162 , \selectp163 ,
    \selectp164 , \selectp165 , \selectp166 , \selectp167 ,
    \selectp168 , \selectp169 , \selectp170 , \selectp171 ,
    \selectp172 , \selectp173 , \selectp174 , \selectp175 ,
    \selectp176 , \selectp177 , \selectp178 , \selectp179 ,
    \selectp180 , \selectp181 , \selectp182 , \selectp183 ,
    \selectp184 , \selectp185 , \selectp186 , \selectp187 ,
    \selectp188 , \selectp189 , \selectp190 , \selectp191 ,
    \selectp192 , \selectp193 , \selectp194 , \selectp195 ,
    \selectp196 , \selectp197 , \selectp198 , \selectp199 ,
    \selectp1100 , \selectp1101 , \selectp1102 , \selectp1103 ,
    \selectp1104 , \selectp1105 , \selectp1106 , \selectp1107 ,
    \selectp1108 , \selectp1109 , \selectp1110 , \selectp1111 ,
    \selectp1112 , \selectp1113 , \selectp1114 , \selectp1115 ,
    \selectp1116 , \selectp1117 , \selectp1118 , \selectp1119 ,
    \selectp1120 , \selectp1121 , \selectp1122 , \selectp1123 ,
    \selectp1124 , \selectp1125 , \selectp1126 , \selectp1127 ,
    \selectp20 , \selectp21 , \selectp22 , \selectp23 ,
    \selectp24 , \selectp25 , \selectp26 , \selectp27 ,
    \selectp28 , \selectp29 , \selectp210 , \selectp211 ,
    \selectp212 , \selectp213 , \selectp214 , \selectp215 ,
    \selectp216 , \selectp217 , \selectp218 , \selectp219 ,
    \selectp220 , \selectp221 , \selectp222 , \selectp223 ,
    \selectp224 , \selectp225 , \selectp226 , \selectp227 ,
    \selectp228 , \selectp229 , \selectp230 , \selectp231 ,
    \selectp232 , \selectp233 , \selectp234 , \selectp235 ,
    \selectp236 , \selectp237 , \selectp238 , \selectp239 ,
    \selectp240 , \selectp241 , \selectp242 , \selectp243 ,
    \selectp244 , \selectp245 , \selectp246 , \selectp247 ,
    \selectp248 , \selectp249 , \selectp250 , \selectp251 ,
    \selectp252 , \selectp253 , \selectp254 , \selectp255 ,
    \selectp256 , \selectp257 , \selectp258 , \selectp259 ,
    \selectp260 , \selectp261 , \selectp262 , \selectp263 ,
    \selectp264 , \selectp265 , \selectp266 , \selectp267 ,
    \selectp268 , \selectp269 , \selectp270 , \selectp271 ,
    \selectp272 , \selectp273 , \selectp274 , \selectp275 ,
    \selectp276 , \selectp277 , \selectp278 , \selectp279 ,
    \selectp280 , \selectp281 , \selectp282 , \selectp283 ,
    \selectp284 , \selectp285 , \selectp286 , \selectp287 ,
    \selectp288 , \selectp289 , \selectp290 , \selectp291 ,
    \selectp292 , \selectp293 , \selectp294 , \selectp295 ,
    \selectp296 , \selectp297 , \selectp298 , \selectp299 ,
    \selectp2100 , \selectp2101 , \selectp2102 , \selectp2103 ,
    \selectp2104 , \selectp2105 , \selectp2106 , \selectp2107 ,
    \selectp2108 , \selectp2109 , \selectp2110 , \selectp2111 ,
    \selectp2112 , \selectp2113 , \selectp2114 , \selectp2115 ,
    \selectp2116 , \selectp2117 , \selectp2118 , \selectp2119 ,
    \selectp2120 , \selectp2121 , \selectp2122 , \selectp2123 ,
    \selectp2124 , \selectp2125 , \selectp2126 , \selectp2127   );
  input  \count0 , \count1 , \count2 , \count3 , \count4 ,
    \count5 , \count6 , \count7 ;
  output \selectp10 , \selectp11 , \selectp12 , \selectp13 ,
    \selectp14 , \selectp15 , \selectp16 , \selectp17 ,
    \selectp18 , \selectp19 , \selectp110 , \selectp111 ,
    \selectp112 , \selectp113 , \selectp114 , \selectp115 ,
    \selectp116 , \selectp117 , \selectp118 , \selectp119 ,
    \selectp120 , \selectp121 , \selectp122 , \selectp123 ,
    \selectp124 , \selectp125 , \selectp126 , \selectp127 ,
    \selectp128 , \selectp129 , \selectp130 , \selectp131 ,
    \selectp132 , \selectp133 , \selectp134 , \selectp135 ,
    \selectp136 , \selectp137 , \selectp138 , \selectp139 ,
    \selectp140 , \selectp141 , \selectp142 , \selectp143 ,
    \selectp144 , \selectp145 , \selectp146 , \selectp147 ,
    \selectp148 , \selectp149 , \selectp150 , \selectp151 ,
    \selectp152 , \selectp153 , \selectp154 , \selectp155 ,
    \selectp156 , \selectp157 , \selectp158 , \selectp159 ,
    \selectp160 , \selectp161 , \selectp162 , \selectp163 ,
    \selectp164 , \selectp165 , \selectp166 , \selectp167 ,
    \selectp168 , \selectp169 , \selectp170 , \selectp171 ,
    \selectp172 , \selectp173 , \selectp174 , \selectp175 ,
    \selectp176 , \selectp177 , \selectp178 , \selectp179 ,
    \selectp180 , \selectp181 , \selectp182 , \selectp183 ,
    \selectp184 , \selectp185 , \selectp186 , \selectp187 ,
    \selectp188 , \selectp189 , \selectp190 , \selectp191 ,
    \selectp192 , \selectp193 , \selectp194 , \selectp195 ,
    \selectp196 , \selectp197 , \selectp198 , \selectp199 ,
    \selectp1100 , \selectp1101 , \selectp1102 , \selectp1103 ,
    \selectp1104 , \selectp1105 , \selectp1106 , \selectp1107 ,
    \selectp1108 , \selectp1109 , \selectp1110 , \selectp1111 ,
    \selectp1112 , \selectp1113 , \selectp1114 , \selectp1115 ,
    \selectp1116 , \selectp1117 , \selectp1118 , \selectp1119 ,
    \selectp1120 , \selectp1121 , \selectp1122 , \selectp1123 ,
    \selectp1124 , \selectp1125 , \selectp1126 , \selectp1127 ,
    \selectp20 , \selectp21 , \selectp22 , \selectp23 ,
    \selectp24 , \selectp25 , \selectp26 , \selectp27 ,
    \selectp28 , \selectp29 , \selectp210 , \selectp211 ,
    \selectp212 , \selectp213 , \selectp214 , \selectp215 ,
    \selectp216 , \selectp217 , \selectp218 , \selectp219 ,
    \selectp220 , \selectp221 , \selectp222 , \selectp223 ,
    \selectp224 , \selectp225 , \selectp226 , \selectp227 ,
    \selectp228 , \selectp229 , \selectp230 , \selectp231 ,
    \selectp232 , \selectp233 , \selectp234 , \selectp235 ,
    \selectp236 , \selectp237 , \selectp238 , \selectp239 ,
    \selectp240 , \selectp241 , \selectp242 , \selectp243 ,
    \selectp244 , \selectp245 , \selectp246 , \selectp247 ,
    \selectp248 , \selectp249 , \selectp250 , \selectp251 ,
    \selectp252 , \selectp253 , \selectp254 , \selectp255 ,
    \selectp256 , \selectp257 , \selectp258 , \selectp259 ,
    \selectp260 , \selectp261 , \selectp262 , \selectp263 ,
    \selectp264 , \selectp265 , \selectp266 , \selectp267 ,
    \selectp268 , \selectp269 , \selectp270 , \selectp271 ,
    \selectp272 , \selectp273 , \selectp274 , \selectp275 ,
    \selectp276 , \selectp277 , \selectp278 , \selectp279 ,
    \selectp280 , \selectp281 , \selectp282 , \selectp283 ,
    \selectp284 , \selectp285 , \selectp286 , \selectp287 ,
    \selectp288 , \selectp289 , \selectp290 , \selectp291 ,
    \selectp292 , \selectp293 , \selectp294 , \selectp295 ,
    \selectp296 , \selectp297 , \selectp298 , \selectp299 ,
    \selectp2100 , \selectp2101 , \selectp2102 , \selectp2103 ,
    \selectp2104 , \selectp2105 , \selectp2106 , \selectp2107 ,
    \selectp2108 , \selectp2109 , \selectp2110 , \selectp2111 ,
    \selectp2112 , \selectp2113 , \selectp2114 , \selectp2115 ,
    \selectp2116 , \selectp2117 , \selectp2118 , \selectp2119 ,
    \selectp2120 , \selectp2121 , \selectp2122 , \selectp2123 ,
    \selectp2124 , \selectp2125 , \selectp2126 , \selectp2127 ;
  wire n265, n266, n267, n268, n269, n270, n272, n273, n275, n276, n278,
    n280, n281, n283, n284, n286, n288, n290, n291, n293, n295, n296, n298,
    n300, n302, n304, n306, n308, n309, n326, n327, n344, n345, n362, n363,
    n380, n397, n414, n431, n432, n449, n466, n483, n500, n501, n518, n535,
    n552;
  assign n265 = ~\count4  & ~\count5 ;
  assign n266 = ~\count6  & \count7 ;
  assign n267 = n265 & n266;
  assign n268 = ~\count0  & ~\count2 ;
  assign n269 = ~\count1  & ~\count3 ;
  assign n270 = n268 & n269;
  assign \selectp10  = n267 & n270;
  assign n272 = \count0  & ~\count2 ;
  assign n273 = n269 & n272;
  assign \selectp11  = n267 & n273;
  assign n275 = \count1  & ~\count3 ;
  assign n276 = n268 & n275;
  assign \selectp12  = n267 & n276;
  assign n278 = n272 & n275;
  assign \selectp13  = n267 & n278;
  assign n280 = ~\count0  & \count2 ;
  assign n281 = n269 & n280;
  assign \selectp14  = n267 & n281;
  assign n283 = \count0  & \count2 ;
  assign n284 = n269 & n283;
  assign \selectp15  = n267 & n284;
  assign n286 = n275 & n280;
  assign \selectp16  = n267 & n286;
  assign n288 = n275 & n283;
  assign \selectp17  = n267 & n288;
  assign n290 = ~\count1  & \count3 ;
  assign n291 = n268 & n290;
  assign \selectp18  = n267 & n291;
  assign n293 = n272 & n290;
  assign \selectp19  = n267 & n293;
  assign n295 = \count1  & \count3 ;
  assign n296 = n268 & n295;
  assign \selectp110  = n267 & n296;
  assign n298 = n272 & n295;
  assign \selectp111  = n267 & n298;
  assign n300 = n280 & n290;
  assign \selectp112  = n267 & n300;
  assign n302 = n283 & n290;
  assign \selectp113  = n267 & n302;
  assign n304 = n280 & n295;
  assign \selectp114  = n267 & n304;
  assign n306 = n283 & n295;
  assign \selectp115  = n267 & n306;
  assign n308 = \count4  & ~\count5 ;
  assign n309 = n266 & n308;
  assign \selectp116  = n270 & n309;
  assign \selectp117  = n273 & n309;
  assign \selectp118  = n276 & n309;
  assign \selectp119  = n278 & n309;
  assign \selectp120  = n281 & n309;
  assign \selectp121  = n284 & n309;
  assign \selectp122  = n286 & n309;
  assign \selectp123  = n288 & n309;
  assign \selectp124  = n291 & n309;
  assign \selectp125  = n293 & n309;
  assign \selectp126  = n296 & n309;
  assign \selectp127  = n298 & n309;
  assign \selectp128  = n300 & n309;
  assign \selectp129  = n302 & n309;
  assign \selectp130  = n304 & n309;
  assign \selectp131  = n306 & n309;
  assign n326 = ~\count4  & \count5 ;
  assign n327 = n266 & n326;
  assign \selectp132  = n270 & n327;
  assign \selectp133  = n273 & n327;
  assign \selectp134  = n276 & n327;
  assign \selectp135  = n278 & n327;
  assign \selectp136  = n281 & n327;
  assign \selectp137  = n284 & n327;
  assign \selectp138  = n286 & n327;
  assign \selectp139  = n288 & n327;
  assign \selectp140  = n291 & n327;
  assign \selectp141  = n293 & n327;
  assign \selectp142  = n296 & n327;
  assign \selectp143  = n298 & n327;
  assign \selectp144  = n300 & n327;
  assign \selectp145  = n302 & n327;
  assign \selectp146  = n304 & n327;
  assign \selectp147  = n306 & n327;
  assign n344 = \count4  & \count5 ;
  assign n345 = n266 & n344;
  assign \selectp148  = n270 & n345;
  assign \selectp149  = n273 & n345;
  assign \selectp150  = n276 & n345;
  assign \selectp151  = n278 & n345;
  assign \selectp152  = n281 & n345;
  assign \selectp153  = n284 & n345;
  assign \selectp154  = n286 & n345;
  assign \selectp155  = n288 & n345;
  assign \selectp156  = n291 & n345;
  assign \selectp157  = n293 & n345;
  assign \selectp158  = n296 & n345;
  assign \selectp159  = n298 & n345;
  assign \selectp160  = n300 & n345;
  assign \selectp161  = n302 & n345;
  assign \selectp162  = n304 & n345;
  assign \selectp163  = n306 & n345;
  assign n362 = \count6  & \count7 ;
  assign n363 = n265 & n362;
  assign \selectp164  = n270 & n363;
  assign \selectp165  = n273 & n363;
  assign \selectp166  = n276 & n363;
  assign \selectp167  = n278 & n363;
  assign \selectp168  = n281 & n363;
  assign \selectp169  = n284 & n363;
  assign \selectp170  = n286 & n363;
  assign \selectp171  = n288 & n363;
  assign \selectp172  = n291 & n363;
  assign \selectp173  = n293 & n363;
  assign \selectp174  = n296 & n363;
  assign \selectp175  = n298 & n363;
  assign \selectp176  = n300 & n363;
  assign \selectp177  = n302 & n363;
  assign \selectp178  = n304 & n363;
  assign \selectp179  = n306 & n363;
  assign n380 = n308 & n362;
  assign \selectp180  = n270 & n380;
  assign \selectp181  = n273 & n380;
  assign \selectp182  = n276 & n380;
  assign \selectp183  = n278 & n380;
  assign \selectp184  = n281 & n380;
  assign \selectp185  = n284 & n380;
  assign \selectp186  = n286 & n380;
  assign \selectp187  = n288 & n380;
  assign \selectp188  = n291 & n380;
  assign \selectp189  = n293 & n380;
  assign \selectp190  = n296 & n380;
  assign \selectp191  = n298 & n380;
  assign \selectp192  = n300 & n380;
  assign \selectp193  = n302 & n380;
  assign \selectp194  = n304 & n380;
  assign \selectp195  = n306 & n380;
  assign n397 = n326 & n362;
  assign \selectp196  = n270 & n397;
  assign \selectp197  = n273 & n397;
  assign \selectp198  = n276 & n397;
  assign \selectp199  = n278 & n397;
  assign \selectp1100  = n281 & n397;
  assign \selectp1101  = n284 & n397;
  assign \selectp1102  = n286 & n397;
  assign \selectp1103  = n288 & n397;
  assign \selectp1104  = n291 & n397;
  assign \selectp1105  = n293 & n397;
  assign \selectp1106  = n296 & n397;
  assign \selectp1107  = n298 & n397;
  assign \selectp1108  = n300 & n397;
  assign \selectp1109  = n302 & n397;
  assign \selectp1110  = n304 & n397;
  assign \selectp1111  = n306 & n397;
  assign n414 = n344 & n362;
  assign \selectp1112  = n270 & n414;
  assign \selectp1113  = n273 & n414;
  assign \selectp1114  = n276 & n414;
  assign \selectp1115  = n278 & n414;
  assign \selectp1116  = n281 & n414;
  assign \selectp1117  = n284 & n414;
  assign \selectp1118  = n286 & n414;
  assign \selectp1119  = n288 & n414;
  assign \selectp1120  = n291 & n414;
  assign \selectp1121  = n293 & n414;
  assign \selectp1122  = n296 & n414;
  assign \selectp1123  = n298 & n414;
  assign \selectp1124  = n300 & n414;
  assign \selectp1125  = n302 & n414;
  assign \selectp1126  = n304 & n414;
  assign \selectp1127  = n306 & n414;
  assign n431 = ~\count6  & ~\count7 ;
  assign n432 = n265 & n431;
  assign \selectp20  = n270 & n432;
  assign \selectp21  = n273 & n432;
  assign \selectp22  = n276 & n432;
  assign \selectp23  = n278 & n432;
  assign \selectp24  = n281 & n432;
  assign \selectp25  = n284 & n432;
  assign \selectp26  = n286 & n432;
  assign \selectp27  = n288 & n432;
  assign \selectp28  = n291 & n432;
  assign \selectp29  = n293 & n432;
  assign \selectp210  = n296 & n432;
  assign \selectp211  = n298 & n432;
  assign \selectp212  = n300 & n432;
  assign \selectp213  = n302 & n432;
  assign \selectp214  = n304 & n432;
  assign \selectp215  = n306 & n432;
  assign n449 = n308 & n431;
  assign \selectp216  = n270 & n449;
  assign \selectp217  = n273 & n449;
  assign \selectp218  = n276 & n449;
  assign \selectp219  = n278 & n449;
  assign \selectp220  = n281 & n449;
  assign \selectp221  = n284 & n449;
  assign \selectp222  = n286 & n449;
  assign \selectp223  = n288 & n449;
  assign \selectp224  = n291 & n449;
  assign \selectp225  = n293 & n449;
  assign \selectp226  = n296 & n449;
  assign \selectp227  = n298 & n449;
  assign \selectp228  = n300 & n449;
  assign \selectp229  = n302 & n449;
  assign \selectp230  = n304 & n449;
  assign \selectp231  = n306 & n449;
  assign n466 = n326 & n431;
  assign \selectp232  = n270 & n466;
  assign \selectp233  = n273 & n466;
  assign \selectp234  = n276 & n466;
  assign \selectp235  = n278 & n466;
  assign \selectp236  = n281 & n466;
  assign \selectp237  = n284 & n466;
  assign \selectp238  = n286 & n466;
  assign \selectp239  = n288 & n466;
  assign \selectp240  = n291 & n466;
  assign \selectp241  = n293 & n466;
  assign \selectp242  = n296 & n466;
  assign \selectp243  = n298 & n466;
  assign \selectp244  = n300 & n466;
  assign \selectp245  = n302 & n466;
  assign \selectp246  = n304 & n466;
  assign \selectp247  = n306 & n466;
  assign n483 = n344 & n431;
  assign \selectp248  = n270 & n483;
  assign \selectp249  = n273 & n483;
  assign \selectp250  = n276 & n483;
  assign \selectp251  = n278 & n483;
  assign \selectp252  = n281 & n483;
  assign \selectp253  = n284 & n483;
  assign \selectp254  = n286 & n483;
  assign \selectp255  = n288 & n483;
  assign \selectp256  = n291 & n483;
  assign \selectp257  = n293 & n483;
  assign \selectp258  = n296 & n483;
  assign \selectp259  = n298 & n483;
  assign \selectp260  = n300 & n483;
  assign \selectp261  = n302 & n483;
  assign \selectp262  = n304 & n483;
  assign \selectp263  = n306 & n483;
  assign n500 = \count6  & ~\count7 ;
  assign n501 = n265 & n500;
  assign \selectp264  = n270 & n501;
  assign \selectp265  = n273 & n501;
  assign \selectp266  = n276 & n501;
  assign \selectp267  = n278 & n501;
  assign \selectp268  = n281 & n501;
  assign \selectp269  = n284 & n501;
  assign \selectp270  = n286 & n501;
  assign \selectp271  = n288 & n501;
  assign \selectp272  = n291 & n501;
  assign \selectp273  = n293 & n501;
  assign \selectp274  = n296 & n501;
  assign \selectp275  = n298 & n501;
  assign \selectp276  = n300 & n501;
  assign \selectp277  = n302 & n501;
  assign \selectp278  = n304 & n501;
  assign \selectp279  = n306 & n501;
  assign n518 = n308 & n500;
  assign \selectp280  = n270 & n518;
  assign \selectp281  = n273 & n518;
  assign \selectp282  = n276 & n518;
  assign \selectp283  = n278 & n518;
  assign \selectp284  = n281 & n518;
  assign \selectp285  = n284 & n518;
  assign \selectp286  = n286 & n518;
  assign \selectp287  = n288 & n518;
  assign \selectp288  = n291 & n518;
  assign \selectp289  = n293 & n518;
  assign \selectp290  = n296 & n518;
  assign \selectp291  = n298 & n518;
  assign \selectp292  = n300 & n518;
  assign \selectp293  = n302 & n518;
  assign \selectp294  = n304 & n518;
  assign \selectp295  = n306 & n518;
  assign n535 = n326 & n500;
  assign \selectp296  = n270 & n535;
  assign \selectp297  = n273 & n535;
  assign \selectp298  = n276 & n535;
  assign \selectp299  = n278 & n535;
  assign \selectp2100  = n281 & n535;
  assign \selectp2101  = n284 & n535;
  assign \selectp2102  = n286 & n535;
  assign \selectp2103  = n288 & n535;
  assign \selectp2104  = n291 & n535;
  assign \selectp2105  = n293 & n535;
  assign \selectp2106  = n296 & n535;
  assign \selectp2107  = n298 & n535;
  assign \selectp2108  = n300 & n535;
  assign \selectp2109  = n302 & n535;
  assign \selectp2110  = n304 & n535;
  assign \selectp2111  = n306 & n535;
  assign n552 = n344 & n500;
  assign \selectp2112  = n270 & n552;
  assign \selectp2113  = n273 & n552;
  assign \selectp2114  = n276 & n552;
  assign \selectp2115  = n278 & n552;
  assign \selectp2116  = n281 & n552;
  assign \selectp2117  = n284 & n552;
  assign \selectp2118  = n286 & n552;
  assign \selectp2119  = n288 & n552;
  assign \selectp2120  = n291 & n552;
  assign \selectp2121  = n293 & n552;
  assign \selectp2122  = n296 & n552;
  assign \selectp2123  = n298 & n552;
  assign \selectp2124  = n300 & n552;
  assign \selectp2125  = n302 & n552;
  assign \selectp2126  = n304 & n552;
  assign \selectp2127  = n306 & n552;
endmodule


